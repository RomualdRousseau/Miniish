// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 27 2022 09:13:54

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    led,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    input [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output [7:0] led;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__33435;
    wire N__33434;
    wire N__33433;
    wire N__33424;
    wire N__33423;
    wire N__33422;
    wire N__33415;
    wire N__33414;
    wire N__33413;
    wire N__33406;
    wire N__33405;
    wire N__33404;
    wire N__33397;
    wire N__33396;
    wire N__33395;
    wire N__33388;
    wire N__33387;
    wire N__33386;
    wire N__33379;
    wire N__33378;
    wire N__33377;
    wire N__33370;
    wire N__33369;
    wire N__33368;
    wire N__33361;
    wire N__33360;
    wire N__33359;
    wire N__33352;
    wire N__33351;
    wire N__33350;
    wire N__33343;
    wire N__33342;
    wire N__33341;
    wire N__33334;
    wire N__33333;
    wire N__33332;
    wire N__33325;
    wire N__33324;
    wire N__33323;
    wire N__33316;
    wire N__33315;
    wire N__33314;
    wire N__33307;
    wire N__33306;
    wire N__33305;
    wire N__33298;
    wire N__33297;
    wire N__33296;
    wire N__33289;
    wire N__33288;
    wire N__33287;
    wire N__33280;
    wire N__33279;
    wire N__33278;
    wire N__33271;
    wire N__33270;
    wire N__33269;
    wire N__33262;
    wire N__33261;
    wire N__33260;
    wire N__33253;
    wire N__33252;
    wire N__33251;
    wire N__33244;
    wire N__33243;
    wire N__33242;
    wire N__33235;
    wire N__33234;
    wire N__33233;
    wire N__33226;
    wire N__33225;
    wire N__33224;
    wire N__33217;
    wire N__33216;
    wire N__33215;
    wire N__33208;
    wire N__33207;
    wire N__33206;
    wire N__33199;
    wire N__33198;
    wire N__33197;
    wire N__33190;
    wire N__33189;
    wire N__33188;
    wire N__33181;
    wire N__33180;
    wire N__33179;
    wire N__33172;
    wire N__33171;
    wire N__33170;
    wire N__33163;
    wire N__33162;
    wire N__33161;
    wire N__33154;
    wire N__33153;
    wire N__33152;
    wire N__33145;
    wire N__33144;
    wire N__33143;
    wire N__33136;
    wire N__33135;
    wire N__33134;
    wire N__33127;
    wire N__33126;
    wire N__33125;
    wire N__33118;
    wire N__33117;
    wire N__33116;
    wire N__33109;
    wire N__33108;
    wire N__33107;
    wire N__33100;
    wire N__33099;
    wire N__33098;
    wire N__33091;
    wire N__33090;
    wire N__33089;
    wire N__33082;
    wire N__33081;
    wire N__33080;
    wire N__33073;
    wire N__33072;
    wire N__33071;
    wire N__33064;
    wire N__33063;
    wire N__33062;
    wire N__33055;
    wire N__33054;
    wire N__33053;
    wire N__33046;
    wire N__33045;
    wire N__33044;
    wire N__33037;
    wire N__33036;
    wire N__33035;
    wire N__33028;
    wire N__33027;
    wire N__33026;
    wire N__33019;
    wire N__33018;
    wire N__33017;
    wire N__33010;
    wire N__33009;
    wire N__33008;
    wire N__33001;
    wire N__33000;
    wire N__32999;
    wire N__32992;
    wire N__32991;
    wire N__32990;
    wire N__32983;
    wire N__32982;
    wire N__32981;
    wire N__32974;
    wire N__32973;
    wire N__32972;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32941;
    wire N__32936;
    wire N__32933;
    wire N__32932;
    wire N__32927;
    wire N__32924;
    wire N__32919;
    wire N__32916;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32908;
    wire N__32905;
    wire N__32904;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32896;
    wire N__32893;
    wire N__32892;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32884;
    wire N__32879;
    wire N__32876;
    wire N__32875;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32858;
    wire N__32855;
    wire N__32850;
    wire N__32845;
    wire N__32840;
    wire N__32833;
    wire N__32830;
    wire N__32827;
    wire N__32826;
    wire N__32823;
    wire N__32820;
    wire N__32819;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32800;
    wire N__32797;
    wire N__32794;
    wire N__32791;
    wire N__32786;
    wire N__32783;
    wire N__32780;
    wire N__32777;
    wire N__32768;
    wire N__32763;
    wire N__32760;
    wire N__32759;
    wire N__32758;
    wire N__32757;
    wire N__32756;
    wire N__32755;
    wire N__32754;
    wire N__32753;
    wire N__32752;
    wire N__32751;
    wire N__32750;
    wire N__32749;
    wire N__32748;
    wire N__32741;
    wire N__32736;
    wire N__32735;
    wire N__32734;
    wire N__32733;
    wire N__32724;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32702;
    wire N__32697;
    wire N__32694;
    wire N__32691;
    wire N__32682;
    wire N__32679;
    wire N__32676;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32664;
    wire N__32663;
    wire N__32662;
    wire N__32661;
    wire N__32660;
    wire N__32659;
    wire N__32658;
    wire N__32657;
    wire N__32656;
    wire N__32655;
    wire N__32654;
    wire N__32653;
    wire N__32652;
    wire N__32651;
    wire N__32650;
    wire N__32649;
    wire N__32648;
    wire N__32647;
    wire N__32646;
    wire N__32645;
    wire N__32644;
    wire N__32643;
    wire N__32642;
    wire N__32641;
    wire N__32640;
    wire N__32639;
    wire N__32638;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32634;
    wire N__32633;
    wire N__32632;
    wire N__32631;
    wire N__32630;
    wire N__32629;
    wire N__32628;
    wire N__32627;
    wire N__32626;
    wire N__32625;
    wire N__32624;
    wire N__32623;
    wire N__32622;
    wire N__32621;
    wire N__32620;
    wire N__32619;
    wire N__32618;
    wire N__32617;
    wire N__32616;
    wire N__32615;
    wire N__32614;
    wire N__32613;
    wire N__32612;
    wire N__32611;
    wire N__32610;
    wire N__32609;
    wire N__32608;
    wire N__32607;
    wire N__32606;
    wire N__32605;
    wire N__32604;
    wire N__32603;
    wire N__32602;
    wire N__32601;
    wire N__32600;
    wire N__32599;
    wire N__32598;
    wire N__32597;
    wire N__32596;
    wire N__32595;
    wire N__32594;
    wire N__32593;
    wire N__32592;
    wire N__32591;
    wire N__32590;
    wire N__32589;
    wire N__32588;
    wire N__32587;
    wire N__32586;
    wire N__32585;
    wire N__32584;
    wire N__32583;
    wire N__32582;
    wire N__32581;
    wire N__32580;
    wire N__32579;
    wire N__32578;
    wire N__32577;
    wire N__32576;
    wire N__32575;
    wire N__32574;
    wire N__32573;
    wire N__32572;
    wire N__32571;
    wire N__32570;
    wire N__32569;
    wire N__32568;
    wire N__32567;
    wire N__32566;
    wire N__32565;
    wire N__32564;
    wire N__32563;
    wire N__32562;
    wire N__32561;
    wire N__32560;
    wire N__32559;
    wire N__32558;
    wire N__32557;
    wire N__32556;
    wire N__32555;
    wire N__32554;
    wire N__32553;
    wire N__32552;
    wire N__32551;
    wire N__32550;
    wire N__32549;
    wire N__32548;
    wire N__32547;
    wire N__32546;
    wire N__32545;
    wire N__32544;
    wire N__32543;
    wire N__32542;
    wire N__32541;
    wire N__32540;
    wire N__32539;
    wire N__32538;
    wire N__32537;
    wire N__32536;
    wire N__32535;
    wire N__32534;
    wire N__32533;
    wire N__32532;
    wire N__32531;
    wire N__32530;
    wire N__32529;
    wire N__32528;
    wire N__32527;
    wire N__32526;
    wire N__32525;
    wire N__32524;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32234;
    wire N__32233;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32177;
    wire N__32176;
    wire N__32175;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32142;
    wire N__32141;
    wire N__32140;
    wire N__32137;
    wire N__32136;
    wire N__32135;
    wire N__32134;
    wire N__32133;
    wire N__32132;
    wire N__32131;
    wire N__32130;
    wire N__32129;
    wire N__32128;
    wire N__32125;
    wire N__32124;
    wire N__32123;
    wire N__32120;
    wire N__32119;
    wire N__32116;
    wire N__32113;
    wire N__32106;
    wire N__32103;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32079;
    wire N__32078;
    wire N__32077;
    wire N__32076;
    wire N__32075;
    wire N__32072;
    wire N__32063;
    wire N__32060;
    wire N__32053;
    wire N__32048;
    wire N__32045;
    wire N__32042;
    wire N__32035;
    wire N__32032;
    wire N__32029;
    wire N__32026;
    wire N__32021;
    wire N__32016;
    wire N__32011;
    wire N__32008;
    wire N__32005;
    wire N__32002;
    wire N__31999;
    wire N__31996;
    wire N__31993;
    wire N__31990;
    wire N__31985;
    wire N__31980;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31966;
    wire N__31965;
    wire N__31964;
    wire N__31961;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31948;
    wire N__31945;
    wire N__31940;
    wire N__31939;
    wire N__31936;
    wire N__31935;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31923;
    wire N__31920;
    wire N__31919;
    wire N__31916;
    wire N__31913;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31901;
    wire N__31898;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31885;
    wire N__31884;
    wire N__31883;
    wire N__31882;
    wire N__31879;
    wire N__31872;
    wire N__31869;
    wire N__31864;
    wire N__31857;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31845;
    wire N__31842;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31825;
    wire N__31820;
    wire N__31815;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31593;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31538;
    wire N__31537;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31522;
    wire N__31519;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31490;
    wire N__31487;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31442;
    wire N__31441;
    wire N__31438;
    wire N__31435;
    wire N__31432;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31358;
    wire N__31357;
    wire N__31356;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31342;
    wire N__31339;
    wire N__31334;
    wire N__31331;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31323;
    wire N__31322;
    wire N__31319;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31300;
    wire N__31297;
    wire N__31296;
    wire N__31295;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31264;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31202;
    wire N__31199;
    wire N__31196;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31104;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31061;
    wire N__31058;
    wire N__31055;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31040;
    wire N__31037;
    wire N__31034;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30977;
    wire N__30974;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30935;
    wire N__30934;
    wire N__30931;
    wire N__30930;
    wire N__30929;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30915;
    wire N__30914;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30863;
    wire N__30858;
    wire N__30855;
    wire N__30850;
    wire N__30847;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30812;
    wire N__30809;
    wire N__30804;
    wire N__30801;
    wire N__30796;
    wire N__30793;
    wire N__30786;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30762;
    wire N__30761;
    wire N__30756;
    wire N__30755;
    wire N__30754;
    wire N__30753;
    wire N__30752;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30740;
    wire N__30739;
    wire N__30734;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30720;
    wire N__30713;
    wire N__30708;
    wire N__30705;
    wire N__30704;
    wire N__30701;
    wire N__30700;
    wire N__30699;
    wire N__30698;
    wire N__30697;
    wire N__30694;
    wire N__30689;
    wire N__30686;
    wire N__30685;
    wire N__30682;
    wire N__30681;
    wire N__30678;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30663;
    wire N__30658;
    wire N__30657;
    wire N__30654;
    wire N__30653;
    wire N__30648;
    wire N__30643;
    wire N__30640;
    wire N__30635;
    wire N__30632;
    wire N__30627;
    wire N__30624;
    wire N__30615;
    wire N__30614;
    wire N__30611;
    wire N__30610;
    wire N__30607;
    wire N__30606;
    wire N__30605;
    wire N__30600;
    wire N__30595;
    wire N__30594;
    wire N__30593;
    wire N__30592;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30577;
    wire N__30574;
    wire N__30573;
    wire N__30572;
    wire N__30569;
    wire N__30564;
    wire N__30561;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30542;
    wire N__30539;
    wire N__30528;
    wire N__30527;
    wire N__30526;
    wire N__30521;
    wire N__30520;
    wire N__30519;
    wire N__30516;
    wire N__30515;
    wire N__30514;
    wire N__30513;
    wire N__30510;
    wire N__30505;
    wire N__30500;
    wire N__30497;
    wire N__30494;
    wire N__30491;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30481;
    wire N__30480;
    wire N__30477;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30447;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30417;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30357;
    wire N__30354;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30281;
    wire N__30280;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30249;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30107;
    wire N__30106;
    wire N__30105;
    wire N__30102;
    wire N__30101;
    wire N__30100;
    wire N__30097;
    wire N__30096;
    wire N__30095;
    wire N__30092;
    wire N__30091;
    wire N__30090;
    wire N__30089;
    wire N__30088;
    wire N__30085;
    wire N__30082;
    wire N__30077;
    wire N__30076;
    wire N__30073;
    wire N__30068;
    wire N__30065;
    wire N__30060;
    wire N__30057;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30045;
    wire N__30042;
    wire N__30037;
    wire N__30036;
    wire N__30035;
    wire N__30032;
    wire N__30027;
    wire N__30024;
    wire N__30015;
    wire N__30012;
    wire N__30007;
    wire N__30002;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29960;
    wire N__29959;
    wire N__29956;
    wire N__29951;
    wire N__29946;
    wire N__29943;
    wire N__29940;
    wire N__29937;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29927;
    wire N__29922;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29910;
    wire N__29909;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29892;
    wire N__29889;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29879;
    wire N__29876;
    wire N__29875;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29859;
    wire N__29856;
    wire N__29853;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29843;
    wire N__29842;
    wire N__29841;
    wire N__29838;
    wire N__29837;
    wire N__29836;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29819;
    wire N__29816;
    wire N__29813;
    wire N__29812;
    wire N__29809;
    wire N__29804;
    wire N__29799;
    wire N__29796;
    wire N__29795;
    wire N__29794;
    wire N__29791;
    wire N__29790;
    wire N__29789;
    wire N__29788;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29780;
    wire N__29779;
    wire N__29778;
    wire N__29775;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29759;
    wire N__29756;
    wire N__29755;
    wire N__29754;
    wire N__29753;
    wire N__29752;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29744;
    wire N__29743;
    wire N__29740;
    wire N__29739;
    wire N__29736;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29725;
    wire N__29722;
    wire N__29721;
    wire N__29720;
    wire N__29711;
    wire N__29706;
    wire N__29703;
    wire N__29702;
    wire N__29699;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29691;
    wire N__29690;
    wire N__29689;
    wire N__29686;
    wire N__29685;
    wire N__29684;
    wire N__29683;
    wire N__29682;
    wire N__29681;
    wire N__29680;
    wire N__29679;
    wire N__29678;
    wire N__29677;
    wire N__29676;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29651;
    wire N__29650;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29630;
    wire N__29629;
    wire N__29628;
    wire N__29625;
    wire N__29620;
    wire N__29617;
    wire N__29614;
    wire N__29599;
    wire N__29596;
    wire N__29593;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29577;
    wire N__29574;
    wire N__29573;
    wire N__29570;
    wire N__29569;
    wire N__29566;
    wire N__29559;
    wire N__29556;
    wire N__29551;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29539;
    wire N__29534;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29520;
    wire N__29519;
    wire N__29516;
    wire N__29515;
    wire N__29514;
    wire N__29513;
    wire N__29512;
    wire N__29511;
    wire N__29510;
    wire N__29505;
    wire N__29502;
    wire N__29497;
    wire N__29488;
    wire N__29481;
    wire N__29468;
    wire N__29463;
    wire N__29454;
    wire N__29451;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29402;
    wire N__29399;
    wire N__29392;
    wire N__29385;
    wire N__29378;
    wire N__29375;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29359;
    wire N__29356;
    wire N__29351;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29328;
    wire N__29319;
    wire N__29316;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29237;
    wire N__29236;
    wire N__29235;
    wire N__29234;
    wire N__29233;
    wire N__29232;
    wire N__29231;
    wire N__29228;
    wire N__29227;
    wire N__29226;
    wire N__29225;
    wire N__29220;
    wire N__29213;
    wire N__29212;
    wire N__29209;
    wire N__29202;
    wire N__29197;
    wire N__29196;
    wire N__29195;
    wire N__29194;
    wire N__29189;
    wire N__29188;
    wire N__29185;
    wire N__29182;
    wire N__29177;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29143;
    wire N__29136;
    wire N__29135;
    wire N__29132;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29109;
    wire N__29108;
    wire N__29105;
    wire N__29104;
    wire N__29103;
    wire N__29102;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29085;
    wire N__29082;
    wire N__29081;
    wire N__29078;
    wire N__29073;
    wire N__29070;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29058;
    wire N__29053;
    wire N__29050;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29025;
    wire N__29022;
    wire N__29021;
    wire N__29020;
    wire N__29017;
    wire N__29012;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28980;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28940;
    wire N__28939;
    wire N__28936;
    wire N__28931;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28910;
    wire N__28907;
    wire N__28904;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28887;
    wire N__28886;
    wire N__28883;
    wire N__28882;
    wire N__28879;
    wire N__28876;
    wire N__28871;
    wire N__28866;
    wire N__28863;
    wire N__28860;
    wire N__28857;
    wire N__28854;
    wire N__28851;
    wire N__28848;
    wire N__28845;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28766;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28720;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28702;
    wire N__28699;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28669;
    wire N__28668;
    wire N__28667;
    wire N__28666;
    wire N__28663;
    wire N__28662;
    wire N__28661;
    wire N__28658;
    wire N__28653;
    wire N__28648;
    wire N__28645;
    wire N__28640;
    wire N__28633;
    wire N__28626;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28511;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28494;
    wire N__28493;
    wire N__28492;
    wire N__28489;
    wire N__28484;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28472;
    wire N__28471;
    wire N__28470;
    wire N__28469;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28455;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28438;
    wire N__28435;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28419;
    wire N__28416;
    wire N__28409;
    wire N__28406;
    wire N__28403;
    wire N__28396;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28326;
    wire N__28325;
    wire N__28324;
    wire N__28321;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28303;
    wire N__28302;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28294;
    wire N__28291;
    wire N__28286;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28276;
    wire N__28275;
    wire N__28270;
    wire N__28267;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28249;
    wire N__28246;
    wire N__28245;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28196;
    wire N__28191;
    wire N__28190;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28179;
    wire N__28176;
    wire N__28171;
    wire N__28168;
    wire N__28167;
    wire N__28166;
    wire N__28163;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28148;
    wire N__28145;
    wire N__28142;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28128;
    wire N__28127;
    wire N__28124;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28109;
    wire N__28108;
    wire N__28105;
    wire N__28100;
    wire N__28097;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28057;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28040;
    wire N__28037;
    wire N__28036;
    wire N__28033;
    wire N__28032;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28015;
    wire N__28014;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27991;
    wire N__27984;
    wire N__27981;
    wire N__27980;
    wire N__27979;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27966;
    wire N__27963;
    wire N__27960;
    wire N__27957;
    wire N__27954;
    wire N__27945;
    wire N__27942;
    wire N__27941;
    wire N__27938;
    wire N__27937;
    wire N__27934;
    wire N__27933;
    wire N__27930;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27916;
    wire N__27913;
    wire N__27912;
    wire N__27911;
    wire N__27908;
    wire N__27907;
    wire N__27902;
    wire N__27899;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27882;
    wire N__27879;
    wire N__27874;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27834;
    wire N__27831;
    wire N__27830;
    wire N__27827;
    wire N__27824;
    wire N__27823;
    wire N__27822;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27804;
    wire N__27803;
    wire N__27800;
    wire N__27799;
    wire N__27796;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27781;
    wire N__27776;
    wire N__27773;
    wire N__27772;
    wire N__27767;
    wire N__27764;
    wire N__27763;
    wire N__27758;
    wire N__27755;
    wire N__27750;
    wire N__27747;
    wire N__27742;
    wire N__27737;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27659;
    wire N__27658;
    wire N__27657;
    wire N__27654;
    wire N__27653;
    wire N__27650;
    wire N__27647;
    wire N__27646;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27634;
    wire N__27631;
    wire N__27628;
    wire N__27625;
    wire N__27612;
    wire N__27611;
    wire N__27608;
    wire N__27607;
    wire N__27604;
    wire N__27603;
    wire N__27602;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27584;
    wire N__27573;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27563;
    wire N__27562;
    wire N__27561;
    wire N__27560;
    wire N__27559;
    wire N__27558;
    wire N__27557;
    wire N__27554;
    wire N__27547;
    wire N__27544;
    wire N__27543;
    wire N__27542;
    wire N__27537;
    wire N__27534;
    wire N__27533;
    wire N__27532;
    wire N__27527;
    wire N__27524;
    wire N__27519;
    wire N__27518;
    wire N__27517;
    wire N__27512;
    wire N__27507;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27450;
    wire N__27447;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27380;
    wire N__27379;
    wire N__27378;
    wire N__27375;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27363;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27336;
    wire N__27333;
    wire N__27330;
    wire N__27327;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27303;
    wire N__27300;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27288;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27247;
    wire N__27246;
    wire N__27241;
    wire N__27238;
    wire N__27237;
    wire N__27234;
    wire N__27233;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27218;
    wire N__27213;
    wire N__27208;
    wire N__27205;
    wire N__27204;
    wire N__27201;
    wire N__27196;
    wire N__27193;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27093;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27074;
    wire N__27071;
    wire N__27070;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26975;
    wire N__26974;
    wire N__26973;
    wire N__26972;
    wire N__26971;
    wire N__26968;
    wire N__26967;
    wire N__26964;
    wire N__26963;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26917;
    wire N__26912;
    wire N__26907;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26876;
    wire N__26875;
    wire N__26872;
    wire N__26871;
    wire N__26868;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26820;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26792;
    wire N__26791;
    wire N__26790;
    wire N__26789;
    wire N__26788;
    wire N__26787;
    wire N__26786;
    wire N__26781;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26726;
    wire N__26721;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26565;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26538;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26484;
    wire N__26481;
    wire N__26478;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26459;
    wire N__26458;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26431;
    wire N__26424;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26400;
    wire N__26397;
    wire N__26394;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26337;
    wire N__26334;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26309;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26301;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26289;
    wire N__26286;
    wire N__26283;
    wire N__26274;
    wire N__26273;
    wire N__26272;
    wire N__26271;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26259;
    wire N__26256;
    wire N__26255;
    wire N__26252;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26226;
    wire N__26225;
    wire N__26224;
    wire N__26223;
    wire N__26222;
    wire N__26219;
    wire N__26218;
    wire N__26215;
    wire N__26214;
    wire N__26213;
    wire N__26212;
    wire N__26211;
    wire N__26210;
    wire N__26209;
    wire N__26208;
    wire N__26207;
    wire N__26206;
    wire N__26205;
    wire N__26204;
    wire N__26203;
    wire N__26202;
    wire N__26201;
    wire N__26200;
    wire N__26199;
    wire N__26198;
    wire N__26197;
    wire N__26196;
    wire N__26195;
    wire N__26194;
    wire N__26193;
    wire N__26192;
    wire N__26191;
    wire N__26190;
    wire N__26189;
    wire N__26188;
    wire N__26187;
    wire N__26186;
    wire N__26185;
    wire N__26184;
    wire N__26183;
    wire N__26182;
    wire N__26181;
    wire N__26180;
    wire N__26175;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26161;
    wire N__26156;
    wire N__26153;
    wire N__26148;
    wire N__26143;
    wire N__26140;
    wire N__26137;
    wire N__26134;
    wire N__26131;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26115;
    wire N__26112;
    wire N__26107;
    wire N__26102;
    wire N__26097;
    wire N__26090;
    wire N__26085;
    wire N__26082;
    wire N__26077;
    wire N__26072;
    wire N__26071;
    wire N__26070;
    wire N__26069;
    wire N__26068;
    wire N__26067;
    wire N__26066;
    wire N__26065;
    wire N__26064;
    wire N__26063;
    wire N__26062;
    wire N__26061;
    wire N__26060;
    wire N__26059;
    wire N__26058;
    wire N__26057;
    wire N__26056;
    wire N__26055;
    wire N__26054;
    wire N__26053;
    wire N__26052;
    wire N__26051;
    wire N__26050;
    wire N__26049;
    wire N__26048;
    wire N__26047;
    wire N__26046;
    wire N__26045;
    wire N__26044;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25857;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25721;
    wire N__25720;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25708;
    wire N__25705;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25590;
    wire N__25589;
    wire N__25588;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25436;
    wire N__25435;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25423;
    wire N__25420;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25356;
    wire N__25353;
    wire N__25352;
    wire N__25347;
    wire N__25346;
    wire N__25345;
    wire N__25344;
    wire N__25343;
    wire N__25340;
    wire N__25331;
    wire N__25330;
    wire N__25327;
    wire N__25324;
    wire N__25321;
    wire N__25314;
    wire N__25313;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25302;
    wire N__25301;
    wire N__25300;
    wire N__25291;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25260;
    wire N__25257;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25200;
    wire N__25197;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25168;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25156;
    wire N__25153;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25033;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24889;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24745;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24708;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24623;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24609;
    wire N__24608;
    wire N__24605;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24585;
    wire N__24584;
    wire N__24581;
    wire N__24580;
    wire N__24577;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24562;
    wire N__24557;
    wire N__24554;
    wire N__24553;
    wire N__24548;
    wire N__24545;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24530;
    wire N__24527;
    wire N__24520;
    wire N__24515;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24503;
    wire N__24502;
    wire N__24499;
    wire N__24498;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24490;
    wire N__24489;
    wire N__24488;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24474;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24463;
    wire N__24462;
    wire N__24459;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24445;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24381;
    wire N__24372;
    wire N__24367;
    wire N__24364;
    wire N__24359;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24317;
    wire N__24314;
    wire N__24313;
    wire N__24310;
    wire N__24309;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24301;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24285;
    wire N__24282;
    wire N__24281;
    wire N__24278;
    wire N__24275;
    wire N__24268;
    wire N__24265;
    wire N__24260;
    wire N__24257;
    wire N__24252;
    wire N__24243;
    wire N__24242;
    wire N__24241;
    wire N__24240;
    wire N__24239;
    wire N__24236;
    wire N__24235;
    wire N__24232;
    wire N__24231;
    wire N__24228;
    wire N__24227;
    wire N__24226;
    wire N__24225;
    wire N__24224;
    wire N__24223;
    wire N__24222;
    wire N__24221;
    wire N__24218;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24192;
    wire N__24187;
    wire N__24180;
    wire N__24179;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24165;
    wire N__24164;
    wire N__24163;
    wire N__24162;
    wire N__24161;
    wire N__24160;
    wire N__24159;
    wire N__24158;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24144;
    wire N__24141;
    wire N__24136;
    wire N__24131;
    wire N__24130;
    wire N__24129;
    wire N__24128;
    wire N__24127;
    wire N__24126;
    wire N__24125;
    wire N__24118;
    wire N__24115;
    wire N__24110;
    wire N__24107;
    wire N__24098;
    wire N__24093;
    wire N__24084;
    wire N__24077;
    wire N__24070;
    wire N__24051;
    wire N__24048;
    wire N__24047;
    wire N__24046;
    wire N__24045;
    wire N__24044;
    wire N__24043;
    wire N__24042;
    wire N__24041;
    wire N__24040;
    wire N__24039;
    wire N__24038;
    wire N__24029;
    wire N__24020;
    wire N__24019;
    wire N__24016;
    wire N__24011;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23999;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23958;
    wire N__23957;
    wire N__23956;
    wire N__23955;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23947;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23922;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23906;
    wire N__23905;
    wire N__23902;
    wire N__23901;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23889;
    wire N__23886;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23841;
    wire N__23838;
    wire N__23835;
    wire N__23832;
    wire N__23829;
    wire N__23828;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23820;
    wire N__23817;
    wire N__23812;
    wire N__23809;
    wire N__23802;
    wire N__23799;
    wire N__23798;
    wire N__23797;
    wire N__23796;
    wire N__23795;
    wire N__23792;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23781;
    wire N__23780;
    wire N__23777;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23762;
    wire N__23757;
    wire N__23752;
    wire N__23745;
    wire N__23740;
    wire N__23733;
    wire N__23732;
    wire N__23731;
    wire N__23728;
    wire N__23727;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23703;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23656;
    wire N__23653;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23576;
    wire N__23573;
    wire N__23572;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23542;
    wire N__23539;
    wire N__23532;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23519;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23495;
    wire N__23492;
    wire N__23491;
    wire N__23490;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23478;
    wire N__23475;
    wire N__23474;
    wire N__23473;
    wire N__23472;
    wire N__23469;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23447;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23429;
    wire N__23428;
    wire N__23425;
    wire N__23420;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23408;
    wire N__23407;
    wire N__23406;
    wire N__23403;
    wire N__23402;
    wire N__23401;
    wire N__23398;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23360;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23326;
    wire N__23319;
    wire N__23318;
    wire N__23317;
    wire N__23316;
    wire N__23315;
    wire N__23314;
    wire N__23313;
    wire N__23312;
    wire N__23311;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23285;
    wire N__23284;
    wire N__23283;
    wire N__23282;
    wire N__23279;
    wire N__23278;
    wire N__23277;
    wire N__23276;
    wire N__23273;
    wire N__23272;
    wire N__23269;
    wire N__23268;
    wire N__23267;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23259;
    wire N__23254;
    wire N__23251;
    wire N__23250;
    wire N__23249;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23237;
    wire N__23234;
    wire N__23229;
    wire N__23222;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23214;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23203;
    wire N__23202;
    wire N__23201;
    wire N__23200;
    wire N__23199;
    wire N__23194;
    wire N__23191;
    wire N__23184;
    wire N__23183;
    wire N__23180;
    wire N__23175;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23159;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23147;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23127;
    wire N__23120;
    wire N__23115;
    wire N__23100;
    wire N__23099;
    wire N__23098;
    wire N__23097;
    wire N__23094;
    wire N__23093;
    wire N__23092;
    wire N__23091;
    wire N__23090;
    wire N__23089;
    wire N__23088;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23077;
    wire N__23074;
    wire N__23073;
    wire N__23070;
    wire N__23069;
    wire N__23066;
    wire N__23065;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23040;
    wire N__23039;
    wire N__23036;
    wire N__23031;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23004;
    wire N__23001;
    wire N__23000;
    wire N__22999;
    wire N__22998;
    wire N__22997;
    wire N__22996;
    wire N__22995;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22983;
    wire N__22980;
    wire N__22971;
    wire N__22966;
    wire N__22957;
    wire N__22952;
    wire N__22935;
    wire N__22934;
    wire N__22933;
    wire N__22930;
    wire N__22929;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22915;
    wire N__22912;
    wire N__22907;
    wire N__22902;
    wire N__22899;
    wire N__22898;
    wire N__22895;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22869;
    wire N__22868;
    wire N__22867;
    wire N__22866;
    wire N__22865;
    wire N__22862;
    wire N__22861;
    wire N__22860;
    wire N__22859;
    wire N__22858;
    wire N__22857;
    wire N__22856;
    wire N__22855;
    wire N__22854;
    wire N__22851;
    wire N__22850;
    wire N__22849;
    wire N__22844;
    wire N__22843;
    wire N__22842;
    wire N__22841;
    wire N__22840;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22816;
    wire N__22813;
    wire N__22808;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22783;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22771;
    wire N__22760;
    wire N__22755;
    wire N__22750;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22725;
    wire N__22716;
    wire N__22715;
    wire N__22714;
    wire N__22713;
    wire N__22710;
    wire N__22709;
    wire N__22708;
    wire N__22707;
    wire N__22706;
    wire N__22705;
    wire N__22704;
    wire N__22703;
    wire N__22702;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22677;
    wire N__22674;
    wire N__22673;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22659;
    wire N__22656;
    wire N__22649;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22613;
    wire N__22610;
    wire N__22605;
    wire N__22600;
    wire N__22593;
    wire N__22584;
    wire N__22583;
    wire N__22582;
    wire N__22581;
    wire N__22580;
    wire N__22579;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22571;
    wire N__22570;
    wire N__22569;
    wire N__22566;
    wire N__22559;
    wire N__22556;
    wire N__22551;
    wire N__22546;
    wire N__22545;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22537;
    wire N__22536;
    wire N__22535;
    wire N__22534;
    wire N__22533;
    wire N__22532;
    wire N__22531;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22503;
    wire N__22502;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22482;
    wire N__22471;
    wire N__22464;
    wire N__22459;
    wire N__22452;
    wire N__22437;
    wire N__22434;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22403;
    wire N__22402;
    wire N__22401;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22393;
    wire N__22392;
    wire N__22391;
    wire N__22388;
    wire N__22387;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22367;
    wire N__22364;
    wire N__22363;
    wire N__22362;
    wire N__22361;
    wire N__22360;
    wire N__22357;
    wire N__22356;
    wire N__22353;
    wire N__22352;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22335;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22320;
    wire N__22317;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22305;
    wire N__22296;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22272;
    wire N__22271;
    wire N__22270;
    wire N__22269;
    wire N__22266;
    wire N__22265;
    wire N__22264;
    wire N__22257;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22237;
    wire N__22228;
    wire N__22225;
    wire N__22220;
    wire N__22213;
    wire N__22200;
    wire N__22197;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22171;
    wire N__22168;
    wire N__22167;
    wire N__22164;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22137;
    wire N__22134;
    wire N__22133;
    wire N__22130;
    wire N__22129;
    wire N__22126;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22097;
    wire N__22094;
    wire N__22093;
    wire N__22092;
    wire N__22087;
    wire N__22084;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22068;
    wire N__22063;
    wire N__22060;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22031;
    wire N__22030;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__22001;
    wire N__22000;
    wire N__21999;
    wire N__21994;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21986;
    wire N__21985;
    wire N__21982;
    wire N__21979;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21967;
    wire N__21964;
    wire N__21963;
    wire N__21962;
    wire N__21957;
    wire N__21952;
    wire N__21951;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21947;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21935;
    wire N__21930;
    wire N__21923;
    wire N__21916;
    wire N__21903;
    wire N__21902;
    wire N__21901;
    wire N__21898;
    wire N__21897;
    wire N__21894;
    wire N__21893;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21882;
    wire N__21879;
    wire N__21874;
    wire N__21873;
    wire N__21872;
    wire N__21871;
    wire N__21868;
    wire N__21863;
    wire N__21862;
    wire N__21861;
    wire N__21860;
    wire N__21857;
    wire N__21852;
    wire N__21847;
    wire N__21844;
    wire N__21839;
    wire N__21832;
    wire N__21819;
    wire N__21818;
    wire N__21815;
    wire N__21814;
    wire N__21813;
    wire N__21812;
    wire N__21811;
    wire N__21810;
    wire N__21807;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21795;
    wire N__21786;
    wire N__21777;
    wire N__21776;
    wire N__21775;
    wire N__21774;
    wire N__21771;
    wire N__21770;
    wire N__21769;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21751;
    wire N__21748;
    wire N__21735;
    wire N__21734;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21719;
    wire N__21716;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21698;
    wire N__21693;
    wire N__21692;
    wire N__21691;
    wire N__21690;
    wire N__21687;
    wire N__21680;
    wire N__21675;
    wire N__21674;
    wire N__21671;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21663;
    wire N__21662;
    wire N__21661;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21643;
    wire N__21640;
    wire N__21639;
    wire N__21638;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21623;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21579;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21539;
    wire N__21538;
    wire N__21537;
    wire N__21536;
    wire N__21531;
    wire N__21526;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21501;
    wire N__21498;
    wire N__21497;
    wire N__21496;
    wire N__21495;
    wire N__21494;
    wire N__21493;
    wire N__21492;
    wire N__21491;
    wire N__21490;
    wire N__21489;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21478;
    wire N__21477;
    wire N__21476;
    wire N__21473;
    wire N__21466;
    wire N__21461;
    wire N__21458;
    wire N__21449;
    wire N__21442;
    wire N__21435;
    wire N__21432;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21402;
    wire N__21393;
    wire N__21390;
    wire N__21389;
    wire N__21386;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21357;
    wire N__21354;
    wire N__21353;
    wire N__21352;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21323;
    wire N__21322;
    wire N__21321;
    wire N__21320;
    wire N__21319;
    wire N__21318;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21299;
    wire N__21292;
    wire N__21289;
    wire N__21284;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21272;
    wire N__21267;
    wire N__21264;
    wire N__21263;
    wire N__21262;
    wire N__21259;
    wire N__21254;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21161;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21101;
    wire N__21100;
    wire N__21099;
    wire N__21094;
    wire N__21093;
    wire N__21090;
    wire N__21089;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21057;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21026;
    wire N__21025;
    wire N__21020;
    wire N__21017;
    wire N__21012;
    wire N__21011;
    wire N__21010;
    wire N__21009;
    wire N__21004;
    wire N__20999;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20978;
    wire N__20977;
    wire N__20976;
    wire N__20971;
    wire N__20966;
    wire N__20961;
    wire N__20958;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20926;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20913;
    wire N__20912;
    wire N__20911;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20894;
    wire N__20891;
    wire N__20886;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20731;
    wire N__20730;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20716;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20670;
    wire N__20667;
    wire N__20666;
    wire N__20663;
    wire N__20662;
    wire N__20661;
    wire N__20660;
    wire N__20657;
    wire N__20656;
    wire N__20655;
    wire N__20654;
    wire N__20653;
    wire N__20652;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20640;
    wire N__20637;
    wire N__20632;
    wire N__20623;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20572;
    wire N__20571;
    wire N__20570;
    wire N__20569;
    wire N__20566;
    wire N__20565;
    wire N__20560;
    wire N__20553;
    wire N__20552;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20520;
    wire N__20519;
    wire N__20518;
    wire N__20515;
    wire N__20514;
    wire N__20513;
    wire N__20510;
    wire N__20509;
    wire N__20508;
    wire N__20505;
    wire N__20504;
    wire N__20503;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20478;
    wire N__20475;
    wire N__20466;
    wire N__20457;
    wire N__20456;
    wire N__20455;
    wire N__20454;
    wire N__20451;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20439;
    wire N__20436;
    wire N__20431;
    wire N__20424;
    wire N__20423;
    wire N__20420;
    wire N__20419;
    wire N__20418;
    wire N__20415;
    wire N__20414;
    wire N__20413;
    wire N__20412;
    wire N__20411;
    wire N__20410;
    wire N__20409;
    wire N__20406;
    wire N__20401;
    wire N__20398;
    wire N__20393;
    wire N__20384;
    wire N__20373;
    wire N__20372;
    wire N__20371;
    wire N__20370;
    wire N__20367;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20355;
    wire N__20352;
    wire N__20351;
    wire N__20348;
    wire N__20343;
    wire N__20342;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20334;
    wire N__20333;
    wire N__20328;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20312;
    wire N__20301;
    wire N__20298;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20248;
    wire N__20247;
    wire N__20246;
    wire N__20245;
    wire N__20240;
    wire N__20239;
    wire N__20238;
    wire N__20237;
    wire N__20234;
    wire N__20233;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20205;
    wire N__20202;
    wire N__20187;
    wire N__20184;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20130;
    wire N__20127;
    wire N__20126;
    wire N__20125;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20113;
    wire N__20110;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20087;
    wire N__20086;
    wire N__20085;
    wire N__20084;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20073;
    wire N__20072;
    wire N__20071;
    wire N__20070;
    wire N__20067;
    wire N__20064;
    wire N__20059;
    wire N__20056;
    wire N__20049;
    wire N__20044;
    wire N__20041;
    wire N__20028;
    wire N__20027;
    wire N__20026;
    wire N__20025;
    wire N__20022;
    wire N__20015;
    wire N__20012;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19934;
    wire N__19933;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19921;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19898;
    wire N__19897;
    wire N__19896;
    wire N__19893;
    wire N__19892;
    wire N__19891;
    wire N__19888;
    wire N__19887;
    wire N__19884;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19876;
    wire N__19873;
    wire N__19872;
    wire N__19869;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19824;
    wire N__19823;
    wire N__19818;
    wire N__19813;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19795;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19777;
    wire N__19774;
    wire N__19767;
    wire N__19764;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19756;
    wire N__19755;
    wire N__19754;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19731;
    wire N__19728;
    wire N__19727;
    wire N__19724;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19707;
    wire N__19706;
    wire N__19705;
    wire N__19704;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19696;
    wire N__19693;
    wire N__19688;
    wire N__19687;
    wire N__19686;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19667;
    wire N__19662;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19629;
    wire N__19628;
    wire N__19627;
    wire N__19626;
    wire N__19625;
    wire N__19624;
    wire N__19621;
    wire N__19620;
    wire N__19619;
    wire N__19616;
    wire N__19611;
    wire N__19606;
    wire N__19603;
    wire N__19598;
    wire N__19593;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19572;
    wire N__19569;
    wire N__19568;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19560;
    wire N__19559;
    wire N__19556;
    wire N__19551;
    wire N__19550;
    wire N__19549;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19491;
    wire N__19490;
    wire N__19489;
    wire N__19488;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19457;
    wire N__19456;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19444;
    wire N__19437;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19427;
    wire N__19424;
    wire N__19423;
    wire N__19422;
    wire N__19419;
    wire N__19416;
    wire N__19411;
    wire N__19404;
    wire N__19403;
    wire N__19400;
    wire N__19399;
    wire N__19396;
    wire N__19395;
    wire N__19394;
    wire N__19391;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19364;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19311;
    wire N__19308;
    wire N__19307;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19290;
    wire N__19287;
    wire N__19286;
    wire N__19285;
    wire N__19282;
    wire N__19275;
    wire N__19266;
    wire N__19263;
    wire N__19258;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19146;
    wire N__19145;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19126;
    wire N__19119;
    wire N__19116;
    wire N__19115;
    wire N__19112;
    wire N__19111;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19099;
    wire N__19092;
    wire N__19091;
    wire N__19088;
    wire N__19087;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19075;
    wire N__19068;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19058;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__19004;
    wire N__19001;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18966;
    wire N__18963;
    wire N__18962;
    wire N__18961;
    wire N__18954;
    wire N__18953;
    wire N__18952;
    wire N__18951;
    wire N__18948;
    wire N__18941;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18884;
    wire N__18883;
    wire N__18882;
    wire N__18879;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18862;
    wire N__18855;
    wire N__18854;
    wire N__18851;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18839;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18818;
    wire N__18817;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18798;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18786;
    wire N__18785;
    wire N__18784;
    wire N__18783;
    wire N__18782;
    wire N__18781;
    wire N__18778;
    wire N__18777;
    wire N__18776;
    wire N__18773;
    wire N__18772;
    wire N__18769;
    wire N__18768;
    wire N__18767;
    wire N__18766;
    wire N__18765;
    wire N__18764;
    wire N__18763;
    wire N__18762;
    wire N__18755;
    wire N__18752;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18738;
    wire N__18731;
    wire N__18726;
    wire N__18721;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18674;
    wire N__18673;
    wire N__18670;
    wire N__18665;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18623;
    wire N__18622;
    wire N__18621;
    wire N__18620;
    wire N__18619;
    wire N__18618;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18610;
    wire N__18609;
    wire N__18608;
    wire N__18605;
    wire N__18602;
    wire N__18601;
    wire N__18600;
    wire N__18599;
    wire N__18598;
    wire N__18597;
    wire N__18596;
    wire N__18593;
    wire N__18592;
    wire N__18591;
    wire N__18590;
    wire N__18589;
    wire N__18588;
    wire N__18587;
    wire N__18586;
    wire N__18585;
    wire N__18584;
    wire N__18583;
    wire N__18582;
    wire N__18581;
    wire N__18580;
    wire N__18579;
    wire N__18578;
    wire N__18577;
    wire N__18576;
    wire N__18575;
    wire N__18572;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18554;
    wire N__18549;
    wire N__18536;
    wire N__18533;
    wire N__18528;
    wire N__18527;
    wire N__18518;
    wire N__18509;
    wire N__18496;
    wire N__18491;
    wire N__18484;
    wire N__18483;
    wire N__18482;
    wire N__18477;
    wire N__18472;
    wire N__18467;
    wire N__18464;
    wire N__18457;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18429;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18408;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18369;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18297;
    wire N__18294;
    wire N__18293;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18260;
    wire N__18259;
    wire N__18258;
    wire N__18257;
    wire N__18252;
    wire N__18251;
    wire N__18250;
    wire N__18249;
    wire N__18248;
    wire N__18247;
    wire N__18244;
    wire N__18243;
    wire N__18242;
    wire N__18237;
    wire N__18236;
    wire N__18235;
    wire N__18234;
    wire N__18233;
    wire N__18232;
    wire N__18231;
    wire N__18230;
    wire N__18229;
    wire N__18226;
    wire N__18215;
    wire N__18212;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18194;
    wire N__18185;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18084;
    wire N__18081;
    wire N__18080;
    wire N__18079;
    wire N__18078;
    wire N__18075;
    wire N__18068;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18012;
    wire N__18009;
    wire N__18008;
    wire N__18007;
    wire N__18004;
    wire N__18003;
    wire N__18000;
    wire N__17995;
    wire N__17992;
    wire N__17985;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17975;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17958;
    wire N__17957;
    wire N__17954;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17944;
    wire N__17939;
    wire N__17934;
    wire N__17933;
    wire N__17930;
    wire N__17929;
    wire N__17928;
    wire N__17925;
    wire N__17920;
    wire N__17917;
    wire N__17910;
    wire N__17907;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17895;
    wire N__17892;
    wire N__17889;
    wire N__17886;
    wire N__17885;
    wire N__17884;
    wire N__17877;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17826;
    wire N__17823;
    wire N__17820;
    wire N__17817;
    wire N__17814;
    wire N__17811;
    wire N__17808;
    wire N__17805;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17784;
    wire N__17781;
    wire N__17778;
    wire N__17775;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17736;
    wire N__17735;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17725;
    wire N__17724;
    wire N__17721;
    wire N__17718;
    wire N__17715;
    wire N__17712;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17693;
    wire N__17688;
    wire N__17685;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17663;
    wire N__17660;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17649;
    wire N__17646;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17625;
    wire N__17622;
    wire N__17617;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17601;
    wire N__17598;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17574;
    wire N__17571;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17556;
    wire N__17553;
    wire N__17550;
    wire N__17547;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17535;
    wire N__17532;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17520;
    wire N__17517;
    wire N__17514;
    wire N__17511;
    wire N__17508;
    wire N__17505;
    wire N__17502;
    wire N__17499;
    wire N__17496;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17468;
    wire N__17467;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17439;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17409;
    wire N__17406;
    wire N__17403;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17391;
    wire N__17388;
    wire N__17385;
    wire N__17382;
    wire N__17379;
    wire N__17376;
    wire N__17373;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17357;
    wire N__17354;
    wire N__17353;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17339;
    wire N__17336;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17304;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17280;
    wire N__17277;
    wire N__17274;
    wire N__17271;
    wire N__17268;
    wire N__17265;
    wire N__17262;
    wire N__17259;
    wire N__17256;
    wire N__17253;
    wire N__17250;
    wire N__17247;
    wire N__17244;
    wire N__17241;
    wire N__17238;
    wire N__17235;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17217;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17196;
    wire N__17193;
    wire N__17190;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17145;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17130;
    wire N__17129;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17121;
    wire N__17120;
    wire N__17119;
    wire N__17118;
    wire N__17115;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17103;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17079;
    wire N__17078;
    wire N__17071;
    wire N__17068;
    wire N__17063;
    wire N__17058;
    wire N__17049;
    wire N__17046;
    wire N__17043;
    wire N__17040;
    wire N__17037;
    wire N__17034;
    wire N__17031;
    wire N__17028;
    wire N__17025;
    wire N__17022;
    wire N__17019;
    wire N__17016;
    wire N__17013;
    wire N__17010;
    wire N__17007;
    wire N__17004;
    wire N__17001;
    wire N__16998;
    wire N__16995;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16982;
    wire N__16979;
    wire N__16978;
    wire N__16975;
    wire N__16974;
    wire N__16973;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16956;
    wire N__16947;
    wire N__16946;
    wire N__16945;
    wire N__16944;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16930;
    wire N__16923;
    wire N__16922;
    wire N__16921;
    wire N__16918;
    wire N__16917;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16887;
    wire N__16886;
    wire N__16885;
    wire N__16882;
    wire N__16877;
    wire N__16876;
    wire N__16873;
    wire N__16872;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16857;
    wire N__16848;
    wire N__16845;
    wire N__16842;
    wire N__16839;
    wire N__16836;
    wire N__16835;
    wire N__16834;
    wire N__16833;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16825;
    wire N__16822;
    wire N__16821;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16804;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16782;
    wire N__16779;
    wire N__16776;
    wire N__16775;
    wire N__16772;
    wire N__16771;
    wire N__16768;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16755;
    wire N__16752;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16731;
    wire N__16722;
    wire N__16721;
    wire N__16720;
    wire N__16713;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16691;
    wire N__16688;
    wire N__16687;
    wire N__16686;
    wire N__16683;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16656;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16638;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16626;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16615;
    wire N__16614;
    wire N__16611;
    wire N__16610;
    wire N__16607;
    wire N__16602;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16584;
    wire N__16583;
    wire N__16582;
    wire N__16579;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16567;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16555;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16520;
    wire N__16517;
    wire N__16516;
    wire N__16513;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16503;
    wire N__16500;
    wire N__16499;
    wire N__16494;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16470;
    wire N__16467;
    wire N__16464;
    wire N__16461;
    wire N__16458;
    wire N__16455;
    wire N__16452;
    wire N__16449;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16437;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16425;
    wire N__16422;
    wire N__16419;
    wire N__16416;
    wire N__16413;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16319;
    wire N__16318;
    wire N__16317;
    wire N__16316;
    wire N__16305;
    wire N__16304;
    wire N__16303;
    wire N__16302;
    wire N__16299;
    wire N__16294;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16280;
    wire N__16277;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16227;
    wire N__16224;
    wire N__16221;
    wire N__16218;
    wire N__16215;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16205;
    wire N__16202;
    wire N__16199;
    wire N__16198;
    wire N__16197;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16176;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16163;
    wire N__16158;
    wire N__16157;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16137;
    wire N__16136;
    wire N__16135;
    wire N__16132;
    wire N__16131;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16123;
    wire N__16122;
    wire N__16121;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16113;
    wire N__16112;
    wire N__16109;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16091;
    wire N__16086;
    wire N__16083;
    wire N__16080;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16064;
    wire N__16061;
    wire N__16056;
    wire N__16053;
    wire N__16050;
    wire N__16049;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16037;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16021;
    wire N__16016;
    wire N__16015;
    wire N__16012;
    wire N__16011;
    wire N__16008;
    wire N__16005;
    wire N__16002;
    wire N__15999;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15985;
    wire N__15982;
    wire N__15977;
    wire N__15972;
    wire N__15965;
    wire N__15962;
    wire N__15957;
    wire N__15954;
    wire N__15951;
    wire N__15948;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15936;
    wire N__15933;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15921;
    wire N__15918;
    wire N__15915;
    wire N__15912;
    wire N__15909;
    wire N__15906;
    wire N__15903;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15882;
    wire N__15879;
    wire N__15876;
    wire N__15873;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15851;
    wire N__15850;
    wire N__15847;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15835;
    wire N__15832;
    wire N__15829;
    wire N__15822;
    wire N__15821;
    wire N__15818;
    wire N__15817;
    wire N__15816;
    wire N__15815;
    wire N__15814;
    wire N__15811;
    wire N__15810;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15790;
    wire N__15787;
    wire N__15782;
    wire N__15779;
    wire N__15774;
    wire N__15773;
    wire N__15772;
    wire N__15771;
    wire N__15768;
    wire N__15765;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15736;
    wire N__15733;
    wire N__15726;
    wire N__15723;
    wire N__15720;
    wire N__15717;
    wire N__15714;
    wire N__15711;
    wire N__15708;
    wire N__15705;
    wire N__15702;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15657;
    wire N__15654;
    wire N__15651;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15597;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15573;
    wire N__15570;
    wire N__15567;
    wire N__15564;
    wire N__15561;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15489;
    wire N__15486;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15462;
    wire N__15459;
    wire N__15456;
    wire N__15453;
    wire N__15452;
    wire N__15447;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15420;
    wire N__15417;
    wire N__15414;
    wire N__15411;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15399;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15374;
    wire N__15373;
    wire N__15370;
    wire N__15367;
    wire N__15364;
    wire N__15357;
    wire N__15356;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15327;
    wire N__15326;
    wire N__15325;
    wire N__15322;
    wire N__15317;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15249;
    wire N__15246;
    wire N__15243;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15213;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15198;
    wire N__15195;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15173;
    wire N__15172;
    wire N__15171;
    wire N__15166;
    wire N__15165;
    wire N__15162;
    wire N__15161;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15144;
    wire N__15141;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15119;
    wire N__15118;
    wire N__15117;
    wire N__15116;
    wire N__15115;
    wire N__15112;
    wire N__15107;
    wire N__15104;
    wire N__15099;
    wire N__15096;
    wire N__15087;
    wire N__15086;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15053;
    wire N__15052;
    wire N__15051;
    wire N__15046;
    wire N__15041;
    wire N__15036;
    wire N__15033;
    wire N__15032;
    wire N__15031;
    wire N__15030;
    wire N__15027;
    wire N__15024;
    wire N__15019;
    wire N__15012;
    wire N__15009;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14985;
    wire N__14982;
    wire N__14979;
    wire N__14976;
    wire N__14973;
    wire N__14972;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14962;
    wire N__14955;
    wire N__14952;
    wire N__14951;
    wire N__14950;
    wire N__14947;
    wire N__14942;
    wire N__14937;
    wire N__14936;
    wire N__14935;
    wire N__14932;
    wire N__14927;
    wire N__14922;
    wire N__14919;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14901;
    wire N__14898;
    wire N__14895;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14849;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14838;
    wire N__14837;
    wire N__14834;
    wire N__14829;
    wire N__14828;
    wire N__14823;
    wire N__14818;
    wire N__14815;
    wire N__14808;
    wire N__14807;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14799;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14789;
    wire N__14784;
    wire N__14783;
    wire N__14776;
    wire N__14773;
    wire N__14772;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14760;
    wire N__14751;
    wire N__14750;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14682;
    wire N__14679;
    wire N__14676;
    wire N__14673;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14661;
    wire N__14658;
    wire N__14657;
    wire N__14652;
    wire N__14649;
    wire N__14648;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14640;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14622;
    wire N__14619;
    wire N__14618;
    wire N__14617;
    wire N__14614;
    wire N__14613;
    wire N__14612;
    wire N__14611;
    wire N__14608;
    wire N__14607;
    wire N__14604;
    wire N__14601;
    wire N__14600;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14579;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14553;
    wire N__14552;
    wire N__14551;
    wire N__14550;
    wire N__14549;
    wire N__14548;
    wire N__14547;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14535;
    wire N__14532;
    wire N__14529;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14521;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14481;
    wire N__14480;
    wire N__14479;
    wire N__14478;
    wire N__14477;
    wire N__14476;
    wire N__14475;
    wire N__14474;
    wire N__14473;
    wire N__14472;
    wire N__14463;
    wire N__14458;
    wire N__14455;
    wire N__14454;
    wire N__14451;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14437;
    wire N__14434;
    wire N__14421;
    wire N__14420;
    wire N__14419;
    wire N__14418;
    wire N__14413;
    wire N__14412;
    wire N__14411;
    wire N__14410;
    wire N__14407;
    wire N__14406;
    wire N__14403;
    wire N__14402;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14387;
    wire N__14378;
    wire N__14367;
    wire N__14364;
    wire N__14363;
    wire N__14360;
    wire N__14359;
    wire N__14356;
    wire N__14353;
    wire N__14352;
    wire N__14351;
    wire N__14350;
    wire N__14349;
    wire N__14348;
    wire N__14347;
    wire N__14346;
    wire N__14343;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14321;
    wire N__14310;
    wire N__14309;
    wire N__14306;
    wire N__14305;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14292;
    wire N__14291;
    wire N__14290;
    wire N__14287;
    wire N__14282;
    wire N__14279;
    wire N__14278;
    wire N__14275;
    wire N__14274;
    wire N__14271;
    wire N__14264;
    wire N__14261;
    wire N__14256;
    wire N__14247;
    wire N__14246;
    wire N__14245;
    wire N__14242;
    wire N__14237;
    wire N__14236;
    wire N__14235;
    wire N__14230;
    wire N__14227;
    wire N__14226;
    wire N__14225;
    wire N__14224;
    wire N__14221;
    wire N__14216;
    wire N__14213;
    wire N__14208;
    wire N__14199;
    wire N__14196;
    wire N__14193;
    wire N__14192;
    wire N__14191;
    wire N__14188;
    wire N__14183;
    wire N__14182;
    wire N__14181;
    wire N__14180;
    wire N__14175;
    wire N__14172;
    wire N__14171;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14159;
    wire N__14156;
    wire N__14151;
    wire N__14142;
    wire N__14139;
    wire N__14136;
    wire N__14133;
    wire N__14130;
    wire N__14127;
    wire N__14124;
    wire N__14121;
    wire N__14118;
    wire N__14115;
    wire N__14112;
    wire N__14109;
    wire N__14106;
    wire N__14103;
    wire N__14100;
    wire N__14097;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14052;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14040;
    wire N__14037;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__14010;
    wire N__14007;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13997;
    wire N__13996;
    wire N__13995;
    wire N__13992;
    wire N__13987;
    wire N__13984;
    wire N__13977;
    wire N__13976;
    wire N__13975;
    wire N__13972;
    wire N__13967;
    wire N__13962;
    wire N__13959;
    wire N__13956;
    wire N__13953;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13929;
    wire N__13928;
    wire N__13927;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13901;
    wire N__13890;
    wire N__13887;
    wire N__13884;
    wire N__13881;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13873;
    wire N__13870;
    wire N__13867;
    wire N__13866;
    wire N__13865;
    wire N__13864;
    wire N__13863;
    wire N__13860;
    wire N__13855;
    wire N__13850;
    wire N__13845;
    wire N__13840;
    wire N__13833;
    wire N__13830;
    wire N__13827;
    wire N__13824;
    wire N__13821;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13797;
    wire N__13796;
    wire N__13793;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13779;
    wire N__13776;
    wire N__13773;
    wire N__13768;
    wire N__13765;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13746;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13734;
    wire N__13733;
    wire N__13732;
    wire N__13729;
    wire N__13728;
    wire N__13725;
    wire N__13722;
    wire N__13717;
    wire N__13710;
    wire N__13709;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13697;
    wire N__13692;
    wire N__13689;
    wire N__13686;
    wire N__13683;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13671;
    wire N__13668;
    wire N__13665;
    wire N__13662;
    wire N__13659;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13644;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13608;
    wire N__13607;
    wire N__13606;
    wire N__13605;
    wire N__13604;
    wire N__13601;
    wire N__13596;
    wire N__13591;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13577;
    wire N__13576;
    wire N__13573;
    wire N__13570;
    wire N__13567;
    wire N__13564;
    wire N__13561;
    wire N__13560;
    wire N__13559;
    wire N__13558;
    wire N__13555;
    wire N__13550;
    wire N__13545;
    wire N__13542;
    wire N__13537;
    wire N__13530;
    wire N__13527;
    wire N__13526;
    wire N__13523;
    wire N__13520;
    wire N__13515;
    wire N__13512;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13494;
    wire N__13491;
    wire N__13488;
    wire N__13485;
    wire N__13482;
    wire N__13479;
    wire N__13476;
    wire N__13473;
    wire N__13470;
    wire N__13467;
    wire N__13464;
    wire N__13461;
    wire N__13458;
    wire N__13457;
    wire N__13452;
    wire N__13449;
    wire N__13446;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13434;
    wire N__13431;
    wire N__13428;
    wire N__13425;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13410;
    wire N__13407;
    wire N__13404;
    wire N__13401;
    wire N__13398;
    wire N__13395;
    wire N__13394;
    wire N__13391;
    wire N__13390;
    wire N__13387;
    wire N__13386;
    wire N__13383;
    wire N__13380;
    wire N__13375;
    wire N__13368;
    wire N__13365;
    wire N__13364;
    wire N__13363;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13351;
    wire N__13344;
    wire N__13341;
    wire N__13338;
    wire N__13335;
    wire N__13332;
    wire N__13329;
    wire N__13326;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13305;
    wire N__13302;
    wire N__13299;
    wire N__13296;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13277;
    wire N__13276;
    wire N__13275;
    wire N__13272;
    wire N__13265;
    wire N__13260;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13248;
    wire N__13245;
    wire N__13242;
    wire N__13241;
    wire N__13236;
    wire N__13233;
    wire N__13230;
    wire N__13227;
    wire N__13224;
    wire N__13221;
    wire N__13218;
    wire N__13215;
    wire N__13212;
    wire N__13209;
    wire N__13206;
    wire N__13203;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13165;
    wire N__13162;
    wire N__13157;
    wire N__13152;
    wire N__13149;
    wire N__13146;
    wire N__13143;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13131;
    wire N__13128;
    wire N__13125;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13113;
    wire N__13112;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13094;
    wire N__13091;
    wire N__13088;
    wire N__13083;
    wire N__13082;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13068;
    wire N__13065;
    wire N__13064;
    wire N__13063;
    wire N__13056;
    wire N__13053;
    wire N__13050;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13042;
    wire N__13041;
    wire N__13040;
    wire N__13039;
    wire N__13038;
    wire N__13035;
    wire N__13032;
    wire N__13023;
    wire N__13020;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__12999;
    wire N__12998;
    wire N__12997;
    wire N__12994;
    wire N__12991;
    wire N__12988;
    wire N__12981;
    wire N__12978;
    wire N__12975;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12963;
    wire N__12960;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12948;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12927;
    wire N__12924;
    wire N__12921;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12813;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12714;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12695;
    wire N__12692;
    wire N__12689;
    wire N__12684;
    wire N__12681;
    wire N__12680;
    wire N__12679;
    wire N__12676;
    wire N__12671;
    wire N__12670;
    wire N__12669;
    wire N__12668;
    wire N__12663;
    wire N__12660;
    wire N__12655;
    wire N__12648;
    wire N__12645;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12602;
    wire N__12601;
    wire N__12594;
    wire N__12593;
    wire N__12592;
    wire N__12589;
    wire N__12584;
    wire N__12583;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12558;
    wire N__12557;
    wire N__12556;
    wire N__12553;
    wire N__12552;
    wire N__12551;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12537;
    wire N__12532;
    wire N__12529;
    wire N__12526;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12507;
    wire N__12506;
    wire N__12505;
    wire N__12502;
    wire N__12501;
    wire N__12498;
    wire N__12497;
    wire N__12496;
    wire N__12489;
    wire N__12484;
    wire N__12481;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12462;
    wire N__12461;
    wire N__12456;
    wire N__12455;
    wire N__12454;
    wire N__12453;
    wire N__12450;
    wire N__12445;
    wire N__12442;
    wire N__12439;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12414;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12380;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12368;
    wire N__12363;
    wire N__12362;
    wire N__12359;
    wire N__12356;
    wire N__12351;
    wire N__12348;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12338;
    wire N__12335;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12276;
    wire N__12273;
    wire N__12270;
    wire N__12267;
    wire N__12264;
    wire N__12261;
    wire N__12258;
    wire N__12255;
    wire N__12252;
    wire N__12249;
    wire N__12246;
    wire N__12243;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12219;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12198;
    wire N__12195;
    wire N__12192;
    wire N__12189;
    wire N__12186;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12171;
    wire N__12168;
    wire N__12165;
    wire N__12162;
    wire N__12159;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12120;
    wire N__12117;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12087;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11967;
    wire N__11964;
    wire N__11961;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11937;
    wire N__11934;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11884;
    wire N__11883;
    wire N__11878;
    wire N__11875;
    wire N__11874;
    wire N__11873;
    wire N__11870;
    wire N__11865;
    wire N__11862;
    wire N__11861;
    wire N__11858;
    wire N__11855;
    wire N__11850;
    wire N__11847;
    wire N__11844;
    wire N__11835;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11730;
    wire N__11727;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11690;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11655;
    wire N__11652;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11613;
    wire N__11610;
    wire N__11607;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11562;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11544;
    wire N__11541;
    wire N__11538;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11520;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11502;
    wire N__11501;
    wire N__11496;
    wire N__11493;
    wire N__11492;
    wire N__11491;
    wire N__11486;
    wire N__11483;
    wire N__11480;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11337;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11319;
    wire N__11316;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11286;
    wire N__11283;
    wire N__11280;
    wire N__11277;
    wire N__11274;
    wire N__11271;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11232;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11217;
    wire N__11214;
    wire N__11211;
    wire N__11208;
    wire N__11205;
    wire N__11202;
    wire N__11199;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11184;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11169;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11151;
    wire N__11148;
    wire N__11145;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11124;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire VCCG0;
    wire GNDG0;
    wire port_nmib_0_i;
    wire this_vga_signals_vvisibility_i;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire rgb_c_2;
    wire port_clk_c;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire M_this_oam_address_qZ0Z_0;
    wire bfn_7_17_0_;
    wire M_this_oam_address_qZ0Z_1;
    wire un1_M_this_oam_address_q_cry_0;
    wire M_this_oam_address_qZ0Z_2;
    wire un1_M_this_oam_address_q_cry_1;
    wire M_this_oam_address_qZ0Z_3;
    wire un1_M_this_oam_address_q_cry_2;
    wire M_this_oam_address_qZ0Z_4;
    wire un1_M_this_oam_address_q_cry_3;
    wire un1_M_this_oam_address_q_cry_4;
    wire M_this_oam_address_qZ0Z_5;
    wire \this_oam_ram.M_this_oam_ram_read_data_19 ;
    wire M_this_data_tmp_qZ0Z_26;
    wire M_this_oam_ram_write_data_26;
    wire M_this_oam_ram_write_data_20;
    wire N_892_0;
    wire rgb_c_0;
    wire rgb_c_3;
    wire rgb_c_4;
    wire N_834_0;
    wire N_818_0;
    wire N_837_0;
    wire M_this_oam_ram_write_data_5;
    wire M_this_oam_ram_write_data_8;
    wire N_836_0;
    wire N_896_0;
    wire M_this_oam_ram_write_data_4;
    wire N_895_0;
    wire N_891_0;
    wire \this_oam_ram.M_this_oam_ram_read_data_10 ;
    wire \this_oam_ram.M_this_oam_ram_read_data_11 ;
    wire M_this_oam_ram_write_data_28;
    wire N_894_0;
    wire N_889_0;
    wire \this_ppu.M_this_oam_ram_read_data_i_16 ;
    wire bfn_9_19_0_;
    wire \this_ppu.un3_sprites_addr_cry_0 ;
    wire \this_ppu.un3_sprites_addr_cry_1 ;
    wire M_this_oam_ram_read_data_i_19;
    wire \this_ppu.un3_sprites_addr_cry_2 ;
    wire \this_ppu.un3_sprites_addr_cry_3 ;
    wire \this_ppu.un3_sprites_addr_cry_4 ;
    wire \this_ppu.un3_sprites_addr_cry_5 ;
    wire M_this_oam_ram_read_data_23;
    wire \this_ppu.un3_sprites_addr_cry_6 ;
    wire \this_oam_ram.M_this_oam_ram_read_data_21 ;
    wire M_this_oam_ram_read_data_i_21;
    wire M_this_oam_ram_write_data_0;
    wire \this_oam_ram.M_this_oam_ram_read_data_12 ;
    wire \this_oam_ram.M_this_oam_ram_read_data_17 ;
    wire M_this_oam_ram_read_data_i_17;
    wire \this_oam_ram.M_this_oam_ram_read_data_18 ;
    wire M_this_oam_ram_read_data_i_18;
    wire \this_oam_ram.M_this_oam_ram_read_data_20 ;
    wire M_this_oam_ram_read_data_i_20;
    wire this_pixel_clk_M_counter_q_i_1;
    wire this_pixel_clk_M_counter_q_0;
    wire rgb_c_1;
    wire M_this_vga_signals_address_1;
    wire N_816_0;
    wire \this_vga_ramdac.N_2612_reto ;
    wire M_this_map_address_qZ0Z_0;
    wire bfn_9_24_0_;
    wire M_this_map_address_qZ0Z_1;
    wire un1_M_this_map_address_q_cry_0;
    wire M_this_map_address_qZ0Z_2;
    wire un1_M_this_map_address_q_cry_1;
    wire M_this_map_address_qZ0Z_3;
    wire un1_M_this_map_address_q_cry_2;
    wire M_this_map_address_qZ0Z_4;
    wire un1_M_this_map_address_q_cry_3;
    wire M_this_map_address_qZ0Z_5;
    wire un1_M_this_map_address_q_cry_4;
    wire M_this_map_address_qZ0Z_6;
    wire un1_M_this_map_address_q_cry_5;
    wire M_this_map_address_qZ0Z_7;
    wire un1_M_this_map_address_q_cry_6;
    wire un1_M_this_map_address_q_cry_7;
    wire M_this_map_address_qZ0Z_8;
    wire bfn_9_25_0_;
    wire un1_M_this_map_address_q_cry_8;
    wire M_this_map_address_qZ0Z_9;
    wire \this_vga_ramdac.i2_mux ;
    wire \this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ;
    wire rgb_c_5;
    wire N_60_0;
    wire M_this_vga_signals_address_5;
    wire M_this_vga_signals_address_2;
    wire M_this_vga_signals_address_4;
    wire M_this_map_ram_read_data_1;
    wire \this_ppu.un3_sprites_addr_cry_6_c_RNIP5LZ0Z8 ;
    wire M_this_ppu_sprites_addr_7;
    wire M_this_data_tmp_qZ0Z_15;
    wire M_this_data_tmp_qZ0Z_8;
    wire M_this_data_tmp_qZ0Z_11;
    wire N_835_0;
    wire N_897_0;
    wire N_53_0;
    wire M_this_oam_ram_write_data_2;
    wire N_890_0;
    wire M_this_oam_ram_write_data_12;
    wire N_831_0;
    wire M_this_oam_ram_write_data_24;
    wire N_832_0;
    wire N_893_0;
    wire M_this_data_tmp_qZ0Z_19;
    wire M_this_data_tmp_qZ0Z_20;
    wire M_this_data_tmp_qZ0Z_21;
    wire M_this_data_tmp_qZ0Z_22;
    wire M_this_data_tmp_qZ0Z_23;
    wire \this_oam_ram.M_this_oam_ram_read_data_22 ;
    wire M_this_oam_ram_read_data_i_22;
    wire \this_vga_signals.mult1_un68_sum_axb1_cascade_ ;
    wire \this_vga_signals.if_m2_0 ;
    wire N_58_0;
    wire N_3_0_cascade_;
    wire G_480_cascade_;
    wire \this_vga_ramdac.N_2614_reto ;
    wire \this_vga_ramdac.N_2611_reto ;
    wire \this_vga_ramdac.N_2610_reto ;
    wire N_2_0;
    wire N_2_0_cascade_;
    wire M_this_vga_signals_pixel_clk_0_0;
    wire \this_vga_ramdac.i2_mux_0_cascade_ ;
    wire \this_vga_ramdac.N_2615_reto ;
    wire \this_vga_ramdac.m16_cascade_ ;
    wire G_480;
    wire \this_vga_ramdac.N_2613_reto ;
    wire N_73_0;
    wire \this_vga_ramdac.N_24_mux ;
    wire \this_vga_ramdac.m19 ;
    wire M_this_vram_read_data_0;
    wire M_this_vram_read_data_3;
    wire M_this_vram_read_data_1;
    wire M_this_vram_read_data_2;
    wire \this_vga_ramdac.m6 ;
    wire M_this_data_tmp_qZ0Z_14;
    wire M_this_data_tmp_qZ0Z_27;
    wire M_this_data_tmp_qZ0Z_3;
    wire M_this_data_tmp_qZ0Z_7;
    wire M_this_data_tmp_qZ0Z_2;
    wire M_this_data_tmp_qZ0Z_4;
    wire M_this_data_tmp_qZ0Z_25;
    wire M_this_data_tmp_qZ0Z_31;
    wire M_this_data_tmp_qZ0Z_28;
    wire N_833_0;
    wire M_this_oam_ram_read_data_16;
    wire M_this_ppu_vram_addr_i_6;
    wire M_this_data_tmp_qZ0Z_18;
    wire M_this_oam_ram_write_data_18;
    wire M_this_ppu_map_addr_4;
    wire M_this_data_tmp_qZ0Z_30;
    wire N_830_0;
    wire M_this_data_tmp_qZ0Z_16;
    wire M_this_oam_ram_write_data_16;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb1 ;
    wire \this_vga_signals.if_i4_mux_0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_0 ;
    wire \this_vga_signals.M_hcounter_q_RNIUULS4Z0Z_3 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.if_m2_2 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_3_1_cascade_ ;
    wire \this_vga_signals.d_N_3_0_i ;
    wire \this_vga_signals.mult1_un82_sum_c2_0 ;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_2_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_c3_0 ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.mult1_un75_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un82_sum_axb1 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_1 ;
    wire \this_vga_signals.mult1_un82_sum_c3 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_axb1 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_ ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2 ;
    wire \this_vga_signals.SUM_3 ;
    wire N_3_0;
    wire \this_vga_signals.M_pcounter_q_3_0 ;
    wire \this_vga_signals.N_17_0 ;
    wire \this_vga_signals.M_hcounter_q_RNI9JJM1Z0Z_0 ;
    wire \this_vga_signals.M_hcounter_q_RNIADGD1Z0Z_5_cascade_ ;
    wire this_vga_signals_hvisibility_i;
    wire \this_vga_signals.i5_mux ;
    wire this_vga_signals_hsync_1_i;
    wire M_this_ppu_map_addr_9;
    wire N_63_0;
    wire \this_vga_signals.mult1_un68_sum_c3_0 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_3 ;
    wire M_this_vga_signals_address_3;
    wire \this_vga_signals.SUM_3_1 ;
    wire M_this_vga_signals_address_6;
    wire M_this_data_tmp_qZ0Z_29;
    wire M_this_data_tmp_qZ0Z_5;
    wire M_this_data_tmp_qZ0Z_12;
    wire M_this_data_tmp_qZ0Z_13;
    wire M_this_data_tmp_qZ0Z_9;
    wire M_this_data_tmp_qZ0Z_0;
    wire M_this_ppu_vram_data_0_cascade_;
    wire \this_ppu.N_134_cascade_ ;
    wire \this_ppu.un1_M_haddress_q_c2_cascade_ ;
    wire \this_ppu.un1_M_haddress_q_c5 ;
    wire M_this_ppu_vram_addr_6;
    wire M_this_ppu_map_addr_2;
    wire \this_ppu.un1_M_haddress_q_c5_cascade_ ;
    wire \this_ppu.M_haddress_qZ0Z_7 ;
    wire bfn_12_21_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_12_22_0_;
    wire \this_vga_signals.M_pcounter_q_i_3_0 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_0 ;
    wire N_815_0;
    wire N_814_0;
    wire this_ppu_M_vaddress_q_i_6;
    wire M_this_data_tmp_qZ0Z_1;
    wire M_this_data_tmp_qZ0Z_24;
    wire M_this_data_tmp_qZ0Z_6;
    wire \this_ppu.un3_sprites_addr_cry_1_c_RNITOBZ0Z8 ;
    wire M_this_ppu_sprites_addr_2;
    wire \this_ppu.un1_M_haddress_q_c1_cascade_ ;
    wire M_this_ppu_vram_en_0;
    wire \this_ppu.N_134 ;
    wire M_this_ppu_map_addr_0;
    wire M_this_ppu_vram_addr_2;
    wire \this_ppu.un1_M_haddress_q_c2 ;
    wire M_this_ppu_map_addr_1;
    wire \this_ppu.N_128 ;
    wire \this_ppu.M_state_qc_1_3 ;
    wire M_this_ppu_vram_data_0;
    wire \this_ppu.M_state_qc_1_1_cascade_ ;
    wire \this_ppu.M_state_qZ0Z_4 ;
    wire \this_ppu.M_state_qZ0Z_5 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.N_18_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.m23_1_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.N_1090_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire G_464;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire M_this_oam_ram_write_data_10;
    wire bfn_14_18_0_;
    wire \this_ppu.un1_M_count_q_1_cry_0_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_1_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_2_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_3_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_4_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_5_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_6_s1 ;
    wire \this_ppu.M_state_d_0_sqmuxa_1_cascade_ ;
    wire \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ;
    wire \this_ppu.N_1456_0_cascade_ ;
    wire \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ;
    wire \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_5 ;
    wire \this_ppu.M_count_qZ0Z_4 ;
    wire \this_ppu.M_count_qZ0Z_1 ;
    wire \this_ppu.M_state_q_RNIE20V4Z0Z_0 ;
    wire M_this_vga_signals_line_clk_0_cascade_;
    wire \this_ppu.M_state_d_0_sqmuxa_cascade_ ;
    wire \this_vga_signals.N_1000_cascade_ ;
    wire \this_reset_cond.M_stage_qZ0Z_3 ;
    wire \this_vga_signals.M_lcounter_qZ0Z_0 ;
    wire \this_vga_signals.i21_mux_cascade_ ;
    wire \this_vga_signals.M_lcounter_qZ0Z_1 ;
    wire N_817_0;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire M_this_data_tmp_qZ0Z_10;
    wire M_this_data_tmp_qZ0Z_17;
    wire \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_3 ;
    wire \this_ppu.M_count_qZ0Z_0 ;
    wire \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_2 ;
    wire M_this_map_ram_read_data_2;
    wire \this_ppu.un10_sprites_addr_axb_0_cascade_ ;
    wire M_this_ppu_sprites_addr_8;
    wire \this_ppu.un10_0 ;
    wire \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ;
    wire \this_ppu.N_1456_0 ;
    wire \this_ppu.M_count_qZ0Z_6 ;
    wire \this_ppu.un3_sprites_addr_cry_2_c_RNIVRCZ0Z8 ;
    wire M_this_ppu_sprites_addr_3;
    wire \this_oam_ram.M_this_oam_ram_read_data_9 ;
    wire M_this_map_ram_read_data_3;
    wire M_this_ppu_sprites_addr_9;
    wire \this_ppu.M_state_d_0_sqmuxa_1 ;
    wire \this_ppu.M_count_q_RNO_0Z0Z_7 ;
    wire \this_ppu.M_count_qZ0Z_7 ;
    wire \this_vga_signals.N_129_mux ;
    wire \this_vga_signals.N_1028 ;
    wire \this_vga_signals.N_1028_cascade_ ;
    wire \this_vga_signals.N_999 ;
    wire \this_vga_signals.N_1004_cascade_ ;
    wire \this_vga_signals.N_1013 ;
    wire \this_vga_signals.N_1013_cascade_ ;
    wire \this_vga_signals.N_105_mux_cascade_ ;
    wire \this_vga_signals.N_113_mux ;
    wire \this_reset_cond.M_stage_qZ0Z_4 ;
    wire \this_reset_cond.M_stage_qZ0Z_5 ;
    wire this_vga_signals_vvisibility;
    wire M_this_reset_cond_out_0;
    wire \this_reset_cond.M_stage_qZ0Z_6 ;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_7 ;
    wire \this_reset_cond.M_stage_qZ0Z_8 ;
    wire \this_vga_signals.vaddress_ac0_9_0_a0_2 ;
    wire \this_ppu.M_vaddress_qZ0Z_6 ;
    wire \this_ppu.un1_M_vaddress_q_c5 ;
    wire \this_ppu.M_vaddress_qZ0Z_7 ;
    wire dma_0_i;
    wire N_1430_0;
    wire M_this_state_q_ns_17_cascade_;
    wire M_this_state_q_ns_0_17;
    wire M_this_map_ram_read_data_6;
    wire M_this_oam_ram_read_data_8;
    wire \this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ;
    wire bfn_16_19_0_;
    wire M_this_oam_ram_read_data_i_9;
    wire \this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5BZ0 ;
    wire \this_ppu.un10_sprites_addr_cry_0 ;
    wire M_this_oam_ram_read_data_i_10;
    wire \this_ppu.un10_sprites_addr_cry_1 ;
    wire M_this_oam_ram_read_data_i_11;
    wire \this_ppu.un10_sprites_addr_cry_2 ;
    wire M_this_oam_ram_read_data_i_12;
    wire \this_ppu.un10_sprites_addr_cry_3_c_RNISS8BZ0 ;
    wire \this_ppu.un10_sprites_addr_cry_3 ;
    wire M_this_oam_ram_read_data_13;
    wire \this_ppu.un10_sprites_addr_cry_4 ;
    wire \this_ppu.M_last_q ;
    wire \this_ppu.M_state_qZ0Z_0 ;
    wire M_this_vga_signals_line_clk_0;
    wire \this_ppu.M_state_d_0_sqmuxa ;
    wire M_this_ppu_vram_addr_7;
    wire M_this_ppu_map_addr_7;
    wire \this_ppu.un1_M_vaddress_q_c3 ;
    wire M_this_ppu_map_addr_5;
    wire M_this_ppu_map_addr_6;
    wire \this_ppu.M_state_q_RNIELANCZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_q_esr_RNI4KCU6Z0Z_9 ;
    wire \this_vga_signals.g1_2_0_0_cascade_ ;
    wire M_this_vga_ramdac_en_0;
    wire \this_vga_signals.mult1_un75_sum_c3_0_0_0_0_cascade_ ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.un6_vvisibilitylt9_0 ;
    wire \this_vga_signals.g2_2 ;
    wire \this_vga_signals.SUM_2_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_1_1_cascade_ ;
    wire \this_vga_signals.N_4_0_0_0 ;
    wire \this_vga_signals.g3_2_0 ;
    wire \this_vga_signals.N_6_cascade_ ;
    wire \this_vga_signals.g4 ;
    wire N_1438_0;
    wire \this_start_data_delay.port_data_rw_0_a2Z0Z_1 ;
    wire port_data_rw_0_i;
    wire \this_sprites_ram.mem_out_bus5_2 ;
    wire \this_sprites_ram.mem_out_bus1_2 ;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire \this_sprites_ram.mem_out_bus4_2 ;
    wire \this_sprites_ram.mem_out_bus0_2 ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ;
    wire M_this_ppu_vram_data_2;
    wire \this_ppu.un10_sprites_addr_cry_2_c_RNIQP7BZ0 ;
    wire M_this_map_ram_read_data_5;
    wire \this_sprites_ram.mem_out_bus7_2 ;
    wire \this_sprites_ram.mem_out_bus3_2 ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ;
    wire \this_ppu.M_state_qZ0Z_1 ;
    wire \this_ppu.M_state_q_srsts_i_a3_5_2 ;
    wire \this_ppu.M_state_q_srsts_i_a3_4_2 ;
    wire N_2_cascade_;
    wire \this_vga_signals.N_6_1_cascade_ ;
    wire \this_vga_signals.vaddress_N_4_0 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un75_sum_axb1_i_1 ;
    wire \this_vga_signals.N_7_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c2_0 ;
    wire \this_vga_signals.if_m2_3_1_cascade_ ;
    wire \this_vga_signals.g2_cascade_ ;
    wire \this_vga_signals.g0_4 ;
    wire \this_vga_signals.g1_0_0 ;
    wire \this_vga_signals.if_m1_0_cascade_ ;
    wire \this_vga_signals.N_129_i ;
    wire \this_vga_signals.if_m1_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0 ;
    wire \this_vga_signals.g0_3_0_a3 ;
    wire \this_vga_signals.g1_0 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_1_0_cascade_ ;
    wire \this_vga_signals.g0_i_x4_7_0_0 ;
    wire \this_vga_signals.g0_9_N_2L1_cascade_ ;
    wire \this_vga_signals.g0_i_x4_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_1_0_0_cascade_ ;
    wire \this_vga_signals.g0_9_N_3L3 ;
    wire \this_vga_signals.g0_i_a4_4_0_0 ;
    wire N_1422_0;
    wire M_this_state_d_0_sqmuxa_2_cascade_;
    wire M_this_state_d_0_sqmuxa_2;
    wire \this_start_data_delay.N_65_cascade_ ;
    wire \this_start_data_delay.N_42_0 ;
    wire \this_start_data_delay.N_43_0 ;
    wire dma_0;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_0_2_cascade_ ;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_cascade_;
    wire \this_vga_signals.mult1_un61_sum_c3_0 ;
    wire \this_vga_signals.if_m2 ;
    wire \this_vga_signals.if_m1_9_0 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_cascade_ ;
    wire \this_vga_signals.if_m2_3_1 ;
    wire \this_vga_signals.if_i4_mux ;
    wire \this_vga_signals.g0_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_0_2_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_0_2_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb2_0_cascade_ ;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d;
    wire \this_vga_signals.g2_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2 ;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_cascade_;
    wire \this_vga_signals.mult1_un61_sum_c3_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3 ;
    wire \this_vga_signals.mult1_un75_sum_axb1_i_0 ;
    wire \this_vga_signals.N_4_2_cascade_ ;
    wire \this_vga_signals.if_m1_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_axb2_0 ;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1;
    wire \this_vga_signals.mult1_un75_sum_axb1_1 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_4_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_cascade_ ;
    wire \this_vga_signals.N_4_3_0_cascade_ ;
    wire \this_vga_signals.N_14_0 ;
    wire \this_vga_signals.g1 ;
    wire \this_vga_signals.g0_10_1 ;
    wire \this_vga_signals.N_24_mux ;
    wire \this_vga_signals.g1_2 ;
    wire \this_vga_signals.g0_3_0_a3_3 ;
    wire \this_vga_signals.mult1_un54_sum_axb1 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_cascade_ ;
    wire \this_vga_signals.if_N_9_i ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i ;
    wire \this_vga_signals.SUM_2_0_1 ;
    wire \this_vga_signals.mult1_un47_sum_c3_1_0 ;
    wire \this_vga_signals.mult1_un47_sum_c3_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire \this_vga_signals.g2_4 ;
    wire \this_vga_signals.m12_0_1 ;
    wire \this_start_data_delay.N_400 ;
    wire led23;
    wire \this_start_data_delay.dmalto4_0_a2Z0Z_1 ;
    wire \this_start_data_delay.N_115 ;
    wire \this_start_data_delay.N_69 ;
    wire port_address_in_5;
    wire port_address_in_6;
    wire \this_start_data_delay.N_47_0_cascade_ ;
    wire \this_start_data_delay.N_48_0_cascade_ ;
    wire N_28_0;
    wire \this_start_data_delay.N_82 ;
    wire \this_start_data_delay.N_82_cascade_ ;
    wire M_this_substate_qZ0;
    wire \this_vga_signals.g0_0_x4_0_0 ;
    wire \this_vga_signals.vaddress_c2_cascade_ ;
    wire \this_vga_signals.N_5_2_1_cascade_ ;
    wire \this_vga_signals.g0_5_0_cascade_ ;
    wire \this_vga_signals.g0_1_1_cascade_ ;
    wire \this_vga_signals.N_3_2 ;
    wire \this_vga_signals.g0_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1 ;
    wire \this_vga_signals.g0_5_2_0 ;
    wire \this_vga_signals.g2_1_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_2_1 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_0_a4 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_0_1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_3_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_602_ns ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_4_x1 ;
    wire \this_vga_signals.mult1_un47_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_2 ;
    wire \this_vga_signals.i1_mux ;
    wire \this_vga_signals.mult1_un47_sum_axbxc1_0 ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_4_x0 ;
    wire \this_vga_signals.g1_7 ;
    wire \this_vga_signals.vaddress_3_6 ;
    wire \this_ppu.un3_sprites_addr_axb_0 ;
    wire M_this_ppu_vram_addr_0;
    wire M_this_ppu_sprites_addr_0;
    wire M_this_state_qZ0Z_15;
    wire M_this_state_qZ0Z_14;
    wire M_this_state_qZ0Z_13;
    wire \this_start_data_delay.N_112_0 ;
    wire \this_start_data_delay.N_80_0 ;
    wire \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_aZ0Z2_cascade_ ;
    wire \this_start_data_delay.N_76_1 ;
    wire \this_start_data_delay.N_127_cascade_ ;
    wire M_this_state_qZ0Z_11;
    wire \this_start_data_delay.N_844_0_cascade_ ;
    wire \this_start_data_delay.N_151_cascade_ ;
    wire \this_start_data_delay.N_89_0 ;
    wire M_this_state_qZ0Z_16;
    wire \this_start_data_delay.N_47_0 ;
    wire \this_start_data_delay.N_909_0_cascade_ ;
    wire led_c_1;
    wire \this_start_data_delay.M_this_state_q_ns_0_i_0_0 ;
    wire \this_start_data_delay.M_this_state_q_ns_0_i_2_0_0 ;
    wire N_822_0;
    wire \this_start_data_delay.N_910_cascade_ ;
    wire M_this_state_qZ0Z_10;
    wire \this_start_data_delay.N_90_0 ;
    wire port_address_in_1;
    wire port_address_in_0;
    wire port_address_in_2;
    wire \this_start_data_delay.N_48_0 ;
    wire \this_start_data_delay.N_71 ;
    wire \this_start_data_delay.N_67 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_2_1_0 ;
    wire \this_vga_signals.N_4558_0 ;
    wire \this_vga_signals.g0_4_i_a3_1_cascade_ ;
    wire \this_vga_signals.g0_4_i_1_cascade_ ;
    wire \this_vga_signals.N_6_2 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_602_x0 ;
    wire \this_vga_signals.vaddress_c2 ;
    wire \this_vga_signals.r_N_4_mux ;
    wire \this_vga_signals.r_N_4_mux_cascade_ ;
    wire \this_vga_signals.SUM_2 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_ns ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x0 ;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_602_x1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_3_x1 ;
    wire \this_vga_signals.N_4_0 ;
    wire \this_vga_signals.g0_6_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_c3 ;
    wire \this_vga_signals.N_4_0_0_1 ;
    wire \this_vga_signals.vaddress_0_5 ;
    wire \this_vga_signals.vaddress_0_6_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_c3_0 ;
    wire \this_vga_signals.M_vcounter_q_5_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z1 ;
    wire \this_vga_signals.vaddress_5 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i ;
    wire \this_vga_signals.g2_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_2 ;
    wire \this_vga_signals.g0_i_x4_0_0 ;
    wire \this_vga_signals.g0_3_0_a3_1 ;
    wire \this_vga_signals.vaddress_1_6 ;
    wire \this_ppu.un3_sprites_addr_cry_0_c_RNIRLAZ0Z8 ;
    wire M_this_ppu_vram_addr_1;
    wire M_this_ppu_sprites_addr_1;
    wire \this_sprites_ram.mem_out_bus4_1 ;
    wire \this_sprites_ram.mem_out_bus0_1 ;
    wire M_this_state_qZ0Z_12;
    wire \this_start_data_delay.N_125 ;
    wire \this_start_data_delay.un30_0_0_cascade_ ;
    wire N_554_0_cascade_;
    wire M_this_state_qZ0Z_2;
    wire \this_start_data_delay.N_109_cascade_ ;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_4 ;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire \this_start_data_delay.M_last_qZ0 ;
    wire port_enb_c;
    wire M_this_delay_clk_out_0;
    wire \this_start_data_delay.N_91_0_cascade_ ;
    wire M_this_state_qZ0Z_1;
    wire \this_start_data_delay.N_110_cascade_ ;
    wire M_this_state_qZ0Z_4;
    wire \this_sprites_ram.mem_out_bus5_1 ;
    wire \this_sprites_ram.mem_out_bus1_1 ;
    wire \this_sprites_ram.mem_out_bus6_1 ;
    wire \this_sprites_ram.mem_out_bus2_1 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0_cascade_ ;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ;
    wire M_this_ppu_vram_data_1;
    wire \this_start_data_delay.M_this_state_q_ns_0_i_2_0 ;
    wire this_vga_signals_M_hcounter_d7_0;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire bfn_21_20_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire G_442;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire bfn_21_21_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire \this_vga_signals.N_4557_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire \this_vga_signals.M_vcounter_q_8_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_7_repZ0Z1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_601 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.N_1090_0 ;
    wire \this_vga_signals.N_1358_g ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire \this_vga_signals.m58_1 ;
    wire \this_vga_signals.m58_0 ;
    wire \this_vga_signals.m58_4_cascade_ ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire this_vga_signals_vsync_1_i;
    wire M_this_state_qZ0Z_3;
    wire \this_start_data_delay.N_123_cascade_ ;
    wire N_812_0;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_7 ;
    wire \this_start_data_delay.N_129_cascade_ ;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_12_cascade_ ;
    wire M_this_state_qZ0Z_8;
    wire \this_start_data_delay.N_821_0_cascade_ ;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_11 ;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_10_cascade_ ;
    wire \this_sprites_ram.mem_out_bus7_1 ;
    wire \this_sprites_ram.mem_out_bus3_1 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ;
    wire \this_start_data_delay.N_55_0 ;
    wire \this_start_data_delay.N_84 ;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_2_cascade_ ;
    wire \this_start_data_delay.N_913_cascade_ ;
    wire M_this_state_qZ0Z_9;
    wire M_this_state_qZ0Z_7;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_3_cascade_ ;
    wire M_this_map_ram_read_data_7;
    wire \this_ppu.un10_sprites_addr_cry_4_c_RNIUV9BZ0 ;
    wire \this_start_data_delay.N_91_0 ;
    wire \this_start_data_delay.N_149_cascade_ ;
    wire M_this_state_qZ0Z_6;
    wire \this_start_data_delay.N_555_0 ;
    wire \this_start_data_delay.M_this_data_count_qlde_i_a3_0 ;
    wire \this_start_data_delay.M_this_data_count_qlde_i_2_tz_0 ;
    wire \this_start_data_delay.N_820_0_cascade_ ;
    wire \this_start_data_delay.N_151 ;
    wire \this_start_data_delay.N_820_0 ;
    wire \this_start_data_delay.M_this_data_count_qlde_i_1_cascade_ ;
    wire \this_start_data_delay.N_68 ;
    wire M_this_state_qZ0Z_5;
    wire N_554_0;
    wire this_start_data_delay_M_this_data_count_q_3_0_a3_0_6_cascade_;
    wire N_911;
    wire M_this_data_count_q_3_0_13;
    wire \this_start_data_delay.N_93_0 ;
    wire \this_start_data_delay.N_122 ;
    wire \this_start_data_delay.N_149 ;
    wire \this_start_data_delay.N_121 ;
    wire \this_start_data_delay.N_938_0 ;
    wire N_813_0;
    wire port_data_c_5;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_6_cascade_ ;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_1_cascade_ ;
    wire \this_start_data_delay.N_993 ;
    wire \this_start_data_delay.N_109 ;
    wire bfn_23_17_0_;
    wire M_this_sprites_address_qZ0Z_1;
    wire un1_M_this_sprites_address_q_cry_0_THRU_CO;
    wire un1_M_this_sprites_address_q_cry_0;
    wire M_this_sprites_address_qZ0Z_2;
    wire un1_M_this_sprites_address_q_cry_1_THRU_CO;
    wire un1_M_this_sprites_address_q_cry_1;
    wire M_this_sprites_address_qZ0Z_3;
    wire un1_M_this_sprites_address_q_cry_2_THRU_CO;
    wire un1_M_this_sprites_address_q_cry_2;
    wire M_this_sprites_address_qZ0Z_4;
    wire un1_M_this_sprites_address_q_cry_3_THRU_CO;
    wire un1_M_this_sprites_address_q_cry_3;
    wire un1_M_this_sprites_address_q_cry_4;
    wire M_this_sprites_address_qZ0Z_6;
    wire un1_M_this_sprites_address_q_cry_5_THRU_CO;
    wire un1_M_this_sprites_address_q_cry_5;
    wire M_this_sprites_address_qZ0Z_7;
    wire un1_M_this_sprites_address_q_cry_6_THRU_CO;
    wire un1_M_this_sprites_address_q_cry_6;
    wire un1_M_this_sprites_address_q_cry_7;
    wire bfn_23_18_0_;
    wire un1_M_this_sprites_address_q_cry_8;
    wire M_this_sprites_address_qZ0Z_10;
    wire un1_M_this_sprites_address_q_cry_9_THRU_CO;
    wire un1_M_this_sprites_address_q_cry_9;
    wire un1_M_this_sprites_address_q_cry_10_THRU_CO;
    wire un1_M_this_sprites_address_q_cry_10;
    wire un1_M_this_sprites_address_q_cry_11_THRU_CO;
    wire un1_M_this_sprites_address_q_cry_11;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_13 ;
    wire un1_M_this_sprites_address_q_cry_12;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_0 ;
    wire un30_0;
    wire M_this_sprites_address_qZ0Z_0;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_9 ;
    wire un1_M_this_sprites_address_q_cry_8_THRU_CO;
    wire M_this_sprites_address_qZ0Z_9;
    wire \this_start_data_delay.N_86_0 ;
    wire M_this_reset_cond_out_g_0;
    wire \this_sprites_ram.mem_out_bus5_3 ;
    wire \this_sprites_ram.mem_out_bus1_3 ;
    wire N_10_0;
    wire \this_start_data_delay.M_this_state_d62Z0Z_11 ;
    wire \this_start_data_delay.M_this_state_d62Z0Z_10 ;
    wire \this_start_data_delay.M_this_state_d62Z0Z_9_cascade_ ;
    wire \this_start_data_delay.M_this_state_d62Z0Z_8 ;
    wire \this_start_data_delay.M_this_state_dZ0Z62 ;
    wire M_this_data_count_q_3_10;
    wire this_start_data_delay_M_this_external_address_q_3_i_0_15;
    wire N_116;
    wire M_this_external_address_q_3_0_13;
    wire M_this_map_ram_read_data_0;
    wire \this_ppu.un3_sprites_addr_cry_5_c_RNI55GZ0Z8 ;
    wire M_this_ppu_sprites_addr_6;
    wire \this_sprites_ram.mem_WE_10 ;
    wire \this_sprites_ram.mem_WE_8 ;
    wire \this_sprites_ram.mem_WE_12 ;
    wire \this_sprites_ram.mem_WE_14 ;
    wire N_811_0;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_5 ;
    wire un1_M_this_sprites_address_q_cry_4_THRU_CO;
    wire M_this_sprites_address_qZ0Z_5;
    wire \this_sprites_ram.mem_WE_6 ;
    wire \this_sprites_ram.mem_out_bus5_0 ;
    wire \this_sprites_ram.mem_out_bus1_0 ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ;
    wire port_data_c_0;
    wire port_data_c_4;
    wire port_data_c_6;
    wire \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3Z0Z_0_cascade_ ;
    wire \this_start_data_delay.N_902_0 ;
    wire \this_start_data_delay.N_821_0 ;
    wire port_data_c_7;
    wire \this_start_data_delay.N_123 ;
    wire N_41_0;
    wire \this_sprites_ram.mem_out_bus4_0 ;
    wire \this_sprites_ram.mem_out_bus0_0 ;
    wire \this_sprites_ram.mem_out_bus4_3 ;
    wire \this_sprites_ram.mem_out_bus0_3 ;
    wire \this_sprites_ram.mem_out_bus6_3 ;
    wire \this_sprites_ram.mem_out_bus2_3 ;
    wire \this_start_data_delay.N_992 ;
    wire \this_start_data_delay.N_110 ;
    wire un1_M_this_sprites_address_q_cry_7_THRU_CO;
    wire \this_start_data_delay.M_this_sprites_address_q_0_0_0_8_cascade_ ;
    wire \this_start_data_delay.N_990 ;
    wire M_this_sprites_address_qZ0Z_8;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ;
    wire M_this_ppu_vram_data_3;
    wire \this_sprites_ram.mem_out_bus6_0 ;
    wire \this_sprites_ram.mem_out_bus2_0 ;
    wire \this_sprites_ram.mem_radregZ0Z_12 ;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0_cascade_ ;
    wire \this_sprites_ram.mem_radregZ0Z_11 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ;
    wire \this_sprites_ram.mem_out_bus6_2 ;
    wire \this_sprites_ram.mem_out_bus2_2 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ;
    wire \this_sprites_ram.mem_WE_4 ;
    wire \this_sprites_ram.mem_out_bus7_0 ;
    wire \this_sprites_ram.mem_out_bus3_0 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ;
    wire M_this_data_count_qZ0Z_0;
    wire bfn_24_21_0_;
    wire M_this_data_count_qZ0Z_1;
    wire M_this_data_count_q_cry_0_THRU_CO;
    wire M_this_data_count_q_cry_0;
    wire M_this_data_count_qZ0Z_2;
    wire M_this_data_count_q_cry_1_THRU_CO;
    wire M_this_data_count_q_cry_1;
    wire M_this_data_count_qZ0Z_3;
    wire M_this_data_count_q_cry_2_THRU_CO;
    wire M_this_data_count_q_cry_2;
    wire M_this_data_count_q_cry_3;
    wire M_this_data_count_qZ0Z_5;
    wire M_this_data_count_q_cry_4_THRU_CO;
    wire M_this_data_count_q_cry_4;
    wire M_this_data_count_qZ0Z_6;
    wire M_this_data_count_q_s_6;
    wire M_this_data_count_q_cry_5;
    wire M_this_data_count_qZ0Z_7;
    wire M_this_data_count_q_cry_6_THRU_CO;
    wire M_this_data_count_q_cry_6;
    wire M_this_data_count_q_cry_7;
    wire M_this_data_count_qZ0Z_8;
    wire M_this_data_count_q_s_8;
    wire bfn_24_22_0_;
    wire M_this_data_count_qZ0Z_9;
    wire M_this_data_count_q_s_9;
    wire M_this_data_count_q_cry_8;
    wire M_this_data_count_qZ0Z_10;
    wire M_this_data_count_q_cry_9_THRU_CO;
    wire M_this_data_count_q_cry_9;
    wire M_this_data_count_qZ0Z_11;
    wire M_this_data_count_q_s_11;
    wire M_this_data_count_q_cry_10;
    wire M_this_data_count_qZ0Z_12;
    wire M_this_data_count_q_s_12;
    wire M_this_data_count_q_cry_11;
    wire M_this_data_count_qZ0Z_13;
    wire M_this_data_count_q_cry_12_THRU_CO;
    wire M_this_data_count_q_cry_12;
    wire CONSTANT_ONE_NET;
    wire M_this_data_count_qZ0Z_14;
    wire M_this_data_count_q_s_14;
    wire M_this_data_count_q_cry_13;
    wire M_this_data_count_qZ0Z_15;
    wire M_this_data_count_q_cry_14;
    wire M_this_data_count_q_s_15;
    wire M_this_data_count_q_cry_3_THRU_CO;
    wire N_33;
    wire M_this_data_count_qZ0Z_4;
    wire N_35;
    wire M_this_external_address_q_3_0_12;
    wire M_this_external_address_q_3_14;
    wire port_data_c_1;
    wire \this_sprites_ram.mem_WE_2 ;
    wire M_this_sprites_ram_write_en_0;
    wire M_this_sprites_address_qZ0Z_12;
    wire M_this_sprites_address_qZ0Z_11;
    wire M_this_sprites_address_qZ0Z_13;
    wire \this_sprites_ram.mem_WE_0 ;
    wire M_this_map_ram_read_data_4;
    wire \this_ppu.un10_sprites_addr_cry_1_c_RNIOM6BZ0 ;
    wire M_this_ppu_sprites_addr_10;
    wire \this_ppu.M_vaddress_qZ0Z_2 ;
    wire \this_ppu.un3_sprites_addr_cry_4_c_RNI32FZ0Z8 ;
    wire M_this_ppu_sprites_addr_5;
    wire \this_sprites_ram.mem_out_bus7_3 ;
    wire \this_sprites_ram.mem_out_bus3_3 ;
    wire \this_sprites_ram.mem_radregZ0Z_13 ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ;
    wire M_this_external_address_qZ0Z_0;
    wire bfn_26_23_0_;
    wire M_this_external_address_qZ0Z_1;
    wire M_this_external_address_q_cry_0;
    wire M_this_external_address_qZ0Z_2;
    wire M_this_external_address_q_cry_1;
    wire M_this_external_address_qZ0Z_3;
    wire M_this_external_address_q_cry_2;
    wire M_this_external_address_qZ0Z_4;
    wire M_this_external_address_q_cry_3;
    wire M_this_external_address_qZ0Z_5;
    wire M_this_external_address_q_cry_4;
    wire M_this_external_address_qZ0Z_6;
    wire M_this_external_address_q_cry_5;
    wire M_this_external_address_qZ0Z_7;
    wire M_this_external_address_q_cry_6;
    wire M_this_external_address_q_cry_7;
    wire M_this_external_address_qZ0Z_8;
    wire M_this_external_address_q_s_8;
    wire bfn_26_24_0_;
    wire M_this_external_address_qZ0Z_9;
    wire M_this_external_address_q_s_9;
    wire M_this_external_address_q_cry_8;
    wire M_this_external_address_q_cry_9;
    wire M_this_external_address_q_cry_10;
    wire M_this_external_address_qZ0Z_12;
    wire M_this_external_address_q_cry_11_THRU_CO;
    wire M_this_external_address_q_cry_11;
    wire M_this_external_address_qZ0Z_13;
    wire M_this_external_address_q_cry_12_THRU_CO;
    wire M_this_external_address_q_cry_12;
    wire M_this_external_address_qZ0Z_14;
    wire M_this_external_address_q_cry_13_THRU_CO;
    wire M_this_external_address_q_cry_13;
    wire M_this_external_address_qZ0Z_15;
    wire M_this_external_address_q_cry_14;
    wire M_this_external_address_q_s_15;
    wire M_this_external_address_q_s_11;
    wire port_data_c_3;
    wire M_this_external_address_qZ0Z_11;
    wire M_this_external_address_q_s_10;
    wire M_this_external_address_d_1_sqmuxa;
    wire port_data_c_2;
    wire N_39;
    wire M_this_external_address_qZ0Z_10;
    wire clk_0_c_g;
    wire N_37;
    wire \this_ppu.M_vaddress_qZ0Z_1 ;
    wire \this_ppu.M_state_qZ0Z_3 ;
    wire \this_ppu.M_state_qZ0Z_2 ;
    wire \this_ppu.un3_sprites_addr_cry_3_c_RNI1VDZ0Z8 ;
    wire M_this_ppu_sprites_addr_4;
    wire port_address_in_7;
    wire port_address_in_4;
    wire port_rw_in;
    wire port_address_in_3;
    wire \this_start_data_delay.un1_M_this_state_q_17_i_o2_1Z0Z_4 ;
    wire _gnd_net_;

    defparam \this_map_ram.mem_mem_0_0_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_0_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,M_this_map_ram_read_data_3,dangling_wire_2,dangling_wire_3,dangling_wire_4,M_this_map_ram_read_data_2,dangling_wire_5,dangling_wire_6,dangling_wire_7,M_this_map_ram_read_data_1,dangling_wire_8,dangling_wire_9,dangling_wire_10,M_this_map_ram_read_data_0,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__13431,N__13662,N__16782,N__16638,N__16701,N__12840,N__12891,N__13584,N__13827,N__13962}),
            .WADDR({dangling_wire_13,N__11931,N__11964,N__11994,N__11589,N__11619,N__11649,N__11679,N__11709,N__11739,N__11766}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__13689,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__11796,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__15012,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__12633,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__32649),
            .RE(N__29819),
            .WCLKE(N__19898),
            .WCLK(N__32650),
            .WE(N__29837));
    defparam \this_map_ram.mem_mem_0_1_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_1_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_42,dangling_wire_43,M_this_map_ram_read_data_7,dangling_wire_44,dangling_wire_45,dangling_wire_46,M_this_map_ram_read_data_6,dangling_wire_47,dangling_wire_48,dangling_wire_49,M_this_map_ram_read_data_5,dangling_wire_50,dangling_wire_51,dangling_wire_52,M_this_map_ram_read_data_4,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__13425,N__13656,N__16776,N__16632,N__16695,N__12834,N__12885,N__13578,N__13821,N__13956}),
            .WADDR({dangling_wire_55,N__11925,N__11958,N__11988,N__11583,N__11613,N__11643,N__11673,N__11703,N__11733,N__11760}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__12405,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__11826,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__13410,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__13677,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__32655),
            .RE(N__29841),
            .WCLKE(N__19899),
            .WCLK(N__32656),
            .WE(N__29836));
    defparam \this_oam_ram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_84,dangling_wire_85,M_this_oam_ram_read_data_13,\this_oam_ram.M_this_oam_ram_read_data_12 ,\this_oam_ram.M_this_oam_ram_read_data_11 ,\this_oam_ram.M_this_oam_ram_read_data_10 ,\this_oam_ram.M_this_oam_ram_read_data_9 ,M_this_oam_ram_read_data_8,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93}),
            .RADDR({dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104}),
            .WADDR({dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,N__11211,N__11241,N__11010,N__11037,N__11067,N__11094}),
            .MASK({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125}),
            .WDATA({N__11301,N__11289,N__11385,N__12258,N__11247,N__14709,N__12039,N__11259,N__11253,N__12018,N__11268,N__11394,N__12030,N__12006,N__11280,N__11559}),
            .RCLKE(),
            .RCLK(N__32605),
            .RE(N__29755),
            .WCLKE(N__18621),
            .WCLK(N__32606),
            .WE(N__29794));
    defparam \this_oam_ram.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,M_this_oam_ram_read_data_23,\this_oam_ram.M_this_oam_ram_read_data_22 ,\this_oam_ram.M_this_oam_ram_read_data_21 ,\this_oam_ram.M_this_oam_ram_read_data_20 ,\this_oam_ram.M_this_oam_ram_read_data_19 ,\this_oam_ram.M_this_oam_ram_read_data_18 ,\this_oam_ram.M_this_oam_ram_read_data_17 ,M_this_oam_ram_read_data_16}),
            .RADDR({dangling_wire_134,dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144}),
            .WADDR({dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,N__11205,N__11235,N__11004,N__11031,N__11061,N__11088}),
            .MASK({dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165}),
            .WDATA({N__11340,N__12801,N__12270,N__11355,N__11376,N__11172,N__12249,N__12237,N__11160,N__12225,N__12213,N__11166,N__11349,N__12855,N__12921,N__12786}),
            .RCLKE(),
            .RCLK(N__32621),
            .RE(N__29790),
            .WCLKE(N__18622),
            .WCLK(N__32622),
            .WE(N__29795));
    defparam \this_sprites_ram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,\this_sprites_ram.mem_out_bus0_1 ,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,\this_sprites_ram.mem_out_bus0_0 ,dangling_wire_177,dangling_wire_178,dangling_wire_179}),
            .RADDR({N__30390,N__15570,N__15291,N__12162,N__26661,N__30234,N__31791,N__15714,N__14121,N__20877,N__19251}),
            .WADDR({N__25539,N__26409,N__27483,N__25689,N__25824,N__27174,N__24852,N__24996,N__25137,N__25272,N__26559}),
            .MASK({dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195}),
            .WDATA({dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,N__22134,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,N__24584,dangling_wire_207,dangling_wire_208,dangling_wire_209}),
            .RCLKE(),
            .RCLK(N__32524),
            .RE(N__29789),
            .WCLKE(N__27282),
            .WCLK(N__32525),
            .WE(N__29787));
    defparam \this_sprites_ram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,\this_sprites_ram.mem_out_bus0_3 ,dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,\this_sprites_ram.mem_out_bus0_2 ,dangling_wire_221,dangling_wire_222,dangling_wire_223}),
            .RADDR({N__30384,N__15564,N__15285,N__12156,N__26655,N__30228,N__31785,N__15708,N__14115,N__20871,N__19245}),
            .WADDR({N__25533,N__26403,N__27477,N__25683,N__25818,N__27168,N__24846,N__24990,N__25131,N__25266,N__26553}),
            .MASK({dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239}),
            .WDATA({dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,N__27803,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,N__27246,dangling_wire_251,dangling_wire_252,dangling_wire_253}),
            .RCLKE(),
            .RCLK(N__32526),
            .RE(N__29788),
            .WCLKE(N__27278),
            .WCLK(N__32527),
            .WE(N__29511));
    defparam \this_sprites_ram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,\this_sprites_ram.mem_out_bus1_1 ,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,\this_sprites_ram.mem_out_bus1_0 ,dangling_wire_265,dangling_wire_266,dangling_wire_267}),
            .RADDR({N__30378,N__15558,N__15279,N__12150,N__26649,N__30222,N__31779,N__15702,N__14109,N__20865,N__19239}),
            .WADDR({N__25527,N__26397,N__27471,N__25677,N__25812,N__27162,N__24840,N__24984,N__25125,N__25260,N__26547}),
            .MASK({dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283}),
            .WDATA({dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,N__22129,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,N__24576,dangling_wire_295,dangling_wire_296,dangling_wire_297}),
            .RCLKE(),
            .RCLK(N__32528),
            .RE(N__29744),
            .WCLKE(N__27303),
            .WCLK(N__32529),
            .WE(N__29739));
    defparam \this_sprites_ram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,\this_sprites_ram.mem_out_bus1_3 ,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,dangling_wire_308,\this_sprites_ram.mem_out_bus1_2 ,dangling_wire_309,dangling_wire_310,dangling_wire_311}),
            .RADDR({N__30372,N__15552,N__15273,N__12144,N__26643,N__30216,N__31773,N__15696,N__14103,N__20859,N__19233}),
            .WADDR({N__25521,N__26391,N__27465,N__25671,N__25806,N__27156,N__24834,N__24978,N__25119,N__25254,N__26541}),
            .MASK({dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327}),
            .WDATA({dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,N__27795,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,N__27233,dangling_wire_339,dangling_wire_340,dangling_wire_341}),
            .RCLKE(),
            .RCLK(N__32532),
            .RE(N__29743),
            .WCLKE(N__27299),
            .WCLK(N__32533),
            .WE(N__29735));
    defparam \this_sprites_ram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,\this_sprites_ram.mem_out_bus2_1 ,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,dangling_wire_352,\this_sprites_ram.mem_out_bus2_0 ,dangling_wire_353,dangling_wire_354,dangling_wire_355}),
            .RADDR({N__30366,N__15546,N__15267,N__12138,N__26637,N__30210,N__31767,N__15690,N__14097,N__20853,N__19227}),
            .WADDR({N__25515,N__26385,N__27459,N__25665,N__25800,N__27150,N__24828,N__24972,N__25113,N__25248,N__26535}),
            .MASK({dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371}),
            .WDATA({dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,N__22118,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,N__24562,dangling_wire_383,dangling_wire_384,dangling_wire_385}),
            .RCLKE(),
            .RCLK(N__32540),
            .RE(N__29651),
            .WCLKE(N__27348),
            .WCLK(N__32539),
            .WE(N__29664));
    defparam \this_sprites_ram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,\this_sprites_ram.mem_out_bus2_3 ,dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,\this_sprites_ram.mem_out_bus2_2 ,dangling_wire_397,dangling_wire_398,dangling_wire_399}),
            .RADDR({N__30360,N__15540,N__15261,N__12132,N__26631,N__30204,N__31761,N__15684,N__14091,N__20847,N__19221}),
            .WADDR({N__25509,N__26379,N__27453,N__25659,N__25794,N__27144,N__24822,N__24966,N__25107,N__25242,N__26529}),
            .MASK({dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415}),
            .WDATA({dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,N__27781,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,N__27218,dangling_wire_427,dangling_wire_428,dangling_wire_429}),
            .RCLKE(),
            .RCLK(N__32558),
            .RE(N__29650),
            .WCLKE(N__27347),
            .WCLK(N__32559),
            .WE(N__29510));
    defparam \this_sprites_ram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,\this_sprites_ram.mem_out_bus3_1 ,dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,dangling_wire_440,\this_sprites_ram.mem_out_bus3_0 ,dangling_wire_441,dangling_wire_442,dangling_wire_443}),
            .RADDR({N__30354,N__15534,N__15255,N__12126,N__26625,N__30198,N__31755,N__15678,N__14085,N__20841,N__19215}),
            .WADDR({N__25503,N__26373,N__27447,N__25653,N__25788,N__27138,N__24816,N__24960,N__25101,N__25236,N__26523}),
            .MASK({dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459}),
            .WDATA({dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,N__22092,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,N__24544,dangling_wire_471,dangling_wire_472,dangling_wire_473}),
            .RCLKE(),
            .RCLK(N__32578),
            .RE(N__29513),
            .WCLKE(N__27326),
            .WCLK(N__32579),
            .WE(N__29539));
    defparam \this_sprites_ram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,\this_sprites_ram.mem_out_bus3_3 ,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,dangling_wire_484,\this_sprites_ram.mem_out_bus3_2 ,dangling_wire_485,dangling_wire_486,dangling_wire_487}),
            .RADDR({N__30348,N__15528,N__15249,N__12120,N__26619,N__30192,N__31749,N__15672,N__14079,N__20835,N__19209}),
            .WADDR({N__25497,N__26367,N__27441,N__25647,N__25782,N__27132,N__24810,N__24954,N__25095,N__25230,N__26517}),
            .MASK({dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503}),
            .WDATA({dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,N__27763,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,dangling_wire_514,N__27204,dangling_wire_515,dangling_wire_516,dangling_wire_517}),
            .RCLKE(),
            .RCLK(N__32595),
            .RE(N__29512),
            .WCLKE(N__27327),
            .WCLK(N__32596),
            .WE(N__29426));
    defparam \this_sprites_ram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,\this_sprites_ram.mem_out_bus4_1 ,dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,dangling_wire_526,dangling_wire_527,dangling_wire_528,\this_sprites_ram.mem_out_bus4_0 ,dangling_wire_529,dangling_wire_530,dangling_wire_531}),
            .RADDR({N__30342,N__15522,N__15243,N__12114,N__26613,N__30186,N__31743,N__15666,N__14073,N__20829,N__19203}),
            .WADDR({N__25491,N__26361,N__27435,N__25641,N__25776,N__27126,N__24804,N__24948,N__25089,N__25224,N__26511}),
            .MASK({dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547}),
            .WDATA({dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,N__22093,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,dangling_wire_558,N__24553,dangling_wire_559,dangling_wire_560,dangling_wire_561}),
            .RCLKE(),
            .RCLK(N__32614),
            .RE(N__29514),
            .WCLKE(N__27035),
            .WCLK(N__32615),
            .WE(N__29519));
    defparam \this_sprites_ram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,\this_sprites_ram.mem_out_bus4_3 ,dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,dangling_wire_570,dangling_wire_571,dangling_wire_572,\this_sprites_ram.mem_out_bus4_2 ,dangling_wire_573,dangling_wire_574,dangling_wire_575}),
            .RADDR({N__30336,N__15516,N__15237,N__12108,N__26607,N__30180,N__31737,N__15660,N__14067,N__20823,N__19197}),
            .WADDR({N__25485,N__26355,N__27429,N__25635,N__25770,N__27120,N__24798,N__24942,N__25083,N__25218,N__26505}),
            .MASK({dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591}),
            .WDATA({dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,N__27772,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,dangling_wire_602,N__27237,dangling_wire_603,dangling_wire_604,dangling_wire_605}),
            .RCLKE(),
            .RCLK(N__32628),
            .RE(N__29515),
            .WCLKE(N__27042),
            .WCLK(N__32629),
            .WE(N__29520));
    defparam \this_sprites_ram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,\this_sprites_ram.mem_out_bus5_1 ,dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,dangling_wire_614,dangling_wire_615,dangling_wire_616,\this_sprites_ram.mem_out_bus5_0 ,dangling_wire_617,dangling_wire_618,dangling_wire_619}),
            .RADDR({N__30330,N__15510,N__15231,N__12102,N__26601,N__30174,N__31731,N__15654,N__14061,N__20817,N__19191}),
            .WADDR({N__25479,N__26349,N__27423,N__25629,N__25764,N__27114,N__24792,N__24936,N__25077,N__25212,N__26499}),
            .MASK({dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635}),
            .WDATA({dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,N__22111,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646,N__24569,dangling_wire_647,dangling_wire_648,dangling_wire_649}),
            .RCLKE(),
            .RCLK(N__32634),
            .RE(N__29702),
            .WCLKE(N__28571),
            .WCLK(N__32635),
            .WE(N__29629));
    defparam \this_sprites_ram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,\this_sprites_ram.mem_out_bus5_3 ,dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,dangling_wire_658,dangling_wire_659,dangling_wire_660,\this_sprites_ram.mem_out_bus5_2 ,dangling_wire_661,dangling_wire_662,dangling_wire_663}),
            .RADDR({N__30324,N__15504,N__15225,N__12096,N__26595,N__30168,N__31725,N__15648,N__14055,N__20811,N__19185}),
            .WADDR({N__25473,N__26343,N__27417,N__25623,N__25758,N__27108,N__24786,N__24930,N__25071,N__25206,N__26493}),
            .MASK({dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679}),
            .WDATA({dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,N__27788,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,N__27247,dangling_wire_691,dangling_wire_692,dangling_wire_693}),
            .RCLKE(),
            .RCLK(N__32645),
            .RE(N__29628),
            .WCLKE(N__28572),
            .WCLK(N__32646),
            .WE(N__29630));
    defparam \this_sprites_ram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,\this_sprites_ram.mem_out_bus6_1 ,dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,dangling_wire_702,dangling_wire_703,dangling_wire_704,\this_sprites_ram.mem_out_bus6_0 ,dangling_wire_705,dangling_wire_706,dangling_wire_707}),
            .RADDR({N__30318,N__15498,N__15219,N__12090,N__26589,N__30162,N__31719,N__15642,N__14049,N__20805,N__19179}),
            .WADDR({N__25467,N__26337,N__27411,N__25617,N__25752,N__27102,N__24780,N__24924,N__25065,N__25200,N__26487}),
            .MASK({dangling_wire_708,dangling_wire_709,dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,dangling_wire_723}),
            .WDATA({dangling_wire_724,dangling_wire_725,dangling_wire_726,dangling_wire_727,N__22125,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,N__24580,dangling_wire_735,dangling_wire_736,dangling_wire_737}),
            .RCLKE(),
            .RCLK(N__32652),
            .RE(N__29754),
            .WCLKE(N__30785),
            .WCLK(N__32653),
            .WE(N__29720));
    defparam \this_sprites_ram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741,\this_sprites_ram.mem_out_bus6_3 ,dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,dangling_wire_746,dangling_wire_747,dangling_wire_748,\this_sprites_ram.mem_out_bus6_2 ,dangling_wire_749,dangling_wire_750,dangling_wire_751}),
            .RADDR({N__30312,N__15492,N__15213,N__12084,N__26583,N__30156,N__31713,N__15636,N__14043,N__20799,N__19173}),
            .WADDR({N__25461,N__26331,N__27405,N__25611,N__25746,N__27096,N__24774,N__24918,N__25059,N__25194,N__26481}),
            .MASK({dangling_wire_752,dangling_wire_753,dangling_wire_754,dangling_wire_755,dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,dangling_wire_767}),
            .WDATA({dangling_wire_768,dangling_wire_769,dangling_wire_770,dangling_wire_771,N__27799,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,dangling_wire_778,N__27254,dangling_wire_779,dangling_wire_780,dangling_wire_781}),
            .RCLKE(),
            .RCLK(N__32657),
            .RE(N__29725),
            .WCLKE(N__30786),
            .WCLK(N__32658),
            .WE(N__29721));
    defparam \this_sprites_ram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785,\this_sprites_ram.mem_out_bus7_1 ,dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,dangling_wire_790,dangling_wire_791,dangling_wire_792,\this_sprites_ram.mem_out_bus7_0 ,dangling_wire_793,dangling_wire_794,dangling_wire_795}),
            .RADDR({N__30306,N__15486,N__15207,N__12078,N__26577,N__30150,N__31707,N__15630,N__14037,N__20793,N__19167}),
            .WADDR({N__25455,N__26325,N__27399,N__25605,N__25740,N__27090,N__24768,N__24912,N__25053,N__25188,N__26475}),
            .MASK({dangling_wire_796,dangling_wire_797,dangling_wire_798,dangling_wire_799,dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,dangling_wire_811}),
            .WDATA({dangling_wire_812,dangling_wire_813,dangling_wire_814,dangling_wire_815,N__22133,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,dangling_wire_822,N__24585,dangling_wire_823,dangling_wire_824,dangling_wire_825}),
            .RCLKE(),
            .RCLK(N__32661),
            .RE(N__29779),
            .WCLKE(N__30446),
            .WCLK(N__32662),
            .WE(N__29778));
    defparam \this_sprites_ram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829,\this_sprites_ram.mem_out_bus7_3 ,dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,dangling_wire_834,dangling_wire_835,dangling_wire_836,\this_sprites_ram.mem_out_bus7_2 ,dangling_wire_837,dangling_wire_838,dangling_wire_839}),
            .RADDR({N__30300,N__15480,N__15201,N__12072,N__26571,N__30144,N__31701,N__15624,N__14031,N__20787,N__19161}),
            .WADDR({N__25449,N__26319,N__27393,N__25599,N__25734,N__27084,N__24762,N__24906,N__25047,N__25182,N__26469}),
            .MASK({dangling_wire_840,dangling_wire_841,dangling_wire_842,dangling_wire_843,dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,dangling_wire_855}),
            .WDATA({dangling_wire_856,dangling_wire_857,dangling_wire_858,dangling_wire_859,N__27804,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,N__27258,dangling_wire_867,dangling_wire_868,dangling_wire_869}),
            .RCLKE(),
            .RCLK(N__32663),
            .RE(N__29780),
            .WCLKE(N__30447),
            .WCLK(N__32664),
            .WE(N__29812));
    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_870,dangling_wire_871,dangling_wire_872,dangling_wire_873,dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,M_this_vram_read_data_3,M_this_vram_read_data_2,M_this_vram_read_data_1,M_this_vram_read_data_0}),
            .RADDR({dangling_wire_882,dangling_wire_883,dangling_wire_884,N__17046,N__13323,N__11820,N__12195,N__13344,N__11805,N__11463,N__13197}),
            .WADDR({dangling_wire_885,dangling_wire_886,dangling_wire_887,N__16848,N__13623,N__13577,N__13820,N__13952,N__13890,N__20940,N__19335}),
            .MASK({dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,dangling_wire_899,dangling_wire_900,dangling_wire_901,dangling_wire_902,dangling_wire_903}),
            .WDATA({dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,dangling_wire_910,dangling_wire_911,dangling_wire_912,dangling_wire_913,dangling_wire_914,dangling_wire_915,N__28790,N__17190,N__21162,N__14685}),
            .RCLKE(),
            .RCLK(N__32659),
            .RE(N__29842),
            .WCLKE(N__14010),
            .WCLK(N__32660),
            .WE(N__29844));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__33433),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__33435),
            .DIN(N__33434),
            .DOUT(N__33433),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__33435),
            .PADOUT(N__33434),
            .PADIN(N__33433),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__33424),
            .DIN(N__33423),
            .DOUT(N__33422),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__33424),
            .PADOUT(N__33423),
            .PADIN(N__33422),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__33415),
            .DIN(N__33414),
            .DOUT(N__33413),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__33415),
            .PADOUT(N__33414),
            .PADIN(N__33413),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__33406),
            .DIN(N__33405),
            .DOUT(N__33404),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__33406),
            .PADOUT(N__33405),
            .PADIN(N__33404),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13224),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__33397),
            .DIN(N__33396),
            .DOUT(N__33395),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__33397),
            .PADOUT(N__33396),
            .PADIN(N__33395),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13443),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_0_iopad (
            .OE(N__33388),
            .DIN(N__33387),
            .DOUT(N__33386),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__33388),
            .PADOUT(N__33387),
            .PADIN(N__33386),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29835),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_1_iopad (
            .OE(N__33379),
            .DIN(N__33378),
            .DOUT(N__33377),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__33379),
            .PADOUT(N__33378),
            .PADIN(N__33377),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__19953),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_2_iopad (
            .OE(N__33370),
            .DIN(N__33369),
            .DOUT(N__33368),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__33370),
            .PADOUT(N__33369),
            .PADIN(N__33368),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_3_iopad (
            .OE(N__33361),
            .DIN(N__33360),
            .DOUT(N__33359),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__33361),
            .PADOUT(N__33360),
            .PADIN(N__33359),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_4_iopad (
            .OE(N__33352),
            .DIN(N__33351),
            .DOUT(N__33350),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__33352),
            .PADOUT(N__33351),
            .PADIN(N__33350),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_5_iopad (
            .OE(N__33343),
            .DIN(N__33342),
            .DOUT(N__33341),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__33343),
            .PADOUT(N__33342),
            .PADIN(N__33341),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_6_iopad (
            .OE(N__33334),
            .DIN(N__33333),
            .DOUT(N__33332),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__33334),
            .PADOUT(N__33333),
            .PADIN(N__33332),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_7_iopad (
            .OE(N__33325),
            .DIN(N__33324),
            .DOUT(N__33323),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__33325),
            .PADOUT(N__33324),
            .PADIN(N__33323),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__33316),
            .DIN(N__33315),
            .DOUT(N__33314),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__33316),
            .PADOUT(N__33315),
            .PADIN(N__33314),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__31191),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16079));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__33307),
            .DIN(N__33306),
            .DOUT(N__33305),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__33307),
            .PADOUT(N__33306),
            .PADIN(N__33305),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__31164),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16048));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__33298),
            .DIN(N__33297),
            .DOUT(N__33296),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__33298),
            .PADOUT(N__33297),
            .PADIN(N__33296),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__31143),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16113));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__33289),
            .DIN(N__33288),
            .DOUT(N__33287),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__33289),
            .PADOUT(N__33288),
            .PADIN(N__33287),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__31116),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16049));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__33280),
            .DIN(N__33279),
            .DOUT(N__33278),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__33280),
            .PADOUT(N__33279),
            .PADIN(N__33278),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__31089),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16122));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__33271),
            .DIN(N__33270),
            .DOUT(N__33269),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__33271),
            .PADOUT(N__33270),
            .PADIN(N__33269),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__31071),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16120));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__33262),
            .DIN(N__33261),
            .DOUT(N__33260),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__33262),
            .PADOUT(N__33261),
            .PADIN(N__33260),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__31047),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16091));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__33253),
            .DIN(N__33252),
            .DOUT(N__33251),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__33253),
            .PADOUT(N__33252),
            .PADIN(N__33251),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__31026),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16136));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__33244),
            .DIN(N__33243),
            .DOUT(N__33242),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__33244),
            .PADOUT(N__33243),
            .PADIN(N__33242),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__32682),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16112));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__33235),
            .DIN(N__33234),
            .DOUT(N__33233),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__33235),
            .PADOUT(N__33234),
            .PADIN(N__33233),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__31212),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16137));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__33226),
            .DIN(N__33225),
            .DOUT(N__33224),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__33226),
            .PADOUT(N__33225),
            .PADIN(N__33224),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__31542),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16123));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__33217),
            .DIN(N__33216),
            .DOUT(N__33215),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__33217),
            .PADOUT(N__33216),
            .PADIN(N__33215),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__31500),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16121));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__33208),
            .DIN(N__33207),
            .DOUT(N__33206),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__33208),
            .PADOUT(N__33207),
            .PADIN(N__33206),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__31452),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16015));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__33199),
            .DIN(N__33198),
            .DOUT(N__33197),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__33199),
            .PADOUT(N__33198),
            .PADIN(N__33197),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__31404),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16135));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__33190),
            .DIN(N__33189),
            .DOUT(N__33188),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__33190),
            .PADOUT(N__33189),
            .PADIN(N__33188),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__30996),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16011));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__33181),
            .DIN(N__33180),
            .DOUT(N__33179),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__33181),
            .PADOUT(N__33180),
            .PADIN(N__33179),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__31584),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16131));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__33172),
            .DIN(N__33171),
            .DOUT(N__33170),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__33172),
            .PADOUT(N__33171),
            .PADIN(N__33170),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__33163),
            .DIN(N__33162),
            .DOUT(N__33161),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__33163),
            .PADOUT(N__33162),
            .PADIN(N__33161),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__33154),
            .DIN(N__33153),
            .DOUT(N__33152),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__33154),
            .PADOUT(N__33153),
            .PADIN(N__33152),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__33145),
            .DIN(N__33144),
            .DOUT(N__33143),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__33145),
            .PADOUT(N__33144),
            .PADIN(N__33143),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__33136),
            .DIN(N__33135),
            .DOUT(N__33134),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__33136),
            .PADOUT(N__33135),
            .PADIN(N__33134),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__33127),
            .DIN(N__33126),
            .DOUT(N__33125),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__33127),
            .PADOUT(N__33126),
            .PADIN(N__33125),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__33118),
            .DIN(N__33117),
            .DOUT(N__33116),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__33118),
            .PADOUT(N__33117),
            .PADIN(N__33116),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__33109),
            .DIN(N__33108),
            .DOUT(N__33107),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__33109),
            .PADOUT(N__33108),
            .PADIN(N__33107),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_7_iopad (
            .OE(N__33100),
            .DIN(N__33099),
            .DOUT(N__33098),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_7_preio (
            .PADOEN(N__33100),
            .PADOUT(N__33099),
            .PADIN(N__33098),
            .CLOCKENABLE(),
            .DIN0(port_data_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__33091),
            .DIN(N__33090),
            .DOUT(N__33089),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__33091),
            .PADOUT(N__33090),
            .PADIN(N__33089),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__17298),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__33082),
            .DIN(N__33081),
            .DOUT(N__33080),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__33082),
            .PADOUT(N__33081),
            .PADIN(N__33080),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__17745),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__33073),
            .DIN(N__33072),
            .DOUT(N__33071),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__33073),
            .PADOUT(N__33072),
            .PADIN(N__33071),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__33064),
            .DIN(N__33063),
            .DOUT(N__33062),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__33064),
            .PADOUT(N__33063),
            .PADIN(N__33062),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__10980),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__33055),
            .DIN(N__33054),
            .DOUT(N__33053),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__33055),
            .PADOUT(N__33054),
            .PADIN(N__33053),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__29843),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16130));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__33046),
            .DIN(N__33045),
            .DOUT(N__33044),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__33046),
            .PADOUT(N__33045),
            .PADIN(N__33044),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11154),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__33037),
            .DIN(N__33036),
            .DOUT(N__33035),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__33037),
            .PADOUT(N__33036),
            .PADIN(N__33035),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11475),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__33028),
            .DIN(N__33027),
            .DOUT(N__33026),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__33028),
            .PADOUT(N__33027),
            .PADIN(N__33026),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11124),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__33019),
            .DIN(N__33018),
            .DOUT(N__33017),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__33019),
            .PADOUT(N__33018),
            .PADIN(N__33017),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11328),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__33010),
            .DIN(N__33009),
            .DOUT(N__33008),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__33010),
            .PADOUT(N__33009),
            .PADIN(N__33008),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11316),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__33001),
            .DIN(N__33000),
            .DOUT(N__32999),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__33001),
            .PADOUT(N__33000),
            .PADIN(N__32999),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11835),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__32992),
            .DIN(N__32991),
            .DOUT(N__32990),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__32992),
            .PADOUT(N__32991),
            .PADIN(N__32990),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__32983),
            .DIN(N__32982),
            .DOUT(N__32981),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__32983),
            .PADOUT(N__32982),
            .PADIN(N__32981),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11139),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__32974),
            .DIN(N__32973),
            .DOUT(N__32972),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__32974),
            .PADOUT(N__32973),
            .PADIN(N__32972),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22200),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__8133 (
            .O(N__32955),
            .I(N__32952));
    LocalMux I__8132 (
            .O(N__32952),
            .I(M_this_external_address_q_s_10));
    InMux I__8131 (
            .O(N__32949),
            .I(N__32945));
    InMux I__8130 (
            .O(N__32948),
            .I(N__32942));
    LocalMux I__8129 (
            .O(N__32945),
            .I(N__32936));
    LocalMux I__8128 (
            .O(N__32942),
            .I(N__32936));
    InMux I__8127 (
            .O(N__32941),
            .I(N__32933));
    Span4Mux_v I__8126 (
            .O(N__32936),
            .I(N__32927));
    LocalMux I__8125 (
            .O(N__32933),
            .I(N__32927));
    InMux I__8124 (
            .O(N__32932),
            .I(N__32924));
    Odrv4 I__8123 (
            .O(N__32927),
            .I(M_this_external_address_d_1_sqmuxa));
    LocalMux I__8122 (
            .O(N__32924),
            .I(M_this_external_address_d_1_sqmuxa));
    InMux I__8121 (
            .O(N__32919),
            .I(N__32916));
    LocalMux I__8120 (
            .O(N__32916),
            .I(N__32912));
    InMux I__8119 (
            .O(N__32915),
            .I(N__32909));
    Span4Mux_v I__8118 (
            .O(N__32912),
            .I(N__32905));
    LocalMux I__8117 (
            .O(N__32909),
            .I(N__32900));
    InMux I__8116 (
            .O(N__32908),
            .I(N__32897));
    Span4Mux_h I__8115 (
            .O(N__32905),
            .I(N__32893));
    InMux I__8114 (
            .O(N__32904),
            .I(N__32888));
    CascadeMux I__8113 (
            .O(N__32903),
            .I(N__32885));
    Span4Mux_h I__8112 (
            .O(N__32900),
            .I(N__32879));
    LocalMux I__8111 (
            .O(N__32897),
            .I(N__32879));
    InMux I__8110 (
            .O(N__32896),
            .I(N__32876));
    Span4Mux_h I__8109 (
            .O(N__32893),
            .I(N__32871));
    InMux I__8108 (
            .O(N__32892),
            .I(N__32868));
    InMux I__8107 (
            .O(N__32891),
            .I(N__32865));
    LocalMux I__8106 (
            .O(N__32888),
            .I(N__32862));
    InMux I__8105 (
            .O(N__32885),
            .I(N__32859));
    CascadeMux I__8104 (
            .O(N__32884),
            .I(N__32855));
    Span4Mux_v I__8103 (
            .O(N__32879),
            .I(N__32850));
    LocalMux I__8102 (
            .O(N__32876),
            .I(N__32850));
    InMux I__8101 (
            .O(N__32875),
            .I(N__32845));
    InMux I__8100 (
            .O(N__32874),
            .I(N__32845));
    Span4Mux_h I__8099 (
            .O(N__32871),
            .I(N__32840));
    LocalMux I__8098 (
            .O(N__32868),
            .I(N__32840));
    LocalMux I__8097 (
            .O(N__32865),
            .I(N__32833));
    Span4Mux_h I__8096 (
            .O(N__32862),
            .I(N__32833));
    LocalMux I__8095 (
            .O(N__32859),
            .I(N__32833));
    InMux I__8094 (
            .O(N__32858),
            .I(N__32830));
    InMux I__8093 (
            .O(N__32855),
            .I(N__32827));
    Span4Mux_v I__8092 (
            .O(N__32850),
            .I(N__32823));
    LocalMux I__8091 (
            .O(N__32845),
            .I(N__32820));
    Span4Mux_h I__8090 (
            .O(N__32840),
            .I(N__32810));
    Span4Mux_v I__8089 (
            .O(N__32833),
            .I(N__32810));
    LocalMux I__8088 (
            .O(N__32830),
            .I(N__32810));
    LocalMux I__8087 (
            .O(N__32827),
            .I(N__32810));
    InMux I__8086 (
            .O(N__32826),
            .I(N__32807));
    Span4Mux_h I__8085 (
            .O(N__32823),
            .I(N__32804));
    Span4Mux_v I__8084 (
            .O(N__32820),
            .I(N__32801));
    CascadeMux I__8083 (
            .O(N__32819),
            .I(N__32797));
    Span4Mux_v I__8082 (
            .O(N__32810),
            .I(N__32794));
    LocalMux I__8081 (
            .O(N__32807),
            .I(N__32791));
    Span4Mux_h I__8080 (
            .O(N__32804),
            .I(N__32786));
    Span4Mux_v I__8079 (
            .O(N__32801),
            .I(N__32786));
    InMux I__8078 (
            .O(N__32800),
            .I(N__32783));
    InMux I__8077 (
            .O(N__32797),
            .I(N__32780));
    Span4Mux_h I__8076 (
            .O(N__32794),
            .I(N__32777));
    Span12Mux_v I__8075 (
            .O(N__32791),
            .I(N__32768));
    Sp12to4 I__8074 (
            .O(N__32786),
            .I(N__32768));
    LocalMux I__8073 (
            .O(N__32783),
            .I(N__32768));
    LocalMux I__8072 (
            .O(N__32780),
            .I(N__32768));
    Sp12to4 I__8071 (
            .O(N__32777),
            .I(N__32763));
    Span12Mux_h I__8070 (
            .O(N__32768),
            .I(N__32763));
    Odrv12 I__8069 (
            .O(N__32763),
            .I(port_data_c_2));
    InMux I__8068 (
            .O(N__32760),
            .I(N__32741));
    InMux I__8067 (
            .O(N__32759),
            .I(N__32741));
    InMux I__8066 (
            .O(N__32758),
            .I(N__32741));
    InMux I__8065 (
            .O(N__32757),
            .I(N__32736));
    InMux I__8064 (
            .O(N__32756),
            .I(N__32736));
    InMux I__8063 (
            .O(N__32755),
            .I(N__32724));
    InMux I__8062 (
            .O(N__32754),
            .I(N__32724));
    InMux I__8061 (
            .O(N__32753),
            .I(N__32724));
    InMux I__8060 (
            .O(N__32752),
            .I(N__32724));
    InMux I__8059 (
            .O(N__32751),
            .I(N__32715));
    InMux I__8058 (
            .O(N__32750),
            .I(N__32715));
    InMux I__8057 (
            .O(N__32749),
            .I(N__32715));
    InMux I__8056 (
            .O(N__32748),
            .I(N__32715));
    LocalMux I__8055 (
            .O(N__32741),
            .I(N__32712));
    LocalMux I__8054 (
            .O(N__32736),
            .I(N__32709));
    InMux I__8053 (
            .O(N__32735),
            .I(N__32702));
    InMux I__8052 (
            .O(N__32734),
            .I(N__32702));
    InMux I__8051 (
            .O(N__32733),
            .I(N__32702));
    LocalMux I__8050 (
            .O(N__32724),
            .I(N__32697));
    LocalMux I__8049 (
            .O(N__32715),
            .I(N__32697));
    Span4Mux_h I__8048 (
            .O(N__32712),
            .I(N__32694));
    Span4Mux_h I__8047 (
            .O(N__32709),
            .I(N__32691));
    LocalMux I__8046 (
            .O(N__32702),
            .I(N_39));
    Odrv12 I__8045 (
            .O(N__32697),
            .I(N_39));
    Odrv4 I__8044 (
            .O(N__32694),
            .I(N_39));
    Odrv4 I__8043 (
            .O(N__32691),
            .I(N_39));
    IoInMux I__8042 (
            .O(N__32682),
            .I(N__32679));
    LocalMux I__8041 (
            .O(N__32679),
            .I(N__32676));
    Span12Mux_s7_v I__8040 (
            .O(N__32676),
            .I(N__32672));
    InMux I__8039 (
            .O(N__32675),
            .I(N__32669));
    Odrv12 I__8038 (
            .O(N__32672),
            .I(M_this_external_address_qZ0Z_10));
    LocalMux I__8037 (
            .O(N__32669),
            .I(M_this_external_address_qZ0Z_10));
    ClkMux I__8036 (
            .O(N__32664),
            .I(N__32241));
    ClkMux I__8035 (
            .O(N__32663),
            .I(N__32241));
    ClkMux I__8034 (
            .O(N__32662),
            .I(N__32241));
    ClkMux I__8033 (
            .O(N__32661),
            .I(N__32241));
    ClkMux I__8032 (
            .O(N__32660),
            .I(N__32241));
    ClkMux I__8031 (
            .O(N__32659),
            .I(N__32241));
    ClkMux I__8030 (
            .O(N__32658),
            .I(N__32241));
    ClkMux I__8029 (
            .O(N__32657),
            .I(N__32241));
    ClkMux I__8028 (
            .O(N__32656),
            .I(N__32241));
    ClkMux I__8027 (
            .O(N__32655),
            .I(N__32241));
    ClkMux I__8026 (
            .O(N__32654),
            .I(N__32241));
    ClkMux I__8025 (
            .O(N__32653),
            .I(N__32241));
    ClkMux I__8024 (
            .O(N__32652),
            .I(N__32241));
    ClkMux I__8023 (
            .O(N__32651),
            .I(N__32241));
    ClkMux I__8022 (
            .O(N__32650),
            .I(N__32241));
    ClkMux I__8021 (
            .O(N__32649),
            .I(N__32241));
    ClkMux I__8020 (
            .O(N__32648),
            .I(N__32241));
    ClkMux I__8019 (
            .O(N__32647),
            .I(N__32241));
    ClkMux I__8018 (
            .O(N__32646),
            .I(N__32241));
    ClkMux I__8017 (
            .O(N__32645),
            .I(N__32241));
    ClkMux I__8016 (
            .O(N__32644),
            .I(N__32241));
    ClkMux I__8015 (
            .O(N__32643),
            .I(N__32241));
    ClkMux I__8014 (
            .O(N__32642),
            .I(N__32241));
    ClkMux I__8013 (
            .O(N__32641),
            .I(N__32241));
    ClkMux I__8012 (
            .O(N__32640),
            .I(N__32241));
    ClkMux I__8011 (
            .O(N__32639),
            .I(N__32241));
    ClkMux I__8010 (
            .O(N__32638),
            .I(N__32241));
    ClkMux I__8009 (
            .O(N__32637),
            .I(N__32241));
    ClkMux I__8008 (
            .O(N__32636),
            .I(N__32241));
    ClkMux I__8007 (
            .O(N__32635),
            .I(N__32241));
    ClkMux I__8006 (
            .O(N__32634),
            .I(N__32241));
    ClkMux I__8005 (
            .O(N__32633),
            .I(N__32241));
    ClkMux I__8004 (
            .O(N__32632),
            .I(N__32241));
    ClkMux I__8003 (
            .O(N__32631),
            .I(N__32241));
    ClkMux I__8002 (
            .O(N__32630),
            .I(N__32241));
    ClkMux I__8001 (
            .O(N__32629),
            .I(N__32241));
    ClkMux I__8000 (
            .O(N__32628),
            .I(N__32241));
    ClkMux I__7999 (
            .O(N__32627),
            .I(N__32241));
    ClkMux I__7998 (
            .O(N__32626),
            .I(N__32241));
    ClkMux I__7997 (
            .O(N__32625),
            .I(N__32241));
    ClkMux I__7996 (
            .O(N__32624),
            .I(N__32241));
    ClkMux I__7995 (
            .O(N__32623),
            .I(N__32241));
    ClkMux I__7994 (
            .O(N__32622),
            .I(N__32241));
    ClkMux I__7993 (
            .O(N__32621),
            .I(N__32241));
    ClkMux I__7992 (
            .O(N__32620),
            .I(N__32241));
    ClkMux I__7991 (
            .O(N__32619),
            .I(N__32241));
    ClkMux I__7990 (
            .O(N__32618),
            .I(N__32241));
    ClkMux I__7989 (
            .O(N__32617),
            .I(N__32241));
    ClkMux I__7988 (
            .O(N__32616),
            .I(N__32241));
    ClkMux I__7987 (
            .O(N__32615),
            .I(N__32241));
    ClkMux I__7986 (
            .O(N__32614),
            .I(N__32241));
    ClkMux I__7985 (
            .O(N__32613),
            .I(N__32241));
    ClkMux I__7984 (
            .O(N__32612),
            .I(N__32241));
    ClkMux I__7983 (
            .O(N__32611),
            .I(N__32241));
    ClkMux I__7982 (
            .O(N__32610),
            .I(N__32241));
    ClkMux I__7981 (
            .O(N__32609),
            .I(N__32241));
    ClkMux I__7980 (
            .O(N__32608),
            .I(N__32241));
    ClkMux I__7979 (
            .O(N__32607),
            .I(N__32241));
    ClkMux I__7978 (
            .O(N__32606),
            .I(N__32241));
    ClkMux I__7977 (
            .O(N__32605),
            .I(N__32241));
    ClkMux I__7976 (
            .O(N__32604),
            .I(N__32241));
    ClkMux I__7975 (
            .O(N__32603),
            .I(N__32241));
    ClkMux I__7974 (
            .O(N__32602),
            .I(N__32241));
    ClkMux I__7973 (
            .O(N__32601),
            .I(N__32241));
    ClkMux I__7972 (
            .O(N__32600),
            .I(N__32241));
    ClkMux I__7971 (
            .O(N__32599),
            .I(N__32241));
    ClkMux I__7970 (
            .O(N__32598),
            .I(N__32241));
    ClkMux I__7969 (
            .O(N__32597),
            .I(N__32241));
    ClkMux I__7968 (
            .O(N__32596),
            .I(N__32241));
    ClkMux I__7967 (
            .O(N__32595),
            .I(N__32241));
    ClkMux I__7966 (
            .O(N__32594),
            .I(N__32241));
    ClkMux I__7965 (
            .O(N__32593),
            .I(N__32241));
    ClkMux I__7964 (
            .O(N__32592),
            .I(N__32241));
    ClkMux I__7963 (
            .O(N__32591),
            .I(N__32241));
    ClkMux I__7962 (
            .O(N__32590),
            .I(N__32241));
    ClkMux I__7961 (
            .O(N__32589),
            .I(N__32241));
    ClkMux I__7960 (
            .O(N__32588),
            .I(N__32241));
    ClkMux I__7959 (
            .O(N__32587),
            .I(N__32241));
    ClkMux I__7958 (
            .O(N__32586),
            .I(N__32241));
    ClkMux I__7957 (
            .O(N__32585),
            .I(N__32241));
    ClkMux I__7956 (
            .O(N__32584),
            .I(N__32241));
    ClkMux I__7955 (
            .O(N__32583),
            .I(N__32241));
    ClkMux I__7954 (
            .O(N__32582),
            .I(N__32241));
    ClkMux I__7953 (
            .O(N__32581),
            .I(N__32241));
    ClkMux I__7952 (
            .O(N__32580),
            .I(N__32241));
    ClkMux I__7951 (
            .O(N__32579),
            .I(N__32241));
    ClkMux I__7950 (
            .O(N__32578),
            .I(N__32241));
    ClkMux I__7949 (
            .O(N__32577),
            .I(N__32241));
    ClkMux I__7948 (
            .O(N__32576),
            .I(N__32241));
    ClkMux I__7947 (
            .O(N__32575),
            .I(N__32241));
    ClkMux I__7946 (
            .O(N__32574),
            .I(N__32241));
    ClkMux I__7945 (
            .O(N__32573),
            .I(N__32241));
    ClkMux I__7944 (
            .O(N__32572),
            .I(N__32241));
    ClkMux I__7943 (
            .O(N__32571),
            .I(N__32241));
    ClkMux I__7942 (
            .O(N__32570),
            .I(N__32241));
    ClkMux I__7941 (
            .O(N__32569),
            .I(N__32241));
    ClkMux I__7940 (
            .O(N__32568),
            .I(N__32241));
    ClkMux I__7939 (
            .O(N__32567),
            .I(N__32241));
    ClkMux I__7938 (
            .O(N__32566),
            .I(N__32241));
    ClkMux I__7937 (
            .O(N__32565),
            .I(N__32241));
    ClkMux I__7936 (
            .O(N__32564),
            .I(N__32241));
    ClkMux I__7935 (
            .O(N__32563),
            .I(N__32241));
    ClkMux I__7934 (
            .O(N__32562),
            .I(N__32241));
    ClkMux I__7933 (
            .O(N__32561),
            .I(N__32241));
    ClkMux I__7932 (
            .O(N__32560),
            .I(N__32241));
    ClkMux I__7931 (
            .O(N__32559),
            .I(N__32241));
    ClkMux I__7930 (
            .O(N__32558),
            .I(N__32241));
    ClkMux I__7929 (
            .O(N__32557),
            .I(N__32241));
    ClkMux I__7928 (
            .O(N__32556),
            .I(N__32241));
    ClkMux I__7927 (
            .O(N__32555),
            .I(N__32241));
    ClkMux I__7926 (
            .O(N__32554),
            .I(N__32241));
    ClkMux I__7925 (
            .O(N__32553),
            .I(N__32241));
    ClkMux I__7924 (
            .O(N__32552),
            .I(N__32241));
    ClkMux I__7923 (
            .O(N__32551),
            .I(N__32241));
    ClkMux I__7922 (
            .O(N__32550),
            .I(N__32241));
    ClkMux I__7921 (
            .O(N__32549),
            .I(N__32241));
    ClkMux I__7920 (
            .O(N__32548),
            .I(N__32241));
    ClkMux I__7919 (
            .O(N__32547),
            .I(N__32241));
    ClkMux I__7918 (
            .O(N__32546),
            .I(N__32241));
    ClkMux I__7917 (
            .O(N__32545),
            .I(N__32241));
    ClkMux I__7916 (
            .O(N__32544),
            .I(N__32241));
    ClkMux I__7915 (
            .O(N__32543),
            .I(N__32241));
    ClkMux I__7914 (
            .O(N__32542),
            .I(N__32241));
    ClkMux I__7913 (
            .O(N__32541),
            .I(N__32241));
    ClkMux I__7912 (
            .O(N__32540),
            .I(N__32241));
    ClkMux I__7911 (
            .O(N__32539),
            .I(N__32241));
    ClkMux I__7910 (
            .O(N__32538),
            .I(N__32241));
    ClkMux I__7909 (
            .O(N__32537),
            .I(N__32241));
    ClkMux I__7908 (
            .O(N__32536),
            .I(N__32241));
    ClkMux I__7907 (
            .O(N__32535),
            .I(N__32241));
    ClkMux I__7906 (
            .O(N__32534),
            .I(N__32241));
    ClkMux I__7905 (
            .O(N__32533),
            .I(N__32241));
    ClkMux I__7904 (
            .O(N__32532),
            .I(N__32241));
    ClkMux I__7903 (
            .O(N__32531),
            .I(N__32241));
    ClkMux I__7902 (
            .O(N__32530),
            .I(N__32241));
    ClkMux I__7901 (
            .O(N__32529),
            .I(N__32241));
    ClkMux I__7900 (
            .O(N__32528),
            .I(N__32241));
    ClkMux I__7899 (
            .O(N__32527),
            .I(N__32241));
    ClkMux I__7898 (
            .O(N__32526),
            .I(N__32241));
    ClkMux I__7897 (
            .O(N__32525),
            .I(N__32241));
    ClkMux I__7896 (
            .O(N__32524),
            .I(N__32241));
    GlobalMux I__7895 (
            .O(N__32241),
            .I(N__32238));
    gio2CtrlBuf I__7894 (
            .O(N__32238),
            .I(clk_0_c_g));
    CEMux I__7893 (
            .O(N__32235),
            .I(N__32230));
    CEMux I__7892 (
            .O(N__32234),
            .I(N__32227));
    CEMux I__7891 (
            .O(N__32233),
            .I(N__32224));
    LocalMux I__7890 (
            .O(N__32230),
            .I(N__32221));
    LocalMux I__7889 (
            .O(N__32227),
            .I(N__32217));
    LocalMux I__7888 (
            .O(N__32224),
            .I(N__32214));
    Span4Mux_h I__7887 (
            .O(N__32221),
            .I(N__32211));
    CEMux I__7886 (
            .O(N__32220),
            .I(N__32208));
    Span4Mux_h I__7885 (
            .O(N__32217),
            .I(N__32205));
    Span4Mux_h I__7884 (
            .O(N__32214),
            .I(N__32202));
    Span4Mux_h I__7883 (
            .O(N__32211),
            .I(N__32199));
    LocalMux I__7882 (
            .O(N__32208),
            .I(N__32196));
    Odrv4 I__7881 (
            .O(N__32205),
            .I(N_37));
    Odrv4 I__7880 (
            .O(N__32202),
            .I(N_37));
    Odrv4 I__7879 (
            .O(N__32199),
            .I(N_37));
    Odrv4 I__7878 (
            .O(N__32196),
            .I(N_37));
    InMux I__7877 (
            .O(N__32187),
            .I(N__32184));
    LocalMux I__7876 (
            .O(N__32184),
            .I(N__32181));
    Span4Mux_h I__7875 (
            .O(N__32181),
            .I(N__32178));
    Sp12to4 I__7874 (
            .O(N__32178),
            .I(N__32171));
    InMux I__7873 (
            .O(N__32177),
            .I(N__32168));
    CascadeMux I__7872 (
            .O(N__32176),
            .I(N__32165));
    InMux I__7871 (
            .O(N__32175),
            .I(N__32160));
    InMux I__7870 (
            .O(N__32174),
            .I(N__32160));
    Span12Mux_v I__7869 (
            .O(N__32171),
            .I(N__32157));
    LocalMux I__7868 (
            .O(N__32168),
            .I(N__32154));
    InMux I__7867 (
            .O(N__32165),
            .I(N__32151));
    LocalMux I__7866 (
            .O(N__32160),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv12 I__7865 (
            .O(N__32157),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv4 I__7864 (
            .O(N__32154),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    LocalMux I__7863 (
            .O(N__32151),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    InMux I__7862 (
            .O(N__32142),
            .I(N__32137));
    InMux I__7861 (
            .O(N__32141),
            .I(N__32125));
    InMux I__7860 (
            .O(N__32140),
            .I(N__32120));
    LocalMux I__7859 (
            .O(N__32137),
            .I(N__32116));
    InMux I__7858 (
            .O(N__32136),
            .I(N__32113));
    InMux I__7857 (
            .O(N__32135),
            .I(N__32106));
    InMux I__7856 (
            .O(N__32134),
            .I(N__32106));
    InMux I__7855 (
            .O(N__32133),
            .I(N__32106));
    InMux I__7854 (
            .O(N__32132),
            .I(N__32103));
    InMux I__7853 (
            .O(N__32131),
            .I(N__32099));
    InMux I__7852 (
            .O(N__32130),
            .I(N__32096));
    InMux I__7851 (
            .O(N__32129),
            .I(N__32091));
    InMux I__7850 (
            .O(N__32128),
            .I(N__32091));
    LocalMux I__7849 (
            .O(N__32125),
            .I(N__32088));
    InMux I__7848 (
            .O(N__32124),
            .I(N__32085));
    InMux I__7847 (
            .O(N__32123),
            .I(N__32082));
    LocalMux I__7846 (
            .O(N__32120),
            .I(N__32079));
    InMux I__7845 (
            .O(N__32119),
            .I(N__32072));
    Span4Mux_h I__7844 (
            .O(N__32116),
            .I(N__32063));
    LocalMux I__7843 (
            .O(N__32113),
            .I(N__32063));
    LocalMux I__7842 (
            .O(N__32106),
            .I(N__32063));
    LocalMux I__7841 (
            .O(N__32103),
            .I(N__32063));
    InMux I__7840 (
            .O(N__32102),
            .I(N__32060));
    LocalMux I__7839 (
            .O(N__32099),
            .I(N__32053));
    LocalMux I__7838 (
            .O(N__32096),
            .I(N__32053));
    LocalMux I__7837 (
            .O(N__32091),
            .I(N__32053));
    Span4Mux_h I__7836 (
            .O(N__32088),
            .I(N__32048));
    LocalMux I__7835 (
            .O(N__32085),
            .I(N__32048));
    LocalMux I__7834 (
            .O(N__32082),
            .I(N__32045));
    Span4Mux_h I__7833 (
            .O(N__32079),
            .I(N__32042));
    InMux I__7832 (
            .O(N__32078),
            .I(N__32035));
    InMux I__7831 (
            .O(N__32077),
            .I(N__32035));
    InMux I__7830 (
            .O(N__32076),
            .I(N__32035));
    InMux I__7829 (
            .O(N__32075),
            .I(N__32032));
    LocalMux I__7828 (
            .O(N__32072),
            .I(N__32029));
    Span4Mux_v I__7827 (
            .O(N__32063),
            .I(N__32026));
    LocalMux I__7826 (
            .O(N__32060),
            .I(N__32021));
    Span4Mux_h I__7825 (
            .O(N__32053),
            .I(N__32021));
    Span4Mux_h I__7824 (
            .O(N__32048),
            .I(N__32016));
    Span4Mux_h I__7823 (
            .O(N__32045),
            .I(N__32016));
    Sp12to4 I__7822 (
            .O(N__32042),
            .I(N__32011));
    LocalMux I__7821 (
            .O(N__32035),
            .I(N__32011));
    LocalMux I__7820 (
            .O(N__32032),
            .I(N__32008));
    Span4Mux_s2_v I__7819 (
            .O(N__32029),
            .I(N__32005));
    Span4Mux_v I__7818 (
            .O(N__32026),
            .I(N__32002));
    Span4Mux_h I__7817 (
            .O(N__32021),
            .I(N__31999));
    Span4Mux_v I__7816 (
            .O(N__32016),
            .I(N__31996));
    Span12Mux_v I__7815 (
            .O(N__32011),
            .I(N__31993));
    Span4Mux_s2_v I__7814 (
            .O(N__32008),
            .I(N__31990));
    Span4Mux_h I__7813 (
            .O(N__32005),
            .I(N__31985));
    Span4Mux_v I__7812 (
            .O(N__32002),
            .I(N__31985));
    Span4Mux_h I__7811 (
            .O(N__31999),
            .I(N__31980));
    Span4Mux_v I__7810 (
            .O(N__31996),
            .I(N__31980));
    Odrv12 I__7809 (
            .O(N__31993),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__7808 (
            .O(N__31990),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__7807 (
            .O(N__31985),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__7806 (
            .O(N__31980),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    CascadeMux I__7805 (
            .O(N__31971),
            .I(N__31966));
    CascadeMux I__7804 (
            .O(N__31970),
            .I(N__31961));
    CascadeMux I__7803 (
            .O(N__31969),
            .I(N__31957));
    InMux I__7802 (
            .O(N__31966),
            .I(N__31954));
    InMux I__7801 (
            .O(N__31965),
            .I(N__31951));
    CascadeMux I__7800 (
            .O(N__31964),
            .I(N__31948));
    InMux I__7799 (
            .O(N__31961),
            .I(N__31945));
    InMux I__7798 (
            .O(N__31960),
            .I(N__31940));
    InMux I__7797 (
            .O(N__31957),
            .I(N__31940));
    LocalMux I__7796 (
            .O(N__31954),
            .I(N__31936));
    LocalMux I__7795 (
            .O(N__31951),
            .I(N__31931));
    InMux I__7794 (
            .O(N__31948),
            .I(N__31928));
    LocalMux I__7793 (
            .O(N__31945),
            .I(N__31923));
    LocalMux I__7792 (
            .O(N__31940),
            .I(N__31923));
    CascadeMux I__7791 (
            .O(N__31939),
            .I(N__31920));
    Span4Mux_v I__7790 (
            .O(N__31936),
            .I(N__31916));
    CascadeMux I__7789 (
            .O(N__31935),
            .I(N__31913));
    CascadeMux I__7788 (
            .O(N__31934),
            .I(N__31909));
    Span4Mux_v I__7787 (
            .O(N__31931),
            .I(N__31906));
    LocalMux I__7786 (
            .O(N__31928),
            .I(N__31901));
    Span4Mux_h I__7785 (
            .O(N__31923),
            .I(N__31901));
    InMux I__7784 (
            .O(N__31920),
            .I(N__31898));
    InMux I__7783 (
            .O(N__31919),
            .I(N__31895));
    Span4Mux_v I__7782 (
            .O(N__31916),
            .I(N__31892));
    InMux I__7781 (
            .O(N__31913),
            .I(N__31889));
    CascadeMux I__7780 (
            .O(N__31912),
            .I(N__31886));
    InMux I__7779 (
            .O(N__31909),
            .I(N__31879));
    Span4Mux_h I__7778 (
            .O(N__31906),
            .I(N__31872));
    Span4Mux_h I__7777 (
            .O(N__31901),
            .I(N__31872));
    LocalMux I__7776 (
            .O(N__31898),
            .I(N__31872));
    LocalMux I__7775 (
            .O(N__31895),
            .I(N__31869));
    Span4Mux_v I__7774 (
            .O(N__31892),
            .I(N__31864));
    LocalMux I__7773 (
            .O(N__31889),
            .I(N__31864));
    InMux I__7772 (
            .O(N__31886),
            .I(N__31857));
    InMux I__7771 (
            .O(N__31885),
            .I(N__31857));
    InMux I__7770 (
            .O(N__31884),
            .I(N__31857));
    InMux I__7769 (
            .O(N__31883),
            .I(N__31853));
    CascadeMux I__7768 (
            .O(N__31882),
            .I(N__31850));
    LocalMux I__7767 (
            .O(N__31879),
            .I(N__31845));
    Sp12to4 I__7766 (
            .O(N__31872),
            .I(N__31845));
    Span4Mux_h I__7765 (
            .O(N__31869),
            .I(N__31842));
    Span4Mux_h I__7764 (
            .O(N__31864),
            .I(N__31837));
    LocalMux I__7763 (
            .O(N__31857),
            .I(N__31837));
    InMux I__7762 (
            .O(N__31856),
            .I(N__31834));
    LocalMux I__7761 (
            .O(N__31853),
            .I(N__31831));
    InMux I__7760 (
            .O(N__31850),
            .I(N__31828));
    Span12Mux_v I__7759 (
            .O(N__31845),
            .I(N__31825));
    Span4Mux_h I__7758 (
            .O(N__31842),
            .I(N__31820));
    Span4Mux_h I__7757 (
            .O(N__31837),
            .I(N__31820));
    LocalMux I__7756 (
            .O(N__31834),
            .I(N__31815));
    Span4Mux_h I__7755 (
            .O(N__31831),
            .I(N__31815));
    LocalMux I__7754 (
            .O(N__31828),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    Odrv12 I__7753 (
            .O(N__31825),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    Odrv4 I__7752 (
            .O(N__31820),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    Odrv4 I__7751 (
            .O(N__31815),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    InMux I__7750 (
            .O(N__31806),
            .I(N__31803));
    LocalMux I__7749 (
            .O(N__31803),
            .I(N__31800));
    Span12Mux_s11_h I__7748 (
            .O(N__31800),
            .I(N__31797));
    Span12Mux_v I__7747 (
            .O(N__31797),
            .I(N__31794));
    Odrv12 I__7746 (
            .O(N__31794),
            .I(\this_ppu.un3_sprites_addr_cry_3_c_RNI1VDZ0Z8 ));
    CascadeMux I__7745 (
            .O(N__31791),
            .I(N__31788));
    CascadeBuf I__7744 (
            .O(N__31788),
            .I(N__31785));
    CascadeMux I__7743 (
            .O(N__31785),
            .I(N__31782));
    CascadeBuf I__7742 (
            .O(N__31782),
            .I(N__31779));
    CascadeMux I__7741 (
            .O(N__31779),
            .I(N__31776));
    CascadeBuf I__7740 (
            .O(N__31776),
            .I(N__31773));
    CascadeMux I__7739 (
            .O(N__31773),
            .I(N__31770));
    CascadeBuf I__7738 (
            .O(N__31770),
            .I(N__31767));
    CascadeMux I__7737 (
            .O(N__31767),
            .I(N__31764));
    CascadeBuf I__7736 (
            .O(N__31764),
            .I(N__31761));
    CascadeMux I__7735 (
            .O(N__31761),
            .I(N__31758));
    CascadeBuf I__7734 (
            .O(N__31758),
            .I(N__31755));
    CascadeMux I__7733 (
            .O(N__31755),
            .I(N__31752));
    CascadeBuf I__7732 (
            .O(N__31752),
            .I(N__31749));
    CascadeMux I__7731 (
            .O(N__31749),
            .I(N__31746));
    CascadeBuf I__7730 (
            .O(N__31746),
            .I(N__31743));
    CascadeMux I__7729 (
            .O(N__31743),
            .I(N__31740));
    CascadeBuf I__7728 (
            .O(N__31740),
            .I(N__31737));
    CascadeMux I__7727 (
            .O(N__31737),
            .I(N__31734));
    CascadeBuf I__7726 (
            .O(N__31734),
            .I(N__31731));
    CascadeMux I__7725 (
            .O(N__31731),
            .I(N__31728));
    CascadeBuf I__7724 (
            .O(N__31728),
            .I(N__31725));
    CascadeMux I__7723 (
            .O(N__31725),
            .I(N__31722));
    CascadeBuf I__7722 (
            .O(N__31722),
            .I(N__31719));
    CascadeMux I__7721 (
            .O(N__31719),
            .I(N__31716));
    CascadeBuf I__7720 (
            .O(N__31716),
            .I(N__31713));
    CascadeMux I__7719 (
            .O(N__31713),
            .I(N__31710));
    CascadeBuf I__7718 (
            .O(N__31710),
            .I(N__31707));
    CascadeMux I__7717 (
            .O(N__31707),
            .I(N__31704));
    CascadeBuf I__7716 (
            .O(N__31704),
            .I(N__31701));
    CascadeMux I__7715 (
            .O(N__31701),
            .I(N__31698));
    InMux I__7714 (
            .O(N__31698),
            .I(N__31695));
    LocalMux I__7713 (
            .O(N__31695),
            .I(N__31692));
    Odrv4 I__7712 (
            .O(N__31692),
            .I(M_this_ppu_sprites_addr_4));
    InMux I__7711 (
            .O(N__31689),
            .I(N__31686));
    LocalMux I__7710 (
            .O(N__31686),
            .I(N__31683));
    Span4Mux_v I__7709 (
            .O(N__31683),
            .I(N__31680));
    Span4Mux_v I__7708 (
            .O(N__31680),
            .I(N__31677));
    Span4Mux_v I__7707 (
            .O(N__31677),
            .I(N__31674));
    Span4Mux_v I__7706 (
            .O(N__31674),
            .I(N__31671));
    Odrv4 I__7705 (
            .O(N__31671),
            .I(port_address_in_7));
    InMux I__7704 (
            .O(N__31668),
            .I(N__31665));
    LocalMux I__7703 (
            .O(N__31665),
            .I(N__31662));
    IoSpan4Mux I__7702 (
            .O(N__31662),
            .I(N__31659));
    Odrv4 I__7701 (
            .O(N__31659),
            .I(port_address_in_4));
    CascadeMux I__7700 (
            .O(N__31656),
            .I(N__31653));
    InMux I__7699 (
            .O(N__31653),
            .I(N__31650));
    LocalMux I__7698 (
            .O(N__31650),
            .I(N__31646));
    InMux I__7697 (
            .O(N__31649),
            .I(N__31643));
    Span4Mux_s2_h I__7696 (
            .O(N__31646),
            .I(N__31640));
    LocalMux I__7695 (
            .O(N__31643),
            .I(N__31637));
    Sp12to4 I__7694 (
            .O(N__31640),
            .I(N__31634));
    Span4Mux_h I__7693 (
            .O(N__31637),
            .I(N__31631));
    Span12Mux_s11_v I__7692 (
            .O(N__31634),
            .I(N__31628));
    Span4Mux_v I__7691 (
            .O(N__31631),
            .I(N__31625));
    Span12Mux_h I__7690 (
            .O(N__31628),
            .I(N__31622));
    Sp12to4 I__7689 (
            .O(N__31625),
            .I(N__31619));
    Span12Mux_h I__7688 (
            .O(N__31622),
            .I(N__31616));
    Span12Mux_h I__7687 (
            .O(N__31619),
            .I(N__31613));
    Odrv12 I__7686 (
            .O(N__31616),
            .I(port_rw_in));
    Odrv12 I__7685 (
            .O(N__31613),
            .I(port_rw_in));
    InMux I__7684 (
            .O(N__31608),
            .I(N__31605));
    LocalMux I__7683 (
            .O(N__31605),
            .I(N__31602));
    Span12Mux_v I__7682 (
            .O(N__31602),
            .I(N__31599));
    Odrv12 I__7681 (
            .O(N__31599),
            .I(port_address_in_3));
    InMux I__7680 (
            .O(N__31596),
            .I(N__31593));
    LocalMux I__7679 (
            .O(N__31593),
            .I(N__31590));
    Span12Mux_h I__7678 (
            .O(N__31590),
            .I(N__31587));
    Odrv12 I__7677 (
            .O(N__31587),
            .I(\this_start_data_delay.un1_M_this_state_q_17_i_o2_1Z0Z_4 ));
    IoInMux I__7676 (
            .O(N__31584),
            .I(N__31581));
    LocalMux I__7675 (
            .O(N__31581),
            .I(N__31578));
    Span4Mux_s1_v I__7674 (
            .O(N__31578),
            .I(N__31574));
    InMux I__7673 (
            .O(N__31577),
            .I(N__31571));
    Span4Mux_v I__7672 (
            .O(N__31574),
            .I(N__31568));
    LocalMux I__7671 (
            .O(N__31571),
            .I(N__31565));
    Odrv4 I__7670 (
            .O(N__31568),
            .I(M_this_external_address_qZ0Z_9));
    Odrv4 I__7669 (
            .O(N__31565),
            .I(M_this_external_address_qZ0Z_9));
    InMux I__7668 (
            .O(N__31560),
            .I(N__31557));
    LocalMux I__7667 (
            .O(N__31557),
            .I(N__31554));
    Odrv12 I__7666 (
            .O(N__31554),
            .I(M_this_external_address_q_s_9));
    InMux I__7665 (
            .O(N__31551),
            .I(M_this_external_address_q_cry_8));
    InMux I__7664 (
            .O(N__31548),
            .I(M_this_external_address_q_cry_9));
    InMux I__7663 (
            .O(N__31545),
            .I(M_this_external_address_q_cry_10));
    IoInMux I__7662 (
            .O(N__31542),
            .I(N__31539));
    LocalMux I__7661 (
            .O(N__31539),
            .I(N__31534));
    CascadeMux I__7660 (
            .O(N__31538),
            .I(N__31531));
    InMux I__7659 (
            .O(N__31537),
            .I(N__31528));
    Sp12to4 I__7658 (
            .O(N__31534),
            .I(N__31525));
    InMux I__7657 (
            .O(N__31531),
            .I(N__31522));
    LocalMux I__7656 (
            .O(N__31528),
            .I(N__31519));
    Odrv12 I__7655 (
            .O(N__31525),
            .I(M_this_external_address_qZ0Z_12));
    LocalMux I__7654 (
            .O(N__31522),
            .I(M_this_external_address_qZ0Z_12));
    Odrv4 I__7653 (
            .O(N__31519),
            .I(M_this_external_address_qZ0Z_12));
    InMux I__7652 (
            .O(N__31512),
            .I(N__31509));
    LocalMux I__7651 (
            .O(N__31509),
            .I(N__31506));
    Odrv4 I__7650 (
            .O(N__31506),
            .I(M_this_external_address_q_cry_11_THRU_CO));
    InMux I__7649 (
            .O(N__31503),
            .I(M_this_external_address_q_cry_11));
    IoInMux I__7648 (
            .O(N__31500),
            .I(N__31497));
    LocalMux I__7647 (
            .O(N__31497),
            .I(N__31494));
    IoSpan4Mux I__7646 (
            .O(N__31494),
            .I(N__31491));
    Span4Mux_s2_h I__7645 (
            .O(N__31491),
            .I(N__31487));
    InMux I__7644 (
            .O(N__31490),
            .I(N__31483));
    Span4Mux_h I__7643 (
            .O(N__31487),
            .I(N__31480));
    InMux I__7642 (
            .O(N__31486),
            .I(N__31477));
    LocalMux I__7641 (
            .O(N__31483),
            .I(N__31474));
    Odrv4 I__7640 (
            .O(N__31480),
            .I(M_this_external_address_qZ0Z_13));
    LocalMux I__7639 (
            .O(N__31477),
            .I(M_this_external_address_qZ0Z_13));
    Odrv12 I__7638 (
            .O(N__31474),
            .I(M_this_external_address_qZ0Z_13));
    CascadeMux I__7637 (
            .O(N__31467),
            .I(N__31464));
    InMux I__7636 (
            .O(N__31464),
            .I(N__31461));
    LocalMux I__7635 (
            .O(N__31461),
            .I(N__31458));
    Odrv12 I__7634 (
            .O(N__31458),
            .I(M_this_external_address_q_cry_12_THRU_CO));
    InMux I__7633 (
            .O(N__31455),
            .I(M_this_external_address_q_cry_12));
    IoInMux I__7632 (
            .O(N__31452),
            .I(N__31449));
    LocalMux I__7631 (
            .O(N__31449),
            .I(N__31446));
    Span4Mux_s3_h I__7630 (
            .O(N__31446),
            .I(N__31443));
    Span4Mux_v I__7629 (
            .O(N__31443),
            .I(N__31438));
    CascadeMux I__7628 (
            .O(N__31442),
            .I(N__31435));
    InMux I__7627 (
            .O(N__31441),
            .I(N__31432));
    Span4Mux_h I__7626 (
            .O(N__31438),
            .I(N__31429));
    InMux I__7625 (
            .O(N__31435),
            .I(N__31426));
    LocalMux I__7624 (
            .O(N__31432),
            .I(N__31423));
    Odrv4 I__7623 (
            .O(N__31429),
            .I(M_this_external_address_qZ0Z_14));
    LocalMux I__7622 (
            .O(N__31426),
            .I(M_this_external_address_qZ0Z_14));
    Odrv4 I__7621 (
            .O(N__31423),
            .I(M_this_external_address_qZ0Z_14));
    InMux I__7620 (
            .O(N__31416),
            .I(N__31413));
    LocalMux I__7619 (
            .O(N__31413),
            .I(N__31410));
    Odrv4 I__7618 (
            .O(N__31410),
            .I(M_this_external_address_q_cry_13_THRU_CO));
    InMux I__7617 (
            .O(N__31407),
            .I(M_this_external_address_q_cry_13));
    IoInMux I__7616 (
            .O(N__31404),
            .I(N__31401));
    LocalMux I__7615 (
            .O(N__31401),
            .I(N__31398));
    Span12Mux_s9_h I__7614 (
            .O(N__31398),
            .I(N__31394));
    InMux I__7613 (
            .O(N__31397),
            .I(N__31391));
    Span12Mux_v I__7612 (
            .O(N__31394),
            .I(N__31388));
    LocalMux I__7611 (
            .O(N__31391),
            .I(N__31385));
    Odrv12 I__7610 (
            .O(N__31388),
            .I(M_this_external_address_qZ0Z_15));
    Odrv12 I__7609 (
            .O(N__31385),
            .I(M_this_external_address_qZ0Z_15));
    InMux I__7608 (
            .O(N__31380),
            .I(M_this_external_address_q_cry_14));
    CascadeMux I__7607 (
            .O(N__31377),
            .I(N__31374));
    InMux I__7606 (
            .O(N__31374),
            .I(N__31371));
    LocalMux I__7605 (
            .O(N__31371),
            .I(N__31368));
    Odrv4 I__7604 (
            .O(N__31368),
            .I(M_this_external_address_q_s_15));
    InMux I__7603 (
            .O(N__31365),
            .I(N__31362));
    LocalMux I__7602 (
            .O(N__31362),
            .I(M_this_external_address_q_s_11));
    InMux I__7601 (
            .O(N__31359),
            .I(N__31352));
    InMux I__7600 (
            .O(N__31358),
            .I(N__31349));
    InMux I__7599 (
            .O(N__31357),
            .I(N__31346));
    InMux I__7598 (
            .O(N__31356),
            .I(N__31343));
    CascadeMux I__7597 (
            .O(N__31355),
            .I(N__31339));
    LocalMux I__7596 (
            .O(N__31352),
            .I(N__31334));
    LocalMux I__7595 (
            .O(N__31349),
            .I(N__31334));
    LocalMux I__7594 (
            .O(N__31346),
            .I(N__31331));
    LocalMux I__7593 (
            .O(N__31343),
            .I(N__31327));
    CascadeMux I__7592 (
            .O(N__31342),
            .I(N__31324));
    InMux I__7591 (
            .O(N__31339),
            .I(N__31319));
    Span4Mux_v I__7590 (
            .O(N__31334),
            .I(N__31314));
    Span4Mux_h I__7589 (
            .O(N__31331),
            .I(N__31314));
    InMux I__7588 (
            .O(N__31330),
            .I(N__31311));
    Span4Mux_v I__7587 (
            .O(N__31327),
            .I(N__31308));
    InMux I__7586 (
            .O(N__31324),
            .I(N__31305));
    InMux I__7585 (
            .O(N__31323),
            .I(N__31300));
    InMux I__7584 (
            .O(N__31322),
            .I(N__31300));
    LocalMux I__7583 (
            .O(N__31319),
            .I(N__31297));
    Span4Mux_v I__7582 (
            .O(N__31314),
            .I(N__31290));
    LocalMux I__7581 (
            .O(N__31311),
            .I(N__31290));
    Span4Mux_h I__7580 (
            .O(N__31308),
            .I(N__31287));
    LocalMux I__7579 (
            .O(N__31305),
            .I(N__31284));
    LocalMux I__7578 (
            .O(N__31300),
            .I(N__31281));
    Span4Mux_h I__7577 (
            .O(N__31297),
            .I(N__31278));
    InMux I__7576 (
            .O(N__31296),
            .I(N__31275));
    CascadeMux I__7575 (
            .O(N__31295),
            .I(N__31272));
    Span4Mux_v I__7574 (
            .O(N__31290),
            .I(N__31269));
    Span4Mux_h I__7573 (
            .O(N__31287),
            .I(N__31264));
    Span4Mux_v I__7572 (
            .O(N__31284),
            .I(N__31264));
    Span4Mux_v I__7571 (
            .O(N__31281),
            .I(N__31257));
    Span4Mux_h I__7570 (
            .O(N__31278),
            .I(N__31257));
    LocalMux I__7569 (
            .O(N__31275),
            .I(N__31257));
    InMux I__7568 (
            .O(N__31272),
            .I(N__31254));
    Span4Mux_h I__7567 (
            .O(N__31269),
            .I(N__31251));
    Sp12to4 I__7566 (
            .O(N__31264),
            .I(N__31248));
    Span4Mux_v I__7565 (
            .O(N__31257),
            .I(N__31245));
    LocalMux I__7564 (
            .O(N__31254),
            .I(N__31242));
    Sp12to4 I__7563 (
            .O(N__31251),
            .I(N__31239));
    Span12Mux_h I__7562 (
            .O(N__31248),
            .I(N__31236));
    Sp12to4 I__7561 (
            .O(N__31245),
            .I(N__31233));
    Span4Mux_h I__7560 (
            .O(N__31242),
            .I(N__31230));
    Span12Mux_h I__7559 (
            .O(N__31239),
            .I(N__31225));
    Span12Mux_v I__7558 (
            .O(N__31236),
            .I(N__31225));
    Span12Mux_h I__7557 (
            .O(N__31233),
            .I(N__31222));
    Span4Mux_v I__7556 (
            .O(N__31230),
            .I(N__31219));
    Odrv12 I__7555 (
            .O(N__31225),
            .I(port_data_c_3));
    Odrv12 I__7554 (
            .O(N__31222),
            .I(port_data_c_3));
    Odrv4 I__7553 (
            .O(N__31219),
            .I(port_data_c_3));
    IoInMux I__7552 (
            .O(N__31212),
            .I(N__31209));
    LocalMux I__7551 (
            .O(N__31209),
            .I(N__31206));
    Span4Mux_s3_v I__7550 (
            .O(N__31206),
            .I(N__31203));
    Span4Mux_v I__7549 (
            .O(N__31203),
            .I(N__31199));
    InMux I__7548 (
            .O(N__31202),
            .I(N__31196));
    Odrv4 I__7547 (
            .O(N__31199),
            .I(M_this_external_address_qZ0Z_11));
    LocalMux I__7546 (
            .O(N__31196),
            .I(M_this_external_address_qZ0Z_11));
    IoInMux I__7545 (
            .O(N__31191),
            .I(N__31188));
    LocalMux I__7544 (
            .O(N__31188),
            .I(N__31185));
    Span4Mux_s1_v I__7543 (
            .O(N__31185),
            .I(N__31182));
    Sp12to4 I__7542 (
            .O(N__31182),
            .I(N__31179));
    Span12Mux_h I__7541 (
            .O(N__31179),
            .I(N__31175));
    InMux I__7540 (
            .O(N__31178),
            .I(N__31172));
    Odrv12 I__7539 (
            .O(N__31175),
            .I(M_this_external_address_qZ0Z_0));
    LocalMux I__7538 (
            .O(N__31172),
            .I(M_this_external_address_qZ0Z_0));
    InMux I__7537 (
            .O(N__31167),
            .I(bfn_26_23_0_));
    IoInMux I__7536 (
            .O(N__31164),
            .I(N__31161));
    LocalMux I__7535 (
            .O(N__31161),
            .I(N__31158));
    Sp12to4 I__7534 (
            .O(N__31158),
            .I(N__31154));
    InMux I__7533 (
            .O(N__31157),
            .I(N__31151));
    Odrv12 I__7532 (
            .O(N__31154),
            .I(M_this_external_address_qZ0Z_1));
    LocalMux I__7531 (
            .O(N__31151),
            .I(M_this_external_address_qZ0Z_1));
    InMux I__7530 (
            .O(N__31146),
            .I(M_this_external_address_q_cry_0));
    IoInMux I__7529 (
            .O(N__31143),
            .I(N__31140));
    LocalMux I__7528 (
            .O(N__31140),
            .I(N__31137));
    IoSpan4Mux I__7527 (
            .O(N__31137),
            .I(N__31134));
    Span4Mux_s2_v I__7526 (
            .O(N__31134),
            .I(N__31131));
    Span4Mux_v I__7525 (
            .O(N__31131),
            .I(N__31127));
    InMux I__7524 (
            .O(N__31130),
            .I(N__31124));
    Odrv4 I__7523 (
            .O(N__31127),
            .I(M_this_external_address_qZ0Z_2));
    LocalMux I__7522 (
            .O(N__31124),
            .I(M_this_external_address_qZ0Z_2));
    InMux I__7521 (
            .O(N__31119),
            .I(M_this_external_address_q_cry_1));
    IoInMux I__7520 (
            .O(N__31116),
            .I(N__31113));
    LocalMux I__7519 (
            .O(N__31113),
            .I(N__31110));
    Span4Mux_s2_h I__7518 (
            .O(N__31110),
            .I(N__31107));
    Span4Mux_h I__7517 (
            .O(N__31107),
            .I(N__31104));
    Span4Mux_v I__7516 (
            .O(N__31104),
            .I(N__31100));
    InMux I__7515 (
            .O(N__31103),
            .I(N__31097));
    Odrv4 I__7514 (
            .O(N__31100),
            .I(M_this_external_address_qZ0Z_3));
    LocalMux I__7513 (
            .O(N__31097),
            .I(M_this_external_address_qZ0Z_3));
    InMux I__7512 (
            .O(N__31092),
            .I(M_this_external_address_q_cry_2));
    IoInMux I__7511 (
            .O(N__31089),
            .I(N__31086));
    LocalMux I__7510 (
            .O(N__31086),
            .I(N__31082));
    InMux I__7509 (
            .O(N__31085),
            .I(N__31079));
    Odrv12 I__7508 (
            .O(N__31082),
            .I(M_this_external_address_qZ0Z_4));
    LocalMux I__7507 (
            .O(N__31079),
            .I(M_this_external_address_qZ0Z_4));
    InMux I__7506 (
            .O(N__31074),
            .I(M_this_external_address_q_cry_3));
    IoInMux I__7505 (
            .O(N__31071),
            .I(N__31068));
    LocalMux I__7504 (
            .O(N__31068),
            .I(N__31065));
    IoSpan4Mux I__7503 (
            .O(N__31065),
            .I(N__31062));
    Sp12to4 I__7502 (
            .O(N__31062),
            .I(N__31058));
    InMux I__7501 (
            .O(N__31061),
            .I(N__31055));
    Odrv12 I__7500 (
            .O(N__31058),
            .I(M_this_external_address_qZ0Z_5));
    LocalMux I__7499 (
            .O(N__31055),
            .I(M_this_external_address_qZ0Z_5));
    InMux I__7498 (
            .O(N__31050),
            .I(M_this_external_address_q_cry_4));
    IoInMux I__7497 (
            .O(N__31047),
            .I(N__31044));
    LocalMux I__7496 (
            .O(N__31044),
            .I(N__31041));
    Span12Mux_s6_h I__7495 (
            .O(N__31041),
            .I(N__31037));
    InMux I__7494 (
            .O(N__31040),
            .I(N__31034));
    Odrv12 I__7493 (
            .O(N__31037),
            .I(M_this_external_address_qZ0Z_6));
    LocalMux I__7492 (
            .O(N__31034),
            .I(M_this_external_address_qZ0Z_6));
    InMux I__7491 (
            .O(N__31029),
            .I(M_this_external_address_q_cry_5));
    IoInMux I__7490 (
            .O(N__31026),
            .I(N__31023));
    LocalMux I__7489 (
            .O(N__31023),
            .I(N__31020));
    Span4Mux_s2_h I__7488 (
            .O(N__31020),
            .I(N__31017));
    Span4Mux_h I__7487 (
            .O(N__31017),
            .I(N__31014));
    Sp12to4 I__7486 (
            .O(N__31014),
            .I(N__31011));
    Span12Mux_v I__7485 (
            .O(N__31011),
            .I(N__31007));
    InMux I__7484 (
            .O(N__31010),
            .I(N__31004));
    Odrv12 I__7483 (
            .O(N__31007),
            .I(M_this_external_address_qZ0Z_7));
    LocalMux I__7482 (
            .O(N__31004),
            .I(M_this_external_address_qZ0Z_7));
    InMux I__7481 (
            .O(N__30999),
            .I(M_this_external_address_q_cry_6));
    IoInMux I__7480 (
            .O(N__30996),
            .I(N__30993));
    LocalMux I__7479 (
            .O(N__30993),
            .I(N__30990));
    Span4Mux_s0_v I__7478 (
            .O(N__30990),
            .I(N__30987));
    Sp12to4 I__7477 (
            .O(N__30987),
            .I(N__30983));
    InMux I__7476 (
            .O(N__30986),
            .I(N__30980));
    Span12Mux_h I__7475 (
            .O(N__30983),
            .I(N__30977));
    LocalMux I__7474 (
            .O(N__30980),
            .I(N__30974));
    Odrv12 I__7473 (
            .O(N__30977),
            .I(M_this_external_address_qZ0Z_8));
    Odrv12 I__7472 (
            .O(N__30974),
            .I(M_this_external_address_qZ0Z_8));
    InMux I__7471 (
            .O(N__30969),
            .I(N__30966));
    LocalMux I__7470 (
            .O(N__30966),
            .I(N__30963));
    Span4Mux_h I__7469 (
            .O(N__30963),
            .I(N__30960));
    Odrv4 I__7468 (
            .O(N__30960),
            .I(M_this_external_address_q_s_8));
    InMux I__7467 (
            .O(N__30957),
            .I(bfn_26_24_0_));
    InMux I__7466 (
            .O(N__30954),
            .I(N__30951));
    LocalMux I__7465 (
            .O(N__30951),
            .I(N__30948));
    Odrv4 I__7464 (
            .O(N__30948),
            .I(M_this_external_address_q_3_0_12));
    InMux I__7463 (
            .O(N__30945),
            .I(N__30942));
    LocalMux I__7462 (
            .O(N__30942),
            .I(N__30939));
    Odrv4 I__7461 (
            .O(N__30939),
            .I(M_this_external_address_q_3_14));
    CascadeMux I__7460 (
            .O(N__30936),
            .I(N__30931));
    InMux I__7459 (
            .O(N__30935),
            .I(N__30925));
    CascadeMux I__7458 (
            .O(N__30934),
            .I(N__30922));
    InMux I__7457 (
            .O(N__30931),
            .I(N__30919));
    InMux I__7456 (
            .O(N__30930),
            .I(N__30916));
    InMux I__7455 (
            .O(N__30929),
            .I(N__30910));
    InMux I__7454 (
            .O(N__30928),
            .I(N__30907));
    LocalMux I__7453 (
            .O(N__30925),
            .I(N__30904));
    InMux I__7452 (
            .O(N__30922),
            .I(N__30901));
    LocalMux I__7451 (
            .O(N__30919),
            .I(N__30896));
    LocalMux I__7450 (
            .O(N__30916),
            .I(N__30896));
    CascadeMux I__7449 (
            .O(N__30915),
            .I(N__30893));
    CascadeMux I__7448 (
            .O(N__30914),
            .I(N__30890));
    InMux I__7447 (
            .O(N__30913),
            .I(N__30887));
    LocalMux I__7446 (
            .O(N__30910),
            .I(N__30884));
    LocalMux I__7445 (
            .O(N__30907),
            .I(N__30881));
    Span4Mux_h I__7444 (
            .O(N__30904),
            .I(N__30876));
    LocalMux I__7443 (
            .O(N__30901),
            .I(N__30876));
    Span4Mux_v I__7442 (
            .O(N__30896),
            .I(N__30873));
    InMux I__7441 (
            .O(N__30893),
            .I(N__30870));
    InMux I__7440 (
            .O(N__30890),
            .I(N__30867));
    LocalMux I__7439 (
            .O(N__30887),
            .I(N__30864));
    Span4Mux_v I__7438 (
            .O(N__30884),
            .I(N__30858));
    Span4Mux_h I__7437 (
            .O(N__30881),
            .I(N__30858));
    Span4Mux_v I__7436 (
            .O(N__30876),
            .I(N__30855));
    Span4Mux_v I__7435 (
            .O(N__30873),
            .I(N__30850));
    LocalMux I__7434 (
            .O(N__30870),
            .I(N__30850));
    LocalMux I__7433 (
            .O(N__30867),
            .I(N__30847));
    Span4Mux_h I__7432 (
            .O(N__30864),
            .I(N__30843));
    InMux I__7431 (
            .O(N__30863),
            .I(N__30840));
    Span4Mux_v I__7430 (
            .O(N__30858),
            .I(N__30837));
    Span4Mux_v I__7429 (
            .O(N__30855),
            .I(N__30832));
    Span4Mux_v I__7428 (
            .O(N__30850),
            .I(N__30832));
    Span4Mux_v I__7427 (
            .O(N__30847),
            .I(N__30829));
    InMux I__7426 (
            .O(N__30846),
            .I(N__30826));
    Span4Mux_v I__7425 (
            .O(N__30843),
            .I(N__30823));
    LocalMux I__7424 (
            .O(N__30840),
            .I(N__30820));
    Span4Mux_v I__7423 (
            .O(N__30837),
            .I(N__30817));
    Sp12to4 I__7422 (
            .O(N__30832),
            .I(N__30812));
    Sp12to4 I__7421 (
            .O(N__30829),
            .I(N__30812));
    LocalMux I__7420 (
            .O(N__30826),
            .I(N__30809));
    Span4Mux_v I__7419 (
            .O(N__30823),
            .I(N__30804));
    Span4Mux_h I__7418 (
            .O(N__30820),
            .I(N__30804));
    Span4Mux_v I__7417 (
            .O(N__30817),
            .I(N__30801));
    Span12Mux_h I__7416 (
            .O(N__30812),
            .I(N__30796));
    Span12Mux_v I__7415 (
            .O(N__30809),
            .I(N__30796));
    Span4Mux_v I__7414 (
            .O(N__30804),
            .I(N__30793));
    Odrv4 I__7413 (
            .O(N__30801),
            .I(port_data_c_1));
    Odrv12 I__7412 (
            .O(N__30796),
            .I(port_data_c_1));
    Odrv4 I__7411 (
            .O(N__30793),
            .I(port_data_c_1));
    CEMux I__7410 (
            .O(N__30786),
            .I(N__30782));
    CEMux I__7409 (
            .O(N__30785),
            .I(N__30779));
    LocalMux I__7408 (
            .O(N__30782),
            .I(N__30776));
    LocalMux I__7407 (
            .O(N__30779),
            .I(N__30773));
    Span4Mux_v I__7406 (
            .O(N__30776),
            .I(N__30770));
    Span4Mux_h I__7405 (
            .O(N__30773),
            .I(N__30767));
    Odrv4 I__7404 (
            .O(N__30770),
            .I(\this_sprites_ram.mem_WE_2 ));
    Odrv4 I__7403 (
            .O(N__30767),
            .I(\this_sprites_ram.mem_WE_2 ));
    InMux I__7402 (
            .O(N__30762),
            .I(N__30756));
    InMux I__7401 (
            .O(N__30761),
            .I(N__30756));
    LocalMux I__7400 (
            .O(N__30756),
            .I(N__30748));
    InMux I__7399 (
            .O(N__30755),
            .I(N__30745));
    InMux I__7398 (
            .O(N__30754),
            .I(N__30740));
    InMux I__7397 (
            .O(N__30753),
            .I(N__30740));
    InMux I__7396 (
            .O(N__30752),
            .I(N__30734));
    InMux I__7395 (
            .O(N__30751),
            .I(N__30734));
    Span4Mux_v I__7394 (
            .O(N__30748),
            .I(N__30729));
    LocalMux I__7393 (
            .O(N__30745),
            .I(N__30729));
    LocalMux I__7392 (
            .O(N__30740),
            .I(N__30726));
    InMux I__7391 (
            .O(N__30739),
            .I(N__30723));
    LocalMux I__7390 (
            .O(N__30734),
            .I(N__30720));
    Span4Mux_v I__7389 (
            .O(N__30729),
            .I(N__30713));
    Span4Mux_v I__7388 (
            .O(N__30726),
            .I(N__30713));
    LocalMux I__7387 (
            .O(N__30723),
            .I(N__30713));
    Span4Mux_h I__7386 (
            .O(N__30720),
            .I(N__30708));
    Span4Mux_h I__7385 (
            .O(N__30713),
            .I(N__30708));
    Odrv4 I__7384 (
            .O(N__30708),
            .I(M_this_sprites_ram_write_en_0));
    CascadeMux I__7383 (
            .O(N__30705),
            .I(N__30701));
    CascadeMux I__7382 (
            .O(N__30704),
            .I(N__30694));
    InMux I__7381 (
            .O(N__30701),
            .I(N__30689));
    InMux I__7380 (
            .O(N__30700),
            .I(N__30689));
    CascadeMux I__7379 (
            .O(N__30699),
            .I(N__30686));
    CascadeMux I__7378 (
            .O(N__30698),
            .I(N__30682));
    CascadeMux I__7377 (
            .O(N__30697),
            .I(N__30678));
    InMux I__7376 (
            .O(N__30694),
            .I(N__30674));
    LocalMux I__7375 (
            .O(N__30689),
            .I(N__30671));
    InMux I__7374 (
            .O(N__30686),
            .I(N__30668));
    InMux I__7373 (
            .O(N__30685),
            .I(N__30663));
    InMux I__7372 (
            .O(N__30682),
            .I(N__30663));
    InMux I__7371 (
            .O(N__30681),
            .I(N__30658));
    InMux I__7370 (
            .O(N__30678),
            .I(N__30658));
    CascadeMux I__7369 (
            .O(N__30677),
            .I(N__30654));
    LocalMux I__7368 (
            .O(N__30674),
            .I(N__30648));
    Span4Mux_v I__7367 (
            .O(N__30671),
            .I(N__30648));
    LocalMux I__7366 (
            .O(N__30668),
            .I(N__30643));
    LocalMux I__7365 (
            .O(N__30663),
            .I(N__30643));
    LocalMux I__7364 (
            .O(N__30658),
            .I(N__30640));
    InMux I__7363 (
            .O(N__30657),
            .I(N__30635));
    InMux I__7362 (
            .O(N__30654),
            .I(N__30635));
    InMux I__7361 (
            .O(N__30653),
            .I(N__30632));
    Span4Mux_v I__7360 (
            .O(N__30648),
            .I(N__30627));
    Span4Mux_v I__7359 (
            .O(N__30643),
            .I(N__30627));
    Span4Mux_h I__7358 (
            .O(N__30640),
            .I(N__30624));
    LocalMux I__7357 (
            .O(N__30635),
            .I(M_this_sprites_address_qZ0Z_12));
    LocalMux I__7356 (
            .O(N__30632),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv4 I__7355 (
            .O(N__30627),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv4 I__7354 (
            .O(N__30624),
            .I(M_this_sprites_address_qZ0Z_12));
    CascadeMux I__7353 (
            .O(N__30615),
            .I(N__30611));
    CascadeMux I__7352 (
            .O(N__30614),
            .I(N__30607));
    InMux I__7351 (
            .O(N__30611),
            .I(N__30600));
    InMux I__7350 (
            .O(N__30610),
            .I(N__30600));
    InMux I__7349 (
            .O(N__30607),
            .I(N__30595));
    InMux I__7348 (
            .O(N__30606),
            .I(N__30595));
    InMux I__7347 (
            .O(N__30605),
            .I(N__30588));
    LocalMux I__7346 (
            .O(N__30600),
            .I(N__30585));
    LocalMux I__7345 (
            .O(N__30595),
            .I(N__30582));
    InMux I__7344 (
            .O(N__30594),
            .I(N__30577));
    InMux I__7343 (
            .O(N__30593),
            .I(N__30577));
    CascadeMux I__7342 (
            .O(N__30592),
            .I(N__30574));
    InMux I__7341 (
            .O(N__30591),
            .I(N__30569));
    LocalMux I__7340 (
            .O(N__30588),
            .I(N__30564));
    Span4Mux_v I__7339 (
            .O(N__30585),
            .I(N__30564));
    Span4Mux_h I__7338 (
            .O(N__30582),
            .I(N__30561));
    LocalMux I__7337 (
            .O(N__30577),
            .I(N__30558));
    InMux I__7336 (
            .O(N__30574),
            .I(N__30555));
    InMux I__7335 (
            .O(N__30573),
            .I(N__30552));
    InMux I__7334 (
            .O(N__30572),
            .I(N__30549));
    LocalMux I__7333 (
            .O(N__30569),
            .I(N__30542));
    Span4Mux_v I__7332 (
            .O(N__30564),
            .I(N__30542));
    Span4Mux_v I__7331 (
            .O(N__30561),
            .I(N__30542));
    Span4Mux_h I__7330 (
            .O(N__30558),
            .I(N__30539));
    LocalMux I__7329 (
            .O(N__30555),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__7328 (
            .O(N__30552),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__7327 (
            .O(N__30549),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv4 I__7326 (
            .O(N__30542),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv4 I__7325 (
            .O(N__30539),
            .I(M_this_sprites_address_qZ0Z_11));
    InMux I__7324 (
            .O(N__30528),
            .I(N__30521));
    InMux I__7323 (
            .O(N__30527),
            .I(N__30521));
    CascadeMux I__7322 (
            .O(N__30526),
            .I(N__30516));
    LocalMux I__7321 (
            .O(N__30521),
            .I(N__30510));
    InMux I__7320 (
            .O(N__30520),
            .I(N__30505));
    InMux I__7319 (
            .O(N__30519),
            .I(N__30505));
    InMux I__7318 (
            .O(N__30516),
            .I(N__30500));
    InMux I__7317 (
            .O(N__30515),
            .I(N__30500));
    InMux I__7316 (
            .O(N__30514),
            .I(N__30497));
    CascadeMux I__7315 (
            .O(N__30513),
            .I(N__30494));
    Span4Mux_v I__7314 (
            .O(N__30510),
            .I(N__30491));
    LocalMux I__7313 (
            .O(N__30505),
            .I(N__30488));
    LocalMux I__7312 (
            .O(N__30500),
            .I(N__30485));
    LocalMux I__7311 (
            .O(N__30497),
            .I(N__30482));
    InMux I__7310 (
            .O(N__30494),
            .I(N__30477));
    Span4Mux_v I__7309 (
            .O(N__30491),
            .I(N__30472));
    Span4Mux_v I__7308 (
            .O(N__30488),
            .I(N__30472));
    Span4Mux_h I__7307 (
            .O(N__30485),
            .I(N__30469));
    Span4Mux_h I__7306 (
            .O(N__30482),
            .I(N__30466));
    InMux I__7305 (
            .O(N__30481),
            .I(N__30463));
    InMux I__7304 (
            .O(N__30480),
            .I(N__30460));
    LocalMux I__7303 (
            .O(N__30477),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__7302 (
            .O(N__30472),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__7301 (
            .O(N__30469),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__7300 (
            .O(N__30466),
            .I(M_this_sprites_address_qZ0Z_13));
    LocalMux I__7299 (
            .O(N__30463),
            .I(M_this_sprites_address_qZ0Z_13));
    LocalMux I__7298 (
            .O(N__30460),
            .I(M_this_sprites_address_qZ0Z_13));
    CEMux I__7297 (
            .O(N__30447),
            .I(N__30443));
    CEMux I__7296 (
            .O(N__30446),
            .I(N__30440));
    LocalMux I__7295 (
            .O(N__30443),
            .I(N__30435));
    LocalMux I__7294 (
            .O(N__30440),
            .I(N__30435));
    Span4Mux_v I__7293 (
            .O(N__30435),
            .I(N__30432));
    Odrv4 I__7292 (
            .O(N__30432),
            .I(\this_sprites_ram.mem_WE_0 ));
    CascadeMux I__7291 (
            .O(N__30429),
            .I(N__30426));
    InMux I__7290 (
            .O(N__30426),
            .I(N__30423));
    LocalMux I__7289 (
            .O(N__30423),
            .I(N__30420));
    Span4Mux_v I__7288 (
            .O(N__30420),
            .I(N__30417));
    Span4Mux_h I__7287 (
            .O(N__30417),
            .I(N__30414));
    Span4Mux_h I__7286 (
            .O(N__30414),
            .I(N__30411));
    Sp12to4 I__7285 (
            .O(N__30411),
            .I(N__30408));
    Odrv12 I__7284 (
            .O(N__30408),
            .I(M_this_map_ram_read_data_4));
    InMux I__7283 (
            .O(N__30405),
            .I(N__30402));
    LocalMux I__7282 (
            .O(N__30402),
            .I(N__30399));
    Span12Mux_s10_h I__7281 (
            .O(N__30399),
            .I(N__30396));
    Span12Mux_v I__7280 (
            .O(N__30396),
            .I(N__30393));
    Odrv12 I__7279 (
            .O(N__30393),
            .I(\this_ppu.un10_sprites_addr_cry_1_c_RNIOM6BZ0 ));
    CascadeMux I__7278 (
            .O(N__30390),
            .I(N__30387));
    CascadeBuf I__7277 (
            .O(N__30387),
            .I(N__30384));
    CascadeMux I__7276 (
            .O(N__30384),
            .I(N__30381));
    CascadeBuf I__7275 (
            .O(N__30381),
            .I(N__30378));
    CascadeMux I__7274 (
            .O(N__30378),
            .I(N__30375));
    CascadeBuf I__7273 (
            .O(N__30375),
            .I(N__30372));
    CascadeMux I__7272 (
            .O(N__30372),
            .I(N__30369));
    CascadeBuf I__7271 (
            .O(N__30369),
            .I(N__30366));
    CascadeMux I__7270 (
            .O(N__30366),
            .I(N__30363));
    CascadeBuf I__7269 (
            .O(N__30363),
            .I(N__30360));
    CascadeMux I__7268 (
            .O(N__30360),
            .I(N__30357));
    CascadeBuf I__7267 (
            .O(N__30357),
            .I(N__30354));
    CascadeMux I__7266 (
            .O(N__30354),
            .I(N__30351));
    CascadeBuf I__7265 (
            .O(N__30351),
            .I(N__30348));
    CascadeMux I__7264 (
            .O(N__30348),
            .I(N__30345));
    CascadeBuf I__7263 (
            .O(N__30345),
            .I(N__30342));
    CascadeMux I__7262 (
            .O(N__30342),
            .I(N__30339));
    CascadeBuf I__7261 (
            .O(N__30339),
            .I(N__30336));
    CascadeMux I__7260 (
            .O(N__30336),
            .I(N__30333));
    CascadeBuf I__7259 (
            .O(N__30333),
            .I(N__30330));
    CascadeMux I__7258 (
            .O(N__30330),
            .I(N__30327));
    CascadeBuf I__7257 (
            .O(N__30327),
            .I(N__30324));
    CascadeMux I__7256 (
            .O(N__30324),
            .I(N__30321));
    CascadeBuf I__7255 (
            .O(N__30321),
            .I(N__30318));
    CascadeMux I__7254 (
            .O(N__30318),
            .I(N__30315));
    CascadeBuf I__7253 (
            .O(N__30315),
            .I(N__30312));
    CascadeMux I__7252 (
            .O(N__30312),
            .I(N__30309));
    CascadeBuf I__7251 (
            .O(N__30309),
            .I(N__30306));
    CascadeMux I__7250 (
            .O(N__30306),
            .I(N__30303));
    CascadeBuf I__7249 (
            .O(N__30303),
            .I(N__30300));
    CascadeMux I__7248 (
            .O(N__30300),
            .I(N__30297));
    InMux I__7247 (
            .O(N__30297),
            .I(N__30294));
    LocalMux I__7246 (
            .O(N__30294),
            .I(M_this_ppu_sprites_addr_10));
    InMux I__7245 (
            .O(N__30291),
            .I(N__30288));
    LocalMux I__7244 (
            .O(N__30288),
            .I(N__30285));
    Span4Mux_s2_v I__7243 (
            .O(N__30285),
            .I(N__30282));
    Sp12to4 I__7242 (
            .O(N__30282),
            .I(N__30276));
    InMux I__7241 (
            .O(N__30281),
            .I(N__30273));
    CascadeMux I__7240 (
            .O(N__30280),
            .I(N__30270));
    InMux I__7239 (
            .O(N__30279),
            .I(N__30267));
    Span12Mux_h I__7238 (
            .O(N__30276),
            .I(N__30264));
    LocalMux I__7237 (
            .O(N__30273),
            .I(N__30261));
    InMux I__7236 (
            .O(N__30270),
            .I(N__30258));
    LocalMux I__7235 (
            .O(N__30267),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    Odrv12 I__7234 (
            .O(N__30264),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    Odrv4 I__7233 (
            .O(N__30261),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    LocalMux I__7232 (
            .O(N__30258),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    InMux I__7231 (
            .O(N__30249),
            .I(N__30246));
    LocalMux I__7230 (
            .O(N__30246),
            .I(N__30243));
    Span12Mux_v I__7229 (
            .O(N__30243),
            .I(N__30240));
    Span12Mux_h I__7228 (
            .O(N__30240),
            .I(N__30237));
    Odrv12 I__7227 (
            .O(N__30237),
            .I(\this_ppu.un3_sprites_addr_cry_4_c_RNI32FZ0Z8 ));
    CascadeMux I__7226 (
            .O(N__30234),
            .I(N__30231));
    CascadeBuf I__7225 (
            .O(N__30231),
            .I(N__30228));
    CascadeMux I__7224 (
            .O(N__30228),
            .I(N__30225));
    CascadeBuf I__7223 (
            .O(N__30225),
            .I(N__30222));
    CascadeMux I__7222 (
            .O(N__30222),
            .I(N__30219));
    CascadeBuf I__7221 (
            .O(N__30219),
            .I(N__30216));
    CascadeMux I__7220 (
            .O(N__30216),
            .I(N__30213));
    CascadeBuf I__7219 (
            .O(N__30213),
            .I(N__30210));
    CascadeMux I__7218 (
            .O(N__30210),
            .I(N__30207));
    CascadeBuf I__7217 (
            .O(N__30207),
            .I(N__30204));
    CascadeMux I__7216 (
            .O(N__30204),
            .I(N__30201));
    CascadeBuf I__7215 (
            .O(N__30201),
            .I(N__30198));
    CascadeMux I__7214 (
            .O(N__30198),
            .I(N__30195));
    CascadeBuf I__7213 (
            .O(N__30195),
            .I(N__30192));
    CascadeMux I__7212 (
            .O(N__30192),
            .I(N__30189));
    CascadeBuf I__7211 (
            .O(N__30189),
            .I(N__30186));
    CascadeMux I__7210 (
            .O(N__30186),
            .I(N__30183));
    CascadeBuf I__7209 (
            .O(N__30183),
            .I(N__30180));
    CascadeMux I__7208 (
            .O(N__30180),
            .I(N__30177));
    CascadeBuf I__7207 (
            .O(N__30177),
            .I(N__30174));
    CascadeMux I__7206 (
            .O(N__30174),
            .I(N__30171));
    CascadeBuf I__7205 (
            .O(N__30171),
            .I(N__30168));
    CascadeMux I__7204 (
            .O(N__30168),
            .I(N__30165));
    CascadeBuf I__7203 (
            .O(N__30165),
            .I(N__30162));
    CascadeMux I__7202 (
            .O(N__30162),
            .I(N__30159));
    CascadeBuf I__7201 (
            .O(N__30159),
            .I(N__30156));
    CascadeMux I__7200 (
            .O(N__30156),
            .I(N__30153));
    CascadeBuf I__7199 (
            .O(N__30153),
            .I(N__30150));
    CascadeMux I__7198 (
            .O(N__30150),
            .I(N__30147));
    CascadeBuf I__7197 (
            .O(N__30147),
            .I(N__30144));
    CascadeMux I__7196 (
            .O(N__30144),
            .I(N__30141));
    InMux I__7195 (
            .O(N__30141),
            .I(N__30138));
    LocalMux I__7194 (
            .O(N__30138),
            .I(M_this_ppu_sprites_addr_5));
    InMux I__7193 (
            .O(N__30135),
            .I(N__30132));
    LocalMux I__7192 (
            .O(N__30132),
            .I(N__30129));
    Span4Mux_v I__7191 (
            .O(N__30129),
            .I(N__30126));
    Span4Mux_v I__7190 (
            .O(N__30126),
            .I(N__30123));
    Span4Mux_v I__7189 (
            .O(N__30123),
            .I(N__30120));
    Odrv4 I__7188 (
            .O(N__30120),
            .I(\this_sprites_ram.mem_out_bus7_3 ));
    InMux I__7187 (
            .O(N__30117),
            .I(N__30114));
    LocalMux I__7186 (
            .O(N__30114),
            .I(N__30111));
    Odrv4 I__7185 (
            .O(N__30111),
            .I(\this_sprites_ram.mem_out_bus3_3 ));
    InMux I__7184 (
            .O(N__30108),
            .I(N__30102));
    InMux I__7183 (
            .O(N__30107),
            .I(N__30097));
    InMux I__7182 (
            .O(N__30106),
            .I(N__30092));
    InMux I__7181 (
            .O(N__30105),
            .I(N__30085));
    LocalMux I__7180 (
            .O(N__30102),
            .I(N__30082));
    InMux I__7179 (
            .O(N__30101),
            .I(N__30077));
    InMux I__7178 (
            .O(N__30100),
            .I(N__30077));
    LocalMux I__7177 (
            .O(N__30097),
            .I(N__30073));
    InMux I__7176 (
            .O(N__30096),
            .I(N__30068));
    InMux I__7175 (
            .O(N__30095),
            .I(N__30068));
    LocalMux I__7174 (
            .O(N__30092),
            .I(N__30065));
    InMux I__7173 (
            .O(N__30091),
            .I(N__30060));
    InMux I__7172 (
            .O(N__30090),
            .I(N__30060));
    InMux I__7171 (
            .O(N__30089),
            .I(N__30057));
    InMux I__7170 (
            .O(N__30088),
            .I(N__30053));
    LocalMux I__7169 (
            .O(N__30085),
            .I(N__30050));
    Span4Mux_v I__7168 (
            .O(N__30082),
            .I(N__30045));
    LocalMux I__7167 (
            .O(N__30077),
            .I(N__30045));
    InMux I__7166 (
            .O(N__30076),
            .I(N__30042));
    Span4Mux_v I__7165 (
            .O(N__30073),
            .I(N__30037));
    LocalMux I__7164 (
            .O(N__30068),
            .I(N__30037));
    Span4Mux_v I__7163 (
            .O(N__30065),
            .I(N__30032));
    LocalMux I__7162 (
            .O(N__30060),
            .I(N__30027));
    LocalMux I__7161 (
            .O(N__30057),
            .I(N__30027));
    InMux I__7160 (
            .O(N__30056),
            .I(N__30024));
    LocalMux I__7159 (
            .O(N__30053),
            .I(N__30015));
    Span4Mux_v I__7158 (
            .O(N__30050),
            .I(N__30015));
    Span4Mux_h I__7157 (
            .O(N__30045),
            .I(N__30015));
    LocalMux I__7156 (
            .O(N__30042),
            .I(N__30015));
    Span4Mux_h I__7155 (
            .O(N__30037),
            .I(N__30012));
    InMux I__7154 (
            .O(N__30036),
            .I(N__30007));
    InMux I__7153 (
            .O(N__30035),
            .I(N__30007));
    Span4Mux_v I__7152 (
            .O(N__30032),
            .I(N__30002));
    Span4Mux_h I__7151 (
            .O(N__30027),
            .I(N__30002));
    LocalMux I__7150 (
            .O(N__30024),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__7149 (
            .O(N__30015),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__7148 (
            .O(N__30012),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    LocalMux I__7147 (
            .O(N__30007),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__7146 (
            .O(N__30002),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    InMux I__7145 (
            .O(N__29991),
            .I(N__29988));
    LocalMux I__7144 (
            .O(N__29988),
            .I(N__29985));
    Span4Mux_h I__7143 (
            .O(N__29985),
            .I(N__29982));
    Odrv4 I__7142 (
            .O(N__29982),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ));
    InMux I__7141 (
            .O(N__29979),
            .I(N__29976));
    LocalMux I__7140 (
            .O(N__29976),
            .I(N__29973));
    Odrv12 I__7139 (
            .O(N__29973),
            .I(M_this_data_count_q_s_9));
    InMux I__7138 (
            .O(N__29970),
            .I(M_this_data_count_q_cry_8));
    CascadeMux I__7137 (
            .O(N__29967),
            .I(N__29964));
    InMux I__7136 (
            .O(N__29964),
            .I(N__29961));
    LocalMux I__7135 (
            .O(N__29961),
            .I(N__29956));
    InMux I__7134 (
            .O(N__29960),
            .I(N__29951));
    InMux I__7133 (
            .O(N__29959),
            .I(N__29951));
    Odrv4 I__7132 (
            .O(N__29956),
            .I(M_this_data_count_qZ0Z_10));
    LocalMux I__7131 (
            .O(N__29951),
            .I(M_this_data_count_qZ0Z_10));
    InMux I__7130 (
            .O(N__29946),
            .I(N__29943));
    LocalMux I__7129 (
            .O(N__29943),
            .I(M_this_data_count_q_cry_9_THRU_CO));
    InMux I__7128 (
            .O(N__29940),
            .I(M_this_data_count_q_cry_9));
    CascadeMux I__7127 (
            .O(N__29937),
            .I(N__29933));
    InMux I__7126 (
            .O(N__29936),
            .I(N__29930));
    InMux I__7125 (
            .O(N__29933),
            .I(N__29927));
    LocalMux I__7124 (
            .O(N__29930),
            .I(M_this_data_count_qZ0Z_11));
    LocalMux I__7123 (
            .O(N__29927),
            .I(M_this_data_count_qZ0Z_11));
    InMux I__7122 (
            .O(N__29922),
            .I(N__29919));
    LocalMux I__7121 (
            .O(N__29919),
            .I(M_this_data_count_q_s_11));
    InMux I__7120 (
            .O(N__29916),
            .I(M_this_data_count_q_cry_10));
    CascadeMux I__7119 (
            .O(N__29913),
            .I(N__29910));
    InMux I__7118 (
            .O(N__29910),
            .I(N__29906));
    InMux I__7117 (
            .O(N__29909),
            .I(N__29903));
    LocalMux I__7116 (
            .O(N__29906),
            .I(N__29900));
    LocalMux I__7115 (
            .O(N__29903),
            .I(N__29897));
    Odrv4 I__7114 (
            .O(N__29900),
            .I(M_this_data_count_qZ0Z_12));
    Odrv4 I__7113 (
            .O(N__29897),
            .I(M_this_data_count_qZ0Z_12));
    InMux I__7112 (
            .O(N__29892),
            .I(N__29889));
    LocalMux I__7111 (
            .O(N__29889),
            .I(N__29886));
    Odrv4 I__7110 (
            .O(N__29886),
            .I(M_this_data_count_q_s_12));
    InMux I__7109 (
            .O(N__29883),
            .I(M_this_data_count_q_cry_11));
    InMux I__7108 (
            .O(N__29880),
            .I(N__29876));
    InMux I__7107 (
            .O(N__29879),
            .I(N__29872));
    LocalMux I__7106 (
            .O(N__29876),
            .I(N__29869));
    InMux I__7105 (
            .O(N__29875),
            .I(N__29866));
    LocalMux I__7104 (
            .O(N__29872),
            .I(M_this_data_count_qZ0Z_13));
    Odrv4 I__7103 (
            .O(N__29869),
            .I(M_this_data_count_qZ0Z_13));
    LocalMux I__7102 (
            .O(N__29866),
            .I(M_this_data_count_qZ0Z_13));
    CascadeMux I__7101 (
            .O(N__29859),
            .I(N__29856));
    InMux I__7100 (
            .O(N__29856),
            .I(N__29853));
    LocalMux I__7099 (
            .O(N__29853),
            .I(N__29850));
    Odrv4 I__7098 (
            .O(N__29850),
            .I(M_this_data_count_q_cry_12_THRU_CO));
    InMux I__7097 (
            .O(N__29847),
            .I(M_this_data_count_q_cry_12));
    SRMux I__7096 (
            .O(N__29844),
            .I(N__29838));
    IoInMux I__7095 (
            .O(N__29843),
            .I(N__29832));
    SRMux I__7094 (
            .O(N__29842),
            .I(N__29829));
    SRMux I__7093 (
            .O(N__29841),
            .I(N__29826));
    LocalMux I__7092 (
            .O(N__29838),
            .I(N__29823));
    SRMux I__7091 (
            .O(N__29837),
            .I(N__29820));
    SRMux I__7090 (
            .O(N__29836),
            .I(N__29816));
    IoInMux I__7089 (
            .O(N__29835),
            .I(N__29813));
    LocalMux I__7088 (
            .O(N__29832),
            .I(N__29809));
    LocalMux I__7087 (
            .O(N__29829),
            .I(N__29804));
    LocalMux I__7086 (
            .O(N__29826),
            .I(N__29804));
    Span4Mux_s3_v I__7085 (
            .O(N__29823),
            .I(N__29799));
    LocalMux I__7084 (
            .O(N__29820),
            .I(N__29799));
    SRMux I__7083 (
            .O(N__29819),
            .I(N__29796));
    LocalMux I__7082 (
            .O(N__29816),
            .I(N__29791));
    LocalMux I__7081 (
            .O(N__29813),
            .I(N__29784));
    SRMux I__7080 (
            .O(N__29812),
            .I(N__29781));
    Span4Mux_s3_h I__7079 (
            .O(N__29809),
            .I(N__29775));
    Span4Mux_v I__7078 (
            .O(N__29804),
            .I(N__29768));
    Span4Mux_v I__7077 (
            .O(N__29799),
            .I(N__29768));
    LocalMux I__7076 (
            .O(N__29796),
            .I(N__29768));
    SRMux I__7075 (
            .O(N__29795),
            .I(N__29765));
    SRMux I__7074 (
            .O(N__29794),
            .I(N__29762));
    Span4Mux_v I__7073 (
            .O(N__29791),
            .I(N__29759));
    SRMux I__7072 (
            .O(N__29790),
            .I(N__29756));
    SRMux I__7071 (
            .O(N__29789),
            .I(N__29748));
    SRMux I__7070 (
            .O(N__29788),
            .I(N__29745));
    SRMux I__7069 (
            .O(N__29787),
            .I(N__29740));
    IoSpan4Mux I__7068 (
            .O(N__29784),
            .I(N__29736));
    LocalMux I__7067 (
            .O(N__29781),
            .I(N__29732));
    SRMux I__7066 (
            .O(N__29780),
            .I(N__29729));
    SRMux I__7065 (
            .O(N__29779),
            .I(N__29726));
    SRMux I__7064 (
            .O(N__29778),
            .I(N__29722));
    Span4Mux_h I__7063 (
            .O(N__29775),
            .I(N__29711));
    Span4Mux_v I__7062 (
            .O(N__29768),
            .I(N__29711));
    LocalMux I__7061 (
            .O(N__29765),
            .I(N__29711));
    LocalMux I__7060 (
            .O(N__29762),
            .I(N__29711));
    Span4Mux_v I__7059 (
            .O(N__29759),
            .I(N__29706));
    LocalMux I__7058 (
            .O(N__29756),
            .I(N__29706));
    SRMux I__7057 (
            .O(N__29755),
            .I(N__29703));
    SRMux I__7056 (
            .O(N__29754),
            .I(N__29699));
    CascadeMux I__7055 (
            .O(N__29753),
            .I(N__29695));
    CascadeMux I__7054 (
            .O(N__29752),
            .I(N__29692));
    CascadeMux I__7053 (
            .O(N__29751),
            .I(N__29686));
    LocalMux I__7052 (
            .O(N__29748),
            .I(N__29671));
    LocalMux I__7051 (
            .O(N__29745),
            .I(N__29671));
    SRMux I__7050 (
            .O(N__29744),
            .I(N__29668));
    SRMux I__7049 (
            .O(N__29743),
            .I(N__29665));
    LocalMux I__7048 (
            .O(N__29740),
            .I(N__29661));
    SRMux I__7047 (
            .O(N__29739),
            .I(N__29658));
    Span4Mux_s2_h I__7046 (
            .O(N__29736),
            .I(N__29655));
    SRMux I__7045 (
            .O(N__29735),
            .I(N__29652));
    Span4Mux_h I__7044 (
            .O(N__29732),
            .I(N__29643));
    LocalMux I__7043 (
            .O(N__29729),
            .I(N__29643));
    LocalMux I__7042 (
            .O(N__29726),
            .I(N__29643));
    SRMux I__7041 (
            .O(N__29725),
            .I(N__29640));
    LocalMux I__7040 (
            .O(N__29722),
            .I(N__29637));
    SRMux I__7039 (
            .O(N__29721),
            .I(N__29634));
    SRMux I__7038 (
            .O(N__29720),
            .I(N__29631));
    Span4Mux_v I__7037 (
            .O(N__29711),
            .I(N__29625));
    Span4Mux_v I__7036 (
            .O(N__29706),
            .I(N__29620));
    LocalMux I__7035 (
            .O(N__29703),
            .I(N__29620));
    SRMux I__7034 (
            .O(N__29702),
            .I(N__29617));
    LocalMux I__7033 (
            .O(N__29699),
            .I(N__29614));
    InMux I__7032 (
            .O(N__29698),
            .I(N__29599));
    InMux I__7031 (
            .O(N__29695),
            .I(N__29599));
    InMux I__7030 (
            .O(N__29692),
            .I(N__29599));
    InMux I__7029 (
            .O(N__29691),
            .I(N__29599));
    InMux I__7028 (
            .O(N__29690),
            .I(N__29599));
    InMux I__7027 (
            .O(N__29689),
            .I(N__29599));
    InMux I__7026 (
            .O(N__29686),
            .I(N__29599));
    CascadeMux I__7025 (
            .O(N__29685),
            .I(N__29596));
    CascadeMux I__7024 (
            .O(N__29684),
            .I(N__29593));
    CascadeMux I__7023 (
            .O(N__29683),
            .I(N__29590));
    CascadeMux I__7022 (
            .O(N__29682),
            .I(N__29587));
    CascadeMux I__7021 (
            .O(N__29681),
            .I(N__29584));
    CascadeMux I__7020 (
            .O(N__29680),
            .I(N__29581));
    CascadeMux I__7019 (
            .O(N__29679),
            .I(N__29578));
    CascadeMux I__7018 (
            .O(N__29678),
            .I(N__29574));
    CascadeMux I__7017 (
            .O(N__29677),
            .I(N__29570));
    CascadeMux I__7016 (
            .O(N__29676),
            .I(N__29566));
    Span4Mux_s3_v I__7015 (
            .O(N__29671),
            .I(N__29559));
    LocalMux I__7014 (
            .O(N__29668),
            .I(N__29559));
    LocalMux I__7013 (
            .O(N__29665),
            .I(N__29559));
    SRMux I__7012 (
            .O(N__29664),
            .I(N__29556));
    Span4Mux_s3_v I__7011 (
            .O(N__29661),
            .I(N__29551));
    LocalMux I__7010 (
            .O(N__29658),
            .I(N__29551));
    Span4Mux_h I__7009 (
            .O(N__29655),
            .I(N__29546));
    LocalMux I__7008 (
            .O(N__29652),
            .I(N__29546));
    SRMux I__7007 (
            .O(N__29651),
            .I(N__29543));
    SRMux I__7006 (
            .O(N__29650),
            .I(N__29540));
    Span4Mux_v I__7005 (
            .O(N__29643),
            .I(N__29534));
    LocalMux I__7004 (
            .O(N__29640),
            .I(N__29534));
    Span4Mux_v I__7003 (
            .O(N__29637),
            .I(N__29527));
    LocalMux I__7002 (
            .O(N__29634),
            .I(N__29527));
    LocalMux I__7001 (
            .O(N__29631),
            .I(N__29527));
    SRMux I__7000 (
            .O(N__29630),
            .I(N__29524));
    SRMux I__6999 (
            .O(N__29629),
            .I(N__29521));
    SRMux I__6998 (
            .O(N__29628),
            .I(N__29516));
    Span4Mux_h I__6997 (
            .O(N__29625),
            .I(N__29505));
    Span4Mux_h I__6996 (
            .O(N__29620),
            .I(N__29505));
    LocalMux I__6995 (
            .O(N__29617),
            .I(N__29502));
    Span4Mux_h I__6994 (
            .O(N__29614),
            .I(N__29497));
    LocalMux I__6993 (
            .O(N__29599),
            .I(N__29497));
    InMux I__6992 (
            .O(N__29596),
            .I(N__29488));
    InMux I__6991 (
            .O(N__29593),
            .I(N__29488));
    InMux I__6990 (
            .O(N__29590),
            .I(N__29488));
    InMux I__6989 (
            .O(N__29587),
            .I(N__29488));
    InMux I__6988 (
            .O(N__29584),
            .I(N__29481));
    InMux I__6987 (
            .O(N__29581),
            .I(N__29481));
    InMux I__6986 (
            .O(N__29578),
            .I(N__29481));
    InMux I__6985 (
            .O(N__29577),
            .I(N__29468));
    InMux I__6984 (
            .O(N__29574),
            .I(N__29468));
    InMux I__6983 (
            .O(N__29573),
            .I(N__29468));
    InMux I__6982 (
            .O(N__29570),
            .I(N__29468));
    InMux I__6981 (
            .O(N__29569),
            .I(N__29468));
    InMux I__6980 (
            .O(N__29566),
            .I(N__29468));
    Span4Mux_v I__6979 (
            .O(N__29559),
            .I(N__29463));
    LocalMux I__6978 (
            .O(N__29556),
            .I(N__29463));
    Span4Mux_v I__6977 (
            .O(N__29551),
            .I(N__29454));
    Span4Mux_h I__6976 (
            .O(N__29546),
            .I(N__29454));
    LocalMux I__6975 (
            .O(N__29543),
            .I(N__29454));
    LocalMux I__6974 (
            .O(N__29540),
            .I(N__29454));
    SRMux I__6973 (
            .O(N__29539),
            .I(N__29451));
    Span4Mux_v I__6972 (
            .O(N__29534),
            .I(N__29442));
    Span4Mux_v I__6971 (
            .O(N__29527),
            .I(N__29442));
    LocalMux I__6970 (
            .O(N__29524),
            .I(N__29442));
    LocalMux I__6969 (
            .O(N__29521),
            .I(N__29442));
    SRMux I__6968 (
            .O(N__29520),
            .I(N__29439));
    SRMux I__6967 (
            .O(N__29519),
            .I(N__29436));
    LocalMux I__6966 (
            .O(N__29516),
            .I(N__29433));
    SRMux I__6965 (
            .O(N__29515),
            .I(N__29430));
    SRMux I__6964 (
            .O(N__29514),
            .I(N__29427));
    SRMux I__6963 (
            .O(N__29513),
            .I(N__29423));
    SRMux I__6962 (
            .O(N__29512),
            .I(N__29420));
    SRMux I__6961 (
            .O(N__29511),
            .I(N__29417));
    SRMux I__6960 (
            .O(N__29510),
            .I(N__29414));
    Span4Mux_h I__6959 (
            .O(N__29505),
            .I(N__29411));
    Span4Mux_h I__6958 (
            .O(N__29502),
            .I(N__29402));
    Span4Mux_v I__6957 (
            .O(N__29497),
            .I(N__29402));
    LocalMux I__6956 (
            .O(N__29488),
            .I(N__29402));
    LocalMux I__6955 (
            .O(N__29481),
            .I(N__29402));
    LocalMux I__6954 (
            .O(N__29468),
            .I(N__29399));
    Span4Mux_v I__6953 (
            .O(N__29463),
            .I(N__29392));
    Span4Mux_v I__6952 (
            .O(N__29454),
            .I(N__29392));
    LocalMux I__6951 (
            .O(N__29451),
            .I(N__29392));
    Span4Mux_v I__6950 (
            .O(N__29442),
            .I(N__29385));
    LocalMux I__6949 (
            .O(N__29439),
            .I(N__29385));
    LocalMux I__6948 (
            .O(N__29436),
            .I(N__29385));
    Span4Mux_v I__6947 (
            .O(N__29433),
            .I(N__29378));
    LocalMux I__6946 (
            .O(N__29430),
            .I(N__29378));
    LocalMux I__6945 (
            .O(N__29427),
            .I(N__29378));
    SRMux I__6944 (
            .O(N__29426),
            .I(N__29375));
    LocalMux I__6943 (
            .O(N__29423),
            .I(N__29370));
    LocalMux I__6942 (
            .O(N__29420),
            .I(N__29370));
    LocalMux I__6941 (
            .O(N__29417),
            .I(N__29367));
    LocalMux I__6940 (
            .O(N__29414),
            .I(N__29364));
    Span4Mux_h I__6939 (
            .O(N__29411),
            .I(N__29359));
    Span4Mux_v I__6938 (
            .O(N__29402),
            .I(N__29359));
    Span4Mux_v I__6937 (
            .O(N__29399),
            .I(N__29356));
    Span4Mux_v I__6936 (
            .O(N__29392),
            .I(N__29351));
    Span4Mux_v I__6935 (
            .O(N__29385),
            .I(N__29351));
    Span4Mux_v I__6934 (
            .O(N__29378),
            .I(N__29344));
    LocalMux I__6933 (
            .O(N__29375),
            .I(N__29344));
    Span4Mux_v I__6932 (
            .O(N__29370),
            .I(N__29344));
    Span12Mux_h I__6931 (
            .O(N__29367),
            .I(N__29341));
    Span12Mux_h I__6930 (
            .O(N__29364),
            .I(N__29338));
    Span4Mux_h I__6929 (
            .O(N__29359),
            .I(N__29335));
    Span4Mux_h I__6928 (
            .O(N__29356),
            .I(N__29328));
    Span4Mux_h I__6927 (
            .O(N__29351),
            .I(N__29328));
    Span4Mux_h I__6926 (
            .O(N__29344),
            .I(N__29328));
    Odrv12 I__6925 (
            .O(N__29341),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__6924 (
            .O(N__29338),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6923 (
            .O(N__29335),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6922 (
            .O(N__29328),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__6921 (
            .O(N__29319),
            .I(N__29316));
    InMux I__6920 (
            .O(N__29316),
            .I(N__29312));
    InMux I__6919 (
            .O(N__29315),
            .I(N__29309));
    LocalMux I__6918 (
            .O(N__29312),
            .I(N__29304));
    LocalMux I__6917 (
            .O(N__29309),
            .I(N__29304));
    Span4Mux_h I__6916 (
            .O(N__29304),
            .I(N__29301));
    Span4Mux_v I__6915 (
            .O(N__29301),
            .I(N__29298));
    Odrv4 I__6914 (
            .O(N__29298),
            .I(M_this_data_count_qZ0Z_14));
    InMux I__6913 (
            .O(N__29295),
            .I(N__29292));
    LocalMux I__6912 (
            .O(N__29292),
            .I(N__29289));
    Span4Mux_h I__6911 (
            .O(N__29289),
            .I(N__29286));
    Span4Mux_v I__6910 (
            .O(N__29286),
            .I(N__29283));
    Span4Mux_h I__6909 (
            .O(N__29283),
            .I(N__29280));
    Odrv4 I__6908 (
            .O(N__29280),
            .I(M_this_data_count_q_s_14));
    InMux I__6907 (
            .O(N__29277),
            .I(M_this_data_count_q_cry_13));
    CascadeMux I__6906 (
            .O(N__29274),
            .I(N__29270));
    InMux I__6905 (
            .O(N__29273),
            .I(N__29267));
    InMux I__6904 (
            .O(N__29270),
            .I(N__29264));
    LocalMux I__6903 (
            .O(N__29267),
            .I(M_this_data_count_qZ0Z_15));
    LocalMux I__6902 (
            .O(N__29264),
            .I(M_this_data_count_qZ0Z_15));
    InMux I__6901 (
            .O(N__29259),
            .I(M_this_data_count_q_cry_14));
    InMux I__6900 (
            .O(N__29256),
            .I(N__29253));
    LocalMux I__6899 (
            .O(N__29253),
            .I(N__29250));
    Odrv4 I__6898 (
            .O(N__29250),
            .I(M_this_data_count_q_s_15));
    InMux I__6897 (
            .O(N__29247),
            .I(N__29244));
    LocalMux I__6896 (
            .O(N__29244),
            .I(N__29241));
    Odrv4 I__6895 (
            .O(N__29241),
            .I(M_this_data_count_q_cry_3_THRU_CO));
    CascadeMux I__6894 (
            .O(N__29238),
            .I(N__29228));
    InMux I__6893 (
            .O(N__29237),
            .I(N__29220));
    InMux I__6892 (
            .O(N__29236),
            .I(N__29220));
    InMux I__6891 (
            .O(N__29235),
            .I(N__29213));
    InMux I__6890 (
            .O(N__29234),
            .I(N__29213));
    InMux I__6889 (
            .O(N__29233),
            .I(N__29213));
    InMux I__6888 (
            .O(N__29232),
            .I(N__29209));
    InMux I__6887 (
            .O(N__29231),
            .I(N__29202));
    InMux I__6886 (
            .O(N__29228),
            .I(N__29202));
    InMux I__6885 (
            .O(N__29227),
            .I(N__29202));
    InMux I__6884 (
            .O(N__29226),
            .I(N__29197));
    InMux I__6883 (
            .O(N__29225),
            .I(N__29197));
    LocalMux I__6882 (
            .O(N__29220),
            .I(N__29189));
    LocalMux I__6881 (
            .O(N__29213),
            .I(N__29189));
    InMux I__6880 (
            .O(N__29212),
            .I(N__29185));
    LocalMux I__6879 (
            .O(N__29209),
            .I(N__29182));
    LocalMux I__6878 (
            .O(N__29202),
            .I(N__29177));
    LocalMux I__6877 (
            .O(N__29197),
            .I(N__29177));
    InMux I__6876 (
            .O(N__29196),
            .I(N__29170));
    InMux I__6875 (
            .O(N__29195),
            .I(N__29170));
    InMux I__6874 (
            .O(N__29194),
            .I(N__29170));
    Span4Mux_h I__6873 (
            .O(N__29189),
            .I(N__29167));
    InMux I__6872 (
            .O(N__29188),
            .I(N__29164));
    LocalMux I__6871 (
            .O(N__29185),
            .I(N__29161));
    Span4Mux_v I__6870 (
            .O(N__29182),
            .I(N__29154));
    Span4Mux_v I__6869 (
            .O(N__29177),
            .I(N__29154));
    LocalMux I__6868 (
            .O(N__29170),
            .I(N__29154));
    Span4Mux_v I__6867 (
            .O(N__29167),
            .I(N__29151));
    LocalMux I__6866 (
            .O(N__29164),
            .I(N__29148));
    Span4Mux_h I__6865 (
            .O(N__29161),
            .I(N__29143));
    Span4Mux_h I__6864 (
            .O(N__29154),
            .I(N__29143));
    Odrv4 I__6863 (
            .O(N__29151),
            .I(N_33));
    Odrv12 I__6862 (
            .O(N__29148),
            .I(N_33));
    Odrv4 I__6861 (
            .O(N__29143),
            .I(N_33));
    InMux I__6860 (
            .O(N__29136),
            .I(N__29132));
    InMux I__6859 (
            .O(N__29135),
            .I(N__29128));
    LocalMux I__6858 (
            .O(N__29132),
            .I(N__29125));
    InMux I__6857 (
            .O(N__29131),
            .I(N__29122));
    LocalMux I__6856 (
            .O(N__29128),
            .I(N__29119));
    Span4Mux_h I__6855 (
            .O(N__29125),
            .I(N__29116));
    LocalMux I__6854 (
            .O(N__29122),
            .I(M_this_data_count_qZ0Z_4));
    Odrv4 I__6853 (
            .O(N__29119),
            .I(M_this_data_count_qZ0Z_4));
    Odrv4 I__6852 (
            .O(N__29116),
            .I(M_this_data_count_qZ0Z_4));
    CEMux I__6851 (
            .O(N__29109),
            .I(N__29105));
    CEMux I__6850 (
            .O(N__29108),
            .I(N__29098));
    LocalMux I__6849 (
            .O(N__29105),
            .I(N__29095));
    CEMux I__6848 (
            .O(N__29104),
            .I(N__29092));
    CEMux I__6847 (
            .O(N__29103),
            .I(N__29089));
    CEMux I__6846 (
            .O(N__29102),
            .I(N__29086));
    CEMux I__6845 (
            .O(N__29101),
            .I(N__29082));
    LocalMux I__6844 (
            .O(N__29098),
            .I(N__29078));
    Span4Mux_h I__6843 (
            .O(N__29095),
            .I(N__29073));
    LocalMux I__6842 (
            .O(N__29092),
            .I(N__29073));
    LocalMux I__6841 (
            .O(N__29089),
            .I(N__29070));
    LocalMux I__6840 (
            .O(N__29086),
            .I(N__29067));
    CEMux I__6839 (
            .O(N__29085),
            .I(N__29064));
    LocalMux I__6838 (
            .O(N__29082),
            .I(N__29061));
    CEMux I__6837 (
            .O(N__29081),
            .I(N__29058));
    Span4Mux_v I__6836 (
            .O(N__29078),
            .I(N__29053));
    Span4Mux_v I__6835 (
            .O(N__29073),
            .I(N__29053));
    Span4Mux_h I__6834 (
            .O(N__29070),
            .I(N__29050));
    Span4Mux_h I__6833 (
            .O(N__29067),
            .I(N__29045));
    LocalMux I__6832 (
            .O(N__29064),
            .I(N__29045));
    Span4Mux_v I__6831 (
            .O(N__29061),
            .I(N__29042));
    LocalMux I__6830 (
            .O(N__29058),
            .I(N__29039));
    Span4Mux_h I__6829 (
            .O(N__29053),
            .I(N__29036));
    Odrv4 I__6828 (
            .O(N__29050),
            .I(N_35));
    Odrv4 I__6827 (
            .O(N__29045),
            .I(N_35));
    Odrv4 I__6826 (
            .O(N__29042),
            .I(N_35));
    Odrv4 I__6825 (
            .O(N__29039),
            .I(N_35));
    Odrv4 I__6824 (
            .O(N__29036),
            .I(N_35));
    InMux I__6823 (
            .O(N__29025),
            .I(M_this_data_count_q_cry_0));
    InMux I__6822 (
            .O(N__29022),
            .I(N__29017));
    InMux I__6821 (
            .O(N__29021),
            .I(N__29012));
    InMux I__6820 (
            .O(N__29020),
            .I(N__29012));
    LocalMux I__6819 (
            .O(N__29017),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__6818 (
            .O(N__29012),
            .I(M_this_data_count_qZ0Z_2));
    InMux I__6817 (
            .O(N__29007),
            .I(N__29004));
    LocalMux I__6816 (
            .O(N__29004),
            .I(N__29001));
    Odrv4 I__6815 (
            .O(N__29001),
            .I(M_this_data_count_q_cry_1_THRU_CO));
    InMux I__6814 (
            .O(N__28998),
            .I(M_this_data_count_q_cry_1));
    CascadeMux I__6813 (
            .O(N__28995),
            .I(N__28991));
    InMux I__6812 (
            .O(N__28994),
            .I(N__28988));
    InMux I__6811 (
            .O(N__28991),
            .I(N__28985));
    LocalMux I__6810 (
            .O(N__28988),
            .I(N__28980));
    LocalMux I__6809 (
            .O(N__28985),
            .I(N__28980));
    Span4Mux_h I__6808 (
            .O(N__28980),
            .I(N__28976));
    InMux I__6807 (
            .O(N__28979),
            .I(N__28973));
    Span4Mux_v I__6806 (
            .O(N__28976),
            .I(N__28970));
    LocalMux I__6805 (
            .O(N__28973),
            .I(M_this_data_count_qZ0Z_3));
    Odrv4 I__6804 (
            .O(N__28970),
            .I(M_this_data_count_qZ0Z_3));
    InMux I__6803 (
            .O(N__28965),
            .I(N__28962));
    LocalMux I__6802 (
            .O(N__28962),
            .I(N__28959));
    Span4Mux_h I__6801 (
            .O(N__28959),
            .I(N__28956));
    Span4Mux_h I__6800 (
            .O(N__28956),
            .I(N__28953));
    Odrv4 I__6799 (
            .O(N__28953),
            .I(M_this_data_count_q_cry_2_THRU_CO));
    InMux I__6798 (
            .O(N__28950),
            .I(M_this_data_count_q_cry_2));
    InMux I__6797 (
            .O(N__28947),
            .I(M_this_data_count_q_cry_3));
    InMux I__6796 (
            .O(N__28944),
            .I(N__28941));
    LocalMux I__6795 (
            .O(N__28941),
            .I(N__28936));
    InMux I__6794 (
            .O(N__28940),
            .I(N__28931));
    InMux I__6793 (
            .O(N__28939),
            .I(N__28931));
    Odrv4 I__6792 (
            .O(N__28936),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__6791 (
            .O(N__28931),
            .I(M_this_data_count_qZ0Z_5));
    InMux I__6790 (
            .O(N__28926),
            .I(N__28923));
    LocalMux I__6789 (
            .O(N__28923),
            .I(N__28920));
    Odrv4 I__6788 (
            .O(N__28920),
            .I(M_this_data_count_q_cry_4_THRU_CO));
    InMux I__6787 (
            .O(N__28917),
            .I(M_this_data_count_q_cry_4));
    InMux I__6786 (
            .O(N__28914),
            .I(N__28911));
    LocalMux I__6785 (
            .O(N__28911),
            .I(N__28907));
    InMux I__6784 (
            .O(N__28910),
            .I(N__28904));
    Odrv4 I__6783 (
            .O(N__28907),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__6782 (
            .O(N__28904),
            .I(M_this_data_count_qZ0Z_6));
    InMux I__6781 (
            .O(N__28899),
            .I(N__28896));
    LocalMux I__6780 (
            .O(N__28896),
            .I(N__28893));
    Odrv12 I__6779 (
            .O(N__28893),
            .I(M_this_data_count_q_s_6));
    InMux I__6778 (
            .O(N__28890),
            .I(M_this_data_count_q_cry_5));
    InMux I__6777 (
            .O(N__28887),
            .I(N__28883));
    CascadeMux I__6776 (
            .O(N__28886),
            .I(N__28879));
    LocalMux I__6775 (
            .O(N__28883),
            .I(N__28876));
    InMux I__6774 (
            .O(N__28882),
            .I(N__28871));
    InMux I__6773 (
            .O(N__28879),
            .I(N__28871));
    Odrv4 I__6772 (
            .O(N__28876),
            .I(M_this_data_count_qZ0Z_7));
    LocalMux I__6771 (
            .O(N__28871),
            .I(M_this_data_count_qZ0Z_7));
    InMux I__6770 (
            .O(N__28866),
            .I(N__28863));
    LocalMux I__6769 (
            .O(N__28863),
            .I(N__28860));
    Odrv4 I__6768 (
            .O(N__28860),
            .I(M_this_data_count_q_cry_6_THRU_CO));
    InMux I__6767 (
            .O(N__28857),
            .I(M_this_data_count_q_cry_6));
    CascadeMux I__6766 (
            .O(N__28854),
            .I(N__28851));
    InMux I__6765 (
            .O(N__28851),
            .I(N__28848));
    LocalMux I__6764 (
            .O(N__28848),
            .I(N__28845));
    Span4Mux_v I__6763 (
            .O(N__28845),
            .I(N__28841));
    InMux I__6762 (
            .O(N__28844),
            .I(N__28838));
    Odrv4 I__6761 (
            .O(N__28841),
            .I(M_this_data_count_qZ0Z_8));
    LocalMux I__6760 (
            .O(N__28838),
            .I(M_this_data_count_qZ0Z_8));
    InMux I__6759 (
            .O(N__28833),
            .I(N__28830));
    LocalMux I__6758 (
            .O(N__28830),
            .I(N__28827));
    Odrv4 I__6757 (
            .O(N__28827),
            .I(M_this_data_count_q_s_8));
    InMux I__6756 (
            .O(N__28824),
            .I(bfn_24_22_0_));
    InMux I__6755 (
            .O(N__28821),
            .I(N__28818));
    LocalMux I__6754 (
            .O(N__28818),
            .I(N__28814));
    InMux I__6753 (
            .O(N__28817),
            .I(N__28811));
    Odrv4 I__6752 (
            .O(N__28814),
            .I(M_this_data_count_qZ0Z_9));
    LocalMux I__6751 (
            .O(N__28811),
            .I(M_this_data_count_qZ0Z_9));
    InMux I__6750 (
            .O(N__28806),
            .I(N__28803));
    LocalMux I__6749 (
            .O(N__28803),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ));
    CascadeMux I__6748 (
            .O(N__28800),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ));
    InMux I__6747 (
            .O(N__28797),
            .I(N__28794));
    LocalMux I__6746 (
            .O(N__28794),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ));
    InMux I__6745 (
            .O(N__28791),
            .I(N__28787));
    InMux I__6744 (
            .O(N__28790),
            .I(N__28784));
    LocalMux I__6743 (
            .O(N__28787),
            .I(N__28780));
    LocalMux I__6742 (
            .O(N__28784),
            .I(N__28777));
    InMux I__6741 (
            .O(N__28783),
            .I(N__28774));
    Span4Mux_v I__6740 (
            .O(N__28780),
            .I(N__28771));
    Span12Mux_s11_h I__6739 (
            .O(N__28777),
            .I(N__28766));
    LocalMux I__6738 (
            .O(N__28774),
            .I(N__28766));
    Sp12to4 I__6737 (
            .O(N__28771),
            .I(N__28761));
    Span12Mux_v I__6736 (
            .O(N__28766),
            .I(N__28761));
    Span12Mux_h I__6735 (
            .O(N__28761),
            .I(N__28758));
    Odrv12 I__6734 (
            .O(N__28758),
            .I(M_this_ppu_vram_data_3));
    InMux I__6733 (
            .O(N__28755),
            .I(N__28752));
    LocalMux I__6732 (
            .O(N__28752),
            .I(N__28749));
    Span4Mux_v I__6731 (
            .O(N__28749),
            .I(N__28746));
    Odrv4 I__6730 (
            .O(N__28746),
            .I(\this_sprites_ram.mem_out_bus6_0 ));
    InMux I__6729 (
            .O(N__28743),
            .I(N__28740));
    LocalMux I__6728 (
            .O(N__28740),
            .I(N__28737));
    Span4Mux_v I__6727 (
            .O(N__28737),
            .I(N__28734));
    Span4Mux_v I__6726 (
            .O(N__28734),
            .I(N__28731));
    Odrv4 I__6725 (
            .O(N__28731),
            .I(\this_sprites_ram.mem_out_bus2_0 ));
    CascadeMux I__6724 (
            .O(N__28728),
            .I(N__28724));
    InMux I__6723 (
            .O(N__28727),
            .I(N__28721));
    InMux I__6722 (
            .O(N__28724),
            .I(N__28716));
    LocalMux I__6721 (
            .O(N__28721),
            .I(N__28713));
    InMux I__6720 (
            .O(N__28720),
            .I(N__28710));
    InMux I__6719 (
            .O(N__28719),
            .I(N__28707));
    LocalMux I__6718 (
            .O(N__28716),
            .I(N__28702));
    Span4Mux_v I__6717 (
            .O(N__28713),
            .I(N__28702));
    LocalMux I__6716 (
            .O(N__28710),
            .I(N__28699));
    LocalMux I__6715 (
            .O(N__28707),
            .I(N__28692));
    Span4Mux_h I__6714 (
            .O(N__28702),
            .I(N__28692));
    Span4Mux_h I__6713 (
            .O(N__28699),
            .I(N__28692));
    Span4Mux_h I__6712 (
            .O(N__28692),
            .I(N__28689));
    Odrv4 I__6711 (
            .O(N__28689),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    InMux I__6710 (
            .O(N__28686),
            .I(N__28683));
    LocalMux I__6709 (
            .O(N__28683),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ));
    CascadeMux I__6708 (
            .O(N__28680),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0_cascade_ ));
    CascadeMux I__6707 (
            .O(N__28677),
            .I(N__28673));
    InMux I__6706 (
            .O(N__28676),
            .I(N__28670));
    InMux I__6705 (
            .O(N__28673),
            .I(N__28663));
    LocalMux I__6704 (
            .O(N__28670),
            .I(N__28658));
    InMux I__6703 (
            .O(N__28669),
            .I(N__28653));
    InMux I__6702 (
            .O(N__28668),
            .I(N__28653));
    InMux I__6701 (
            .O(N__28667),
            .I(N__28648));
    InMux I__6700 (
            .O(N__28666),
            .I(N__28648));
    LocalMux I__6699 (
            .O(N__28663),
            .I(N__28645));
    InMux I__6698 (
            .O(N__28662),
            .I(N__28640));
    InMux I__6697 (
            .O(N__28661),
            .I(N__28640));
    Sp12to4 I__6696 (
            .O(N__28658),
            .I(N__28633));
    LocalMux I__6695 (
            .O(N__28653),
            .I(N__28633));
    LocalMux I__6694 (
            .O(N__28648),
            .I(N__28633));
    Odrv12 I__6693 (
            .O(N__28645),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    LocalMux I__6692 (
            .O(N__28640),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    Odrv12 I__6691 (
            .O(N__28633),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    InMux I__6690 (
            .O(N__28626),
            .I(N__28623));
    LocalMux I__6689 (
            .O(N__28623),
            .I(N__28620));
    Span12Mux_h I__6688 (
            .O(N__28620),
            .I(N__28617));
    Odrv12 I__6687 (
            .O(N__28617),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ));
    InMux I__6686 (
            .O(N__28614),
            .I(N__28611));
    LocalMux I__6685 (
            .O(N__28611),
            .I(N__28608));
    Sp12to4 I__6684 (
            .O(N__28608),
            .I(N__28605));
    Odrv12 I__6683 (
            .O(N__28605),
            .I(\this_sprites_ram.mem_out_bus6_2 ));
    InMux I__6682 (
            .O(N__28602),
            .I(N__28599));
    LocalMux I__6681 (
            .O(N__28599),
            .I(N__28596));
    Span4Mux_v I__6680 (
            .O(N__28596),
            .I(N__28593));
    Span4Mux_v I__6679 (
            .O(N__28593),
            .I(N__28590));
    Odrv4 I__6678 (
            .O(N__28590),
            .I(\this_sprites_ram.mem_out_bus2_2 ));
    InMux I__6677 (
            .O(N__28587),
            .I(N__28584));
    LocalMux I__6676 (
            .O(N__28584),
            .I(N__28581));
    Span4Mux_v I__6675 (
            .O(N__28581),
            .I(N__28578));
    Span4Mux_h I__6674 (
            .O(N__28578),
            .I(N__28575));
    Odrv4 I__6673 (
            .O(N__28575),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ));
    CEMux I__6672 (
            .O(N__28572),
            .I(N__28568));
    CEMux I__6671 (
            .O(N__28571),
            .I(N__28565));
    LocalMux I__6670 (
            .O(N__28568),
            .I(N__28560));
    LocalMux I__6669 (
            .O(N__28565),
            .I(N__28560));
    Span4Mux_v I__6668 (
            .O(N__28560),
            .I(N__28557));
    Odrv4 I__6667 (
            .O(N__28557),
            .I(\this_sprites_ram.mem_WE_4 ));
    InMux I__6666 (
            .O(N__28554),
            .I(N__28551));
    LocalMux I__6665 (
            .O(N__28551),
            .I(N__28548));
    Span4Mux_v I__6664 (
            .O(N__28548),
            .I(N__28545));
    Span4Mux_v I__6663 (
            .O(N__28545),
            .I(N__28542));
    Odrv4 I__6662 (
            .O(N__28542),
            .I(\this_sprites_ram.mem_out_bus7_0 ));
    InMux I__6661 (
            .O(N__28539),
            .I(N__28536));
    LocalMux I__6660 (
            .O(N__28536),
            .I(N__28533));
    Span4Mux_v I__6659 (
            .O(N__28533),
            .I(N__28530));
    Odrv4 I__6658 (
            .O(N__28530),
            .I(\this_sprites_ram.mem_out_bus3_0 ));
    InMux I__6657 (
            .O(N__28527),
            .I(N__28524));
    LocalMux I__6656 (
            .O(N__28524),
            .I(N__28521));
    Span12Mux_v I__6655 (
            .O(N__28521),
            .I(N__28518));
    Span12Mux_h I__6654 (
            .O(N__28518),
            .I(N__28515));
    Odrv12 I__6653 (
            .O(N__28515),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ));
    InMux I__6652 (
            .O(N__28512),
            .I(N__28507));
    InMux I__6651 (
            .O(N__28511),
            .I(N__28504));
    InMux I__6650 (
            .O(N__28510),
            .I(N__28501));
    LocalMux I__6649 (
            .O(N__28507),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__6648 (
            .O(N__28504),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__6647 (
            .O(N__28501),
            .I(M_this_data_count_qZ0Z_0));
    InMux I__6646 (
            .O(N__28494),
            .I(N__28489));
    InMux I__6645 (
            .O(N__28493),
            .I(N__28484));
    InMux I__6644 (
            .O(N__28492),
            .I(N__28484));
    LocalMux I__6643 (
            .O(N__28489),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__6642 (
            .O(N__28484),
            .I(M_this_data_count_qZ0Z_1));
    InMux I__6641 (
            .O(N__28479),
            .I(N__28476));
    LocalMux I__6640 (
            .O(N__28476),
            .I(M_this_data_count_q_cry_0_THRU_CO));
    InMux I__6639 (
            .O(N__28473),
            .I(N__28465));
    InMux I__6638 (
            .O(N__28472),
            .I(N__28462));
    InMux I__6637 (
            .O(N__28471),
            .I(N__28459));
    CascadeMux I__6636 (
            .O(N__28470),
            .I(N__28456));
    InMux I__6635 (
            .O(N__28469),
            .I(N__28451));
    InMux I__6634 (
            .O(N__28468),
            .I(N__28448));
    LocalMux I__6633 (
            .O(N__28465),
            .I(N__28444));
    LocalMux I__6632 (
            .O(N__28462),
            .I(N__28441));
    LocalMux I__6631 (
            .O(N__28459),
            .I(N__28438));
    InMux I__6630 (
            .O(N__28456),
            .I(N__28435));
    CascadeMux I__6629 (
            .O(N__28455),
            .I(N__28432));
    InMux I__6628 (
            .O(N__28454),
            .I(N__28429));
    LocalMux I__6627 (
            .O(N__28451),
            .I(N__28426));
    LocalMux I__6626 (
            .O(N__28448),
            .I(N__28423));
    InMux I__6625 (
            .O(N__28447),
            .I(N__28420));
    Span4Mux_v I__6624 (
            .O(N__28444),
            .I(N__28416));
    Span4Mux_v I__6623 (
            .O(N__28441),
            .I(N__28409));
    Span4Mux_v I__6622 (
            .O(N__28438),
            .I(N__28409));
    LocalMux I__6621 (
            .O(N__28435),
            .I(N__28409));
    InMux I__6620 (
            .O(N__28432),
            .I(N__28406));
    LocalMux I__6619 (
            .O(N__28429),
            .I(N__28403));
    Span4Mux_v I__6618 (
            .O(N__28426),
            .I(N__28396));
    Span4Mux_v I__6617 (
            .O(N__28423),
            .I(N__28396));
    LocalMux I__6616 (
            .O(N__28420),
            .I(N__28396));
    InMux I__6615 (
            .O(N__28419),
            .I(N__28392));
    Span4Mux_v I__6614 (
            .O(N__28416),
            .I(N__28389));
    Span4Mux_v I__6613 (
            .O(N__28409),
            .I(N__28386));
    LocalMux I__6612 (
            .O(N__28406),
            .I(N__28383));
    Span4Mux_v I__6611 (
            .O(N__28403),
            .I(N__28378));
    Span4Mux_h I__6610 (
            .O(N__28396),
            .I(N__28378));
    InMux I__6609 (
            .O(N__28395),
            .I(N__28375));
    LocalMux I__6608 (
            .O(N__28392),
            .I(N__28372));
    Span4Mux_v I__6607 (
            .O(N__28389),
            .I(N__28369));
    Span4Mux_v I__6606 (
            .O(N__28386),
            .I(N__28364));
    Span4Mux_v I__6605 (
            .O(N__28383),
            .I(N__28364));
    Span4Mux_v I__6604 (
            .O(N__28378),
            .I(N__28361));
    LocalMux I__6603 (
            .O(N__28375),
            .I(N__28358));
    Span12Mux_h I__6602 (
            .O(N__28372),
            .I(N__28355));
    Sp12to4 I__6601 (
            .O(N__28369),
            .I(N__28350));
    Sp12to4 I__6600 (
            .O(N__28364),
            .I(N__28350));
    Span4Mux_v I__6599 (
            .O(N__28361),
            .I(N__28347));
    Span4Mux_h I__6598 (
            .O(N__28358),
            .I(N__28344));
    Span12Mux_v I__6597 (
            .O(N__28355),
            .I(N__28339));
    Span12Mux_h I__6596 (
            .O(N__28350),
            .I(N__28339));
    Span4Mux_v I__6595 (
            .O(N__28347),
            .I(N__28336));
    Span4Mux_v I__6594 (
            .O(N__28344),
            .I(N__28333));
    Odrv12 I__6593 (
            .O(N__28339),
            .I(port_data_c_0));
    Odrv4 I__6592 (
            .O(N__28336),
            .I(port_data_c_0));
    Odrv4 I__6591 (
            .O(N__28333),
            .I(port_data_c_0));
    InMux I__6590 (
            .O(N__28326),
            .I(N__28321));
    InMux I__6589 (
            .O(N__28325),
            .I(N__28317));
    InMux I__6588 (
            .O(N__28324),
            .I(N__28314));
    LocalMux I__6587 (
            .O(N__28321),
            .I(N__28311));
    CascadeMux I__6586 (
            .O(N__28320),
            .I(N__28308));
    LocalMux I__6585 (
            .O(N__28317),
            .I(N__28303));
    LocalMux I__6584 (
            .O(N__28314),
            .I(N__28303));
    Span4Mux_v I__6583 (
            .O(N__28311),
            .I(N__28298));
    InMux I__6582 (
            .O(N__28308),
            .I(N__28295));
    Span4Mux_h I__6581 (
            .O(N__28303),
            .I(N__28291));
    InMux I__6580 (
            .O(N__28302),
            .I(N__28286));
    InMux I__6579 (
            .O(N__28301),
            .I(N__28286));
    Span4Mux_h I__6578 (
            .O(N__28298),
            .I(N__28282));
    LocalMux I__6577 (
            .O(N__28295),
            .I(N__28279));
    CascadeMux I__6576 (
            .O(N__28294),
            .I(N__28276));
    Span4Mux_h I__6575 (
            .O(N__28291),
            .I(N__28270));
    LocalMux I__6574 (
            .O(N__28286),
            .I(N__28270));
    InMux I__6573 (
            .O(N__28285),
            .I(N__28267));
    Span4Mux_h I__6572 (
            .O(N__28282),
            .I(N__28263));
    Span4Mux_h I__6571 (
            .O(N__28279),
            .I(N__28260));
    InMux I__6570 (
            .O(N__28276),
            .I(N__28257));
    CascadeMux I__6569 (
            .O(N__28275),
            .I(N__28254));
    Span4Mux_h I__6568 (
            .O(N__28270),
            .I(N__28249));
    LocalMux I__6567 (
            .O(N__28267),
            .I(N__28249));
    InMux I__6566 (
            .O(N__28266),
            .I(N__28246));
    Span4Mux_h I__6565 (
            .O(N__28263),
            .I(N__28238));
    Span4Mux_v I__6564 (
            .O(N__28260),
            .I(N__28238));
    LocalMux I__6563 (
            .O(N__28257),
            .I(N__28238));
    InMux I__6562 (
            .O(N__28254),
            .I(N__28235));
    Span4Mux_h I__6561 (
            .O(N__28249),
            .I(N__28232));
    LocalMux I__6560 (
            .O(N__28246),
            .I(N__28229));
    InMux I__6559 (
            .O(N__28245),
            .I(N__28226));
    Span4Mux_v I__6558 (
            .O(N__28238),
            .I(N__28223));
    LocalMux I__6557 (
            .O(N__28235),
            .I(N__28220));
    Sp12to4 I__6556 (
            .O(N__28232),
            .I(N__28217));
    Span12Mux_v I__6555 (
            .O(N__28229),
            .I(N__28212));
    LocalMux I__6554 (
            .O(N__28226),
            .I(N__28212));
    Span4Mux_v I__6553 (
            .O(N__28223),
            .I(N__28209));
    Span4Mux_v I__6552 (
            .O(N__28220),
            .I(N__28206));
    Span12Mux_v I__6551 (
            .O(N__28217),
            .I(N__28203));
    Span12Mux_h I__6550 (
            .O(N__28212),
            .I(N__28196));
    Sp12to4 I__6549 (
            .O(N__28209),
            .I(N__28196));
    Sp12to4 I__6548 (
            .O(N__28206),
            .I(N__28196));
    Odrv12 I__6547 (
            .O(N__28203),
            .I(port_data_c_4));
    Odrv12 I__6546 (
            .O(N__28196),
            .I(port_data_c_4));
    InMux I__6545 (
            .O(N__28191),
            .I(N__28186));
    InMux I__6544 (
            .O(N__28190),
            .I(N__28183));
    InMux I__6543 (
            .O(N__28189),
            .I(N__28180));
    LocalMux I__6542 (
            .O(N__28186),
            .I(N__28176));
    LocalMux I__6541 (
            .O(N__28183),
            .I(N__28171));
    LocalMux I__6540 (
            .O(N__28180),
            .I(N__28171));
    InMux I__6539 (
            .O(N__28179),
            .I(N__28168));
    Span4Mux_v I__6538 (
            .O(N__28176),
            .I(N__28163));
    Span4Mux_v I__6537 (
            .O(N__28171),
            .I(N__28158));
    LocalMux I__6536 (
            .O(N__28168),
            .I(N__28158));
    CascadeMux I__6535 (
            .O(N__28167),
            .I(N__28155));
    CascadeMux I__6534 (
            .O(N__28166),
            .I(N__28152));
    Span4Mux_h I__6533 (
            .O(N__28163),
            .I(N__28149));
    Span4Mux_h I__6532 (
            .O(N__28158),
            .I(N__28145));
    InMux I__6531 (
            .O(N__28155),
            .I(N__28142));
    InMux I__6530 (
            .O(N__28152),
            .I(N__28139));
    Span4Mux_v I__6529 (
            .O(N__28149),
            .I(N__28136));
    InMux I__6528 (
            .O(N__28148),
            .I(N__28133));
    Span4Mux_h I__6527 (
            .O(N__28145),
            .I(N__28128));
    LocalMux I__6526 (
            .O(N__28142),
            .I(N__28128));
    LocalMux I__6525 (
            .O(N__28139),
            .I(N__28124));
    Span4Mux_v I__6524 (
            .O(N__28136),
            .I(N__28119));
    LocalMux I__6523 (
            .O(N__28133),
            .I(N__28119));
    Span4Mux_v I__6522 (
            .O(N__28128),
            .I(N__28116));
    InMux I__6521 (
            .O(N__28127),
            .I(N__28113));
    Span4Mux_v I__6520 (
            .O(N__28124),
            .I(N__28110));
    Span4Mux_v I__6519 (
            .O(N__28119),
            .I(N__28105));
    Span4Mux_h I__6518 (
            .O(N__28116),
            .I(N__28100));
    LocalMux I__6517 (
            .O(N__28113),
            .I(N__28100));
    Span4Mux_h I__6516 (
            .O(N__28110),
            .I(N__28097));
    InMux I__6515 (
            .O(N__28109),
            .I(N__28093));
    CascadeMux I__6514 (
            .O(N__28108),
            .I(N__28090));
    Span4Mux_v I__6513 (
            .O(N__28105),
            .I(N__28087));
    Span4Mux_v I__6512 (
            .O(N__28100),
            .I(N__28084));
    Sp12to4 I__6511 (
            .O(N__28097),
            .I(N__28081));
    InMux I__6510 (
            .O(N__28096),
            .I(N__28078));
    LocalMux I__6509 (
            .O(N__28093),
            .I(N__28075));
    InMux I__6508 (
            .O(N__28090),
            .I(N__28072));
    Sp12to4 I__6507 (
            .O(N__28087),
            .I(N__28069));
    Span4Mux_v I__6506 (
            .O(N__28084),
            .I(N__28066));
    Span12Mux_s8_h I__6505 (
            .O(N__28081),
            .I(N__28057));
    LocalMux I__6504 (
            .O(N__28078),
            .I(N__28057));
    Sp12to4 I__6503 (
            .O(N__28075),
            .I(N__28057));
    LocalMux I__6502 (
            .O(N__28072),
            .I(N__28057));
    Span12Mux_h I__6501 (
            .O(N__28069),
            .I(N__28050));
    Sp12to4 I__6500 (
            .O(N__28066),
            .I(N__28050));
    Span12Mux_v I__6499 (
            .O(N__28057),
            .I(N__28050));
    Odrv12 I__6498 (
            .O(N__28050),
            .I(port_data_c_6));
    CascadeMux I__6497 (
            .O(N__28047),
            .I(\this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3Z0Z_0_cascade_ ));
    CascadeMux I__6496 (
            .O(N__28044),
            .I(N__28041));
    InMux I__6495 (
            .O(N__28041),
            .I(N__28037));
    CascadeMux I__6494 (
            .O(N__28040),
            .I(N__28033));
    LocalMux I__6493 (
            .O(N__28037),
            .I(N__28029));
    InMux I__6492 (
            .O(N__28036),
            .I(N__28026));
    InMux I__6491 (
            .O(N__28033),
            .I(N__28023));
    InMux I__6490 (
            .O(N__28032),
            .I(N__28020));
    Span4Mux_v I__6489 (
            .O(N__28029),
            .I(N__28015));
    LocalMux I__6488 (
            .O(N__28026),
            .I(N__28015));
    LocalMux I__6487 (
            .O(N__28023),
            .I(N__28011));
    LocalMux I__6486 (
            .O(N__28020),
            .I(N__28008));
    Span4Mux_v I__6485 (
            .O(N__28015),
            .I(N__28005));
    InMux I__6484 (
            .O(N__28014),
            .I(N__28002));
    Span4Mux_v I__6483 (
            .O(N__28011),
            .I(N__27999));
    Span4Mux_h I__6482 (
            .O(N__28008),
            .I(N__27996));
    Sp12to4 I__6481 (
            .O(N__28005),
            .I(N__27991));
    LocalMux I__6480 (
            .O(N__28002),
            .I(N__27991));
    Odrv4 I__6479 (
            .O(N__27999),
            .I(\this_start_data_delay.N_902_0 ));
    Odrv4 I__6478 (
            .O(N__27996),
            .I(\this_start_data_delay.N_902_0 ));
    Odrv12 I__6477 (
            .O(N__27991),
            .I(\this_start_data_delay.N_902_0 ));
    InMux I__6476 (
            .O(N__27984),
            .I(N__27981));
    LocalMux I__6475 (
            .O(N__27981),
            .I(N__27975));
    InMux I__6474 (
            .O(N__27980),
            .I(N__27972));
    InMux I__6473 (
            .O(N__27979),
            .I(N__27969));
    InMux I__6472 (
            .O(N__27978),
            .I(N__27966));
    Span4Mux_h I__6471 (
            .O(N__27975),
            .I(N__27963));
    LocalMux I__6470 (
            .O(N__27972),
            .I(N__27960));
    LocalMux I__6469 (
            .O(N__27969),
            .I(N__27957));
    LocalMux I__6468 (
            .O(N__27966),
            .I(N__27954));
    Odrv4 I__6467 (
            .O(N__27963),
            .I(\this_start_data_delay.N_821_0 ));
    Odrv4 I__6466 (
            .O(N__27960),
            .I(\this_start_data_delay.N_821_0 ));
    Odrv4 I__6465 (
            .O(N__27957),
            .I(\this_start_data_delay.N_821_0 ));
    Odrv4 I__6464 (
            .O(N__27954),
            .I(\this_start_data_delay.N_821_0 ));
    InMux I__6463 (
            .O(N__27945),
            .I(N__27942));
    LocalMux I__6462 (
            .O(N__27942),
            .I(N__27938));
    CascadeMux I__6461 (
            .O(N__27941),
            .I(N__27934));
    Span4Mux_h I__6460 (
            .O(N__27938),
            .I(N__27930));
    InMux I__6459 (
            .O(N__27937),
            .I(N__27926));
    InMux I__6458 (
            .O(N__27934),
            .I(N__27923));
    InMux I__6457 (
            .O(N__27933),
            .I(N__27920));
    Span4Mux_h I__6456 (
            .O(N__27930),
            .I(N__27917));
    CascadeMux I__6455 (
            .O(N__27929),
            .I(N__27913));
    LocalMux I__6454 (
            .O(N__27926),
            .I(N__27908));
    LocalMux I__6453 (
            .O(N__27923),
            .I(N__27902));
    LocalMux I__6452 (
            .O(N__27920),
            .I(N__27902));
    Span4Mux_h I__6451 (
            .O(N__27917),
            .I(N__27899));
    InMux I__6450 (
            .O(N__27916),
            .I(N__27894));
    InMux I__6449 (
            .O(N__27913),
            .I(N__27894));
    InMux I__6448 (
            .O(N__27912),
            .I(N__27891));
    InMux I__6447 (
            .O(N__27911),
            .I(N__27888));
    Span4Mux_h I__6446 (
            .O(N__27908),
            .I(N__27885));
    InMux I__6445 (
            .O(N__27907),
            .I(N__27882));
    Span4Mux_v I__6444 (
            .O(N__27902),
            .I(N__27879));
    Span4Mux_h I__6443 (
            .O(N__27899),
            .I(N__27874));
    LocalMux I__6442 (
            .O(N__27894),
            .I(N__27874));
    LocalMux I__6441 (
            .O(N__27891),
            .I(N__27865));
    LocalMux I__6440 (
            .O(N__27888),
            .I(N__27865));
    Sp12to4 I__6439 (
            .O(N__27885),
            .I(N__27865));
    LocalMux I__6438 (
            .O(N__27882),
            .I(N__27865));
    Sp12to4 I__6437 (
            .O(N__27879),
            .I(N__27862));
    Span4Mux_v I__6436 (
            .O(N__27874),
            .I(N__27859));
    Span12Mux_v I__6435 (
            .O(N__27865),
            .I(N__27856));
    Span12Mux_h I__6434 (
            .O(N__27862),
            .I(N__27853));
    Span4Mux_h I__6433 (
            .O(N__27859),
            .I(N__27850));
    Span12Mux_h I__6432 (
            .O(N__27856),
            .I(N__27847));
    Span12Mux_v I__6431 (
            .O(N__27853),
            .I(N__27844));
    IoSpan4Mux I__6430 (
            .O(N__27850),
            .I(N__27841));
    Odrv12 I__6429 (
            .O(N__27847),
            .I(port_data_c_7));
    Odrv12 I__6428 (
            .O(N__27844),
            .I(port_data_c_7));
    Odrv4 I__6427 (
            .O(N__27841),
            .I(port_data_c_7));
    InMux I__6426 (
            .O(N__27834),
            .I(N__27831));
    LocalMux I__6425 (
            .O(N__27831),
            .I(N__27827));
    InMux I__6424 (
            .O(N__27830),
            .I(N__27824));
    Span4Mux_v I__6423 (
            .O(N__27827),
            .I(N__27817));
    LocalMux I__6422 (
            .O(N__27824),
            .I(N__27817));
    InMux I__6421 (
            .O(N__27823),
            .I(N__27814));
    InMux I__6420 (
            .O(N__27822),
            .I(N__27811));
    Odrv4 I__6419 (
            .O(N__27817),
            .I(\this_start_data_delay.N_123 ));
    LocalMux I__6418 (
            .O(N__27814),
            .I(\this_start_data_delay.N_123 ));
    LocalMux I__6417 (
            .O(N__27811),
            .I(\this_start_data_delay.N_123 ));
    InMux I__6416 (
            .O(N__27804),
            .I(N__27800));
    InMux I__6415 (
            .O(N__27803),
            .I(N__27796));
    LocalMux I__6414 (
            .O(N__27800),
            .I(N__27792));
    InMux I__6413 (
            .O(N__27799),
            .I(N__27789));
    LocalMux I__6412 (
            .O(N__27796),
            .I(N__27785));
    InMux I__6411 (
            .O(N__27795),
            .I(N__27782));
    Span4Mux_v I__6410 (
            .O(N__27792),
            .I(N__27776));
    LocalMux I__6409 (
            .O(N__27789),
            .I(N__27776));
    InMux I__6408 (
            .O(N__27788),
            .I(N__27773));
    Span4Mux_v I__6407 (
            .O(N__27785),
            .I(N__27767));
    LocalMux I__6406 (
            .O(N__27782),
            .I(N__27767));
    InMux I__6405 (
            .O(N__27781),
            .I(N__27764));
    Span4Mux_v I__6404 (
            .O(N__27776),
            .I(N__27758));
    LocalMux I__6403 (
            .O(N__27773),
            .I(N__27758));
    InMux I__6402 (
            .O(N__27772),
            .I(N__27755));
    Span4Mux_v I__6401 (
            .O(N__27767),
            .I(N__27750));
    LocalMux I__6400 (
            .O(N__27764),
            .I(N__27750));
    InMux I__6399 (
            .O(N__27763),
            .I(N__27747));
    Span4Mux_v I__6398 (
            .O(N__27758),
            .I(N__27742));
    LocalMux I__6397 (
            .O(N__27755),
            .I(N__27742));
    Span4Mux_v I__6396 (
            .O(N__27750),
            .I(N__27737));
    LocalMux I__6395 (
            .O(N__27747),
            .I(N__27737));
    Odrv4 I__6394 (
            .O(N__27742),
            .I(N_41_0));
    Odrv4 I__6393 (
            .O(N__27737),
            .I(N_41_0));
    InMux I__6392 (
            .O(N__27732),
            .I(N__27729));
    LocalMux I__6391 (
            .O(N__27729),
            .I(\this_sprites_ram.mem_out_bus4_0 ));
    InMux I__6390 (
            .O(N__27726),
            .I(N__27723));
    LocalMux I__6389 (
            .O(N__27723),
            .I(N__27720));
    Sp12to4 I__6388 (
            .O(N__27720),
            .I(N__27717));
    Span12Mux_v I__6387 (
            .O(N__27717),
            .I(N__27714));
    Odrv12 I__6386 (
            .O(N__27714),
            .I(\this_sprites_ram.mem_out_bus0_0 ));
    InMux I__6385 (
            .O(N__27711),
            .I(N__27708));
    LocalMux I__6384 (
            .O(N__27708),
            .I(\this_sprites_ram.mem_out_bus4_3 ));
    InMux I__6383 (
            .O(N__27705),
            .I(N__27702));
    LocalMux I__6382 (
            .O(N__27702),
            .I(N__27699));
    Span4Mux_v I__6381 (
            .O(N__27699),
            .I(N__27696));
    Span4Mux_v I__6380 (
            .O(N__27696),
            .I(N__27693));
    Span4Mux_v I__6379 (
            .O(N__27693),
            .I(N__27690));
    Odrv4 I__6378 (
            .O(N__27690),
            .I(\this_sprites_ram.mem_out_bus0_3 ));
    InMux I__6377 (
            .O(N__27687),
            .I(N__27684));
    LocalMux I__6376 (
            .O(N__27684),
            .I(N__27681));
    Sp12to4 I__6375 (
            .O(N__27681),
            .I(N__27678));
    Odrv12 I__6374 (
            .O(N__27678),
            .I(\this_sprites_ram.mem_out_bus6_3 ));
    InMux I__6373 (
            .O(N__27675),
            .I(N__27672));
    LocalMux I__6372 (
            .O(N__27672),
            .I(N__27669));
    Span4Mux_v I__6371 (
            .O(N__27669),
            .I(N__27666));
    Odrv4 I__6370 (
            .O(N__27666),
            .I(\this_sprites_ram.mem_out_bus2_3 ));
    InMux I__6369 (
            .O(N__27663),
            .I(N__27660));
    LocalMux I__6368 (
            .O(N__27660),
            .I(N__27654));
    CascadeMux I__6367 (
            .O(N__27659),
            .I(N__27650));
    CascadeMux I__6366 (
            .O(N__27658),
            .I(N__27647));
    InMux I__6365 (
            .O(N__27657),
            .I(N__27642));
    Span4Mux_h I__6364 (
            .O(N__27654),
            .I(N__27639));
    InMux I__6363 (
            .O(N__27653),
            .I(N__27634));
    InMux I__6362 (
            .O(N__27650),
            .I(N__27634));
    InMux I__6361 (
            .O(N__27647),
            .I(N__27631));
    InMux I__6360 (
            .O(N__27646),
            .I(N__27628));
    InMux I__6359 (
            .O(N__27645),
            .I(N__27625));
    LocalMux I__6358 (
            .O(N__27642),
            .I(\this_start_data_delay.N_992 ));
    Odrv4 I__6357 (
            .O(N__27639),
            .I(\this_start_data_delay.N_992 ));
    LocalMux I__6356 (
            .O(N__27634),
            .I(\this_start_data_delay.N_992 ));
    LocalMux I__6355 (
            .O(N__27631),
            .I(\this_start_data_delay.N_992 ));
    LocalMux I__6354 (
            .O(N__27628),
            .I(\this_start_data_delay.N_992 ));
    LocalMux I__6353 (
            .O(N__27625),
            .I(\this_start_data_delay.N_992 ));
    InMux I__6352 (
            .O(N__27612),
            .I(N__27608));
    InMux I__6351 (
            .O(N__27611),
            .I(N__27604));
    LocalMux I__6350 (
            .O(N__27608),
            .I(N__27598));
    InMux I__6349 (
            .O(N__27607),
            .I(N__27595));
    LocalMux I__6348 (
            .O(N__27604),
            .I(N__27592));
    InMux I__6347 (
            .O(N__27603),
            .I(N__27589));
    InMux I__6346 (
            .O(N__27602),
            .I(N__27584));
    InMux I__6345 (
            .O(N__27601),
            .I(N__27584));
    Odrv4 I__6344 (
            .O(N__27598),
            .I(\this_start_data_delay.N_110 ));
    LocalMux I__6343 (
            .O(N__27595),
            .I(\this_start_data_delay.N_110 ));
    Odrv4 I__6342 (
            .O(N__27592),
            .I(\this_start_data_delay.N_110 ));
    LocalMux I__6341 (
            .O(N__27589),
            .I(\this_start_data_delay.N_110 ));
    LocalMux I__6340 (
            .O(N__27584),
            .I(\this_start_data_delay.N_110 ));
    InMux I__6339 (
            .O(N__27573),
            .I(N__27570));
    LocalMux I__6338 (
            .O(N__27570),
            .I(un1_M_this_sprites_address_q_cry_7_THRU_CO));
    CascadeMux I__6337 (
            .O(N__27567),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_8_cascade_ ));
    InMux I__6336 (
            .O(N__27564),
            .I(N__27554));
    InMux I__6335 (
            .O(N__27563),
            .I(N__27547));
    InMux I__6334 (
            .O(N__27562),
            .I(N__27547));
    InMux I__6333 (
            .O(N__27561),
            .I(N__27547));
    InMux I__6332 (
            .O(N__27560),
            .I(N__27544));
    InMux I__6331 (
            .O(N__27559),
            .I(N__27537));
    InMux I__6330 (
            .O(N__27558),
            .I(N__27537));
    InMux I__6329 (
            .O(N__27557),
            .I(N__27534));
    LocalMux I__6328 (
            .O(N__27554),
            .I(N__27527));
    LocalMux I__6327 (
            .O(N__27547),
            .I(N__27527));
    LocalMux I__6326 (
            .O(N__27544),
            .I(N__27524));
    InMux I__6325 (
            .O(N__27543),
            .I(N__27519));
    InMux I__6324 (
            .O(N__27542),
            .I(N__27519));
    LocalMux I__6323 (
            .O(N__27537),
            .I(N__27512));
    LocalMux I__6322 (
            .O(N__27534),
            .I(N__27512));
    InMux I__6321 (
            .O(N__27533),
            .I(N__27507));
    InMux I__6320 (
            .O(N__27532),
            .I(N__27507));
    Span4Mux_v I__6319 (
            .O(N__27527),
            .I(N__27500));
    Span4Mux_h I__6318 (
            .O(N__27524),
            .I(N__27500));
    LocalMux I__6317 (
            .O(N__27519),
            .I(N__27500));
    InMux I__6316 (
            .O(N__27518),
            .I(N__27497));
    InMux I__6315 (
            .O(N__27517),
            .I(N__27494));
    Odrv4 I__6314 (
            .O(N__27512),
            .I(\this_start_data_delay.N_990 ));
    LocalMux I__6313 (
            .O(N__27507),
            .I(\this_start_data_delay.N_990 ));
    Odrv4 I__6312 (
            .O(N__27500),
            .I(\this_start_data_delay.N_990 ));
    LocalMux I__6311 (
            .O(N__27497),
            .I(\this_start_data_delay.N_990 ));
    LocalMux I__6310 (
            .O(N__27494),
            .I(\this_start_data_delay.N_990 ));
    CascadeMux I__6309 (
            .O(N__27483),
            .I(N__27480));
    CascadeBuf I__6308 (
            .O(N__27480),
            .I(N__27477));
    CascadeMux I__6307 (
            .O(N__27477),
            .I(N__27474));
    CascadeBuf I__6306 (
            .O(N__27474),
            .I(N__27471));
    CascadeMux I__6305 (
            .O(N__27471),
            .I(N__27468));
    CascadeBuf I__6304 (
            .O(N__27468),
            .I(N__27465));
    CascadeMux I__6303 (
            .O(N__27465),
            .I(N__27462));
    CascadeBuf I__6302 (
            .O(N__27462),
            .I(N__27459));
    CascadeMux I__6301 (
            .O(N__27459),
            .I(N__27456));
    CascadeBuf I__6300 (
            .O(N__27456),
            .I(N__27453));
    CascadeMux I__6299 (
            .O(N__27453),
            .I(N__27450));
    CascadeBuf I__6298 (
            .O(N__27450),
            .I(N__27447));
    CascadeMux I__6297 (
            .O(N__27447),
            .I(N__27444));
    CascadeBuf I__6296 (
            .O(N__27444),
            .I(N__27441));
    CascadeMux I__6295 (
            .O(N__27441),
            .I(N__27438));
    CascadeBuf I__6294 (
            .O(N__27438),
            .I(N__27435));
    CascadeMux I__6293 (
            .O(N__27435),
            .I(N__27432));
    CascadeBuf I__6292 (
            .O(N__27432),
            .I(N__27429));
    CascadeMux I__6291 (
            .O(N__27429),
            .I(N__27426));
    CascadeBuf I__6290 (
            .O(N__27426),
            .I(N__27423));
    CascadeMux I__6289 (
            .O(N__27423),
            .I(N__27420));
    CascadeBuf I__6288 (
            .O(N__27420),
            .I(N__27417));
    CascadeMux I__6287 (
            .O(N__27417),
            .I(N__27414));
    CascadeBuf I__6286 (
            .O(N__27414),
            .I(N__27411));
    CascadeMux I__6285 (
            .O(N__27411),
            .I(N__27408));
    CascadeBuf I__6284 (
            .O(N__27408),
            .I(N__27405));
    CascadeMux I__6283 (
            .O(N__27405),
            .I(N__27402));
    CascadeBuf I__6282 (
            .O(N__27402),
            .I(N__27399));
    CascadeMux I__6281 (
            .O(N__27399),
            .I(N__27396));
    CascadeBuf I__6280 (
            .O(N__27396),
            .I(N__27393));
    CascadeMux I__6279 (
            .O(N__27393),
            .I(N__27390));
    InMux I__6278 (
            .O(N__27390),
            .I(N__27387));
    LocalMux I__6277 (
            .O(N__27387),
            .I(N__27384));
    Span4Mux_s3_v I__6276 (
            .O(N__27384),
            .I(N__27381));
    Span4Mux_v I__6275 (
            .O(N__27381),
            .I(N__27375));
    InMux I__6274 (
            .O(N__27380),
            .I(N__27372));
    InMux I__6273 (
            .O(N__27379),
            .I(N__27369));
    InMux I__6272 (
            .O(N__27378),
            .I(N__27366));
    Span4Mux_v I__6271 (
            .O(N__27375),
            .I(N__27363));
    LocalMux I__6270 (
            .O(N__27372),
            .I(M_this_sprites_address_qZ0Z_8));
    LocalMux I__6269 (
            .O(N__27369),
            .I(M_this_sprites_address_qZ0Z_8));
    LocalMux I__6268 (
            .O(N__27366),
            .I(M_this_sprites_address_qZ0Z_8));
    Odrv4 I__6267 (
            .O(N__27363),
            .I(M_this_sprites_address_qZ0Z_8));
    InMux I__6266 (
            .O(N__27354),
            .I(N__27351));
    LocalMux I__6265 (
            .O(N__27351),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ));
    CEMux I__6264 (
            .O(N__27348),
            .I(N__27344));
    CEMux I__6263 (
            .O(N__27347),
            .I(N__27341));
    LocalMux I__6262 (
            .O(N__27344),
            .I(N__27336));
    LocalMux I__6261 (
            .O(N__27341),
            .I(N__27336));
    Span4Mux_v I__6260 (
            .O(N__27336),
            .I(N__27333));
    Span4Mux_h I__6259 (
            .O(N__27333),
            .I(N__27330));
    Odrv4 I__6258 (
            .O(N__27330),
            .I(\this_sprites_ram.mem_WE_10 ));
    CEMux I__6257 (
            .O(N__27327),
            .I(N__27323));
    CEMux I__6256 (
            .O(N__27326),
            .I(N__27320));
    LocalMux I__6255 (
            .O(N__27323),
            .I(N__27317));
    LocalMux I__6254 (
            .O(N__27320),
            .I(N__27314));
    Span4Mux_h I__6253 (
            .O(N__27317),
            .I(N__27311));
    Span4Mux_h I__6252 (
            .O(N__27314),
            .I(N__27308));
    Odrv4 I__6251 (
            .O(N__27311),
            .I(\this_sprites_ram.mem_WE_8 ));
    Odrv4 I__6250 (
            .O(N__27308),
            .I(\this_sprites_ram.mem_WE_8 ));
    CEMux I__6249 (
            .O(N__27303),
            .I(N__27300));
    LocalMux I__6248 (
            .O(N__27300),
            .I(N__27296));
    CEMux I__6247 (
            .O(N__27299),
            .I(N__27293));
    Span4Mux_v I__6246 (
            .O(N__27296),
            .I(N__27288));
    LocalMux I__6245 (
            .O(N__27293),
            .I(N__27288));
    Span4Mux_v I__6244 (
            .O(N__27288),
            .I(N__27285));
    Odrv4 I__6243 (
            .O(N__27285),
            .I(\this_sprites_ram.mem_WE_12 ));
    CEMux I__6242 (
            .O(N__27282),
            .I(N__27279));
    LocalMux I__6241 (
            .O(N__27279),
            .I(N__27275));
    CEMux I__6240 (
            .O(N__27278),
            .I(N__27272));
    Span4Mux_s1_v I__6239 (
            .O(N__27275),
            .I(N__27267));
    LocalMux I__6238 (
            .O(N__27272),
            .I(N__27267));
    Span4Mux_v I__6237 (
            .O(N__27267),
            .I(N__27264));
    Span4Mux_v I__6236 (
            .O(N__27264),
            .I(N__27261));
    Odrv4 I__6235 (
            .O(N__27261),
            .I(\this_sprites_ram.mem_WE_14 ));
    InMux I__6234 (
            .O(N__27258),
            .I(N__27255));
    LocalMux I__6233 (
            .O(N__27255),
            .I(N__27251));
    InMux I__6232 (
            .O(N__27254),
            .I(N__27248));
    Span4Mux_v I__6231 (
            .O(N__27251),
            .I(N__27241));
    LocalMux I__6230 (
            .O(N__27248),
            .I(N__27241));
    InMux I__6229 (
            .O(N__27247),
            .I(N__27238));
    InMux I__6228 (
            .O(N__27246),
            .I(N__27234));
    Span4Mux_v I__6227 (
            .O(N__27241),
            .I(N__27228));
    LocalMux I__6226 (
            .O(N__27238),
            .I(N__27228));
    InMux I__6225 (
            .O(N__27237),
            .I(N__27225));
    LocalMux I__6224 (
            .O(N__27234),
            .I(N__27222));
    InMux I__6223 (
            .O(N__27233),
            .I(N__27219));
    Span4Mux_v I__6222 (
            .O(N__27228),
            .I(N__27213));
    LocalMux I__6221 (
            .O(N__27225),
            .I(N__27213));
    Span4Mux_v I__6220 (
            .O(N__27222),
            .I(N__27208));
    LocalMux I__6219 (
            .O(N__27219),
            .I(N__27208));
    InMux I__6218 (
            .O(N__27218),
            .I(N__27205));
    Span4Mux_v I__6217 (
            .O(N__27213),
            .I(N__27201));
    Span4Mux_v I__6216 (
            .O(N__27208),
            .I(N__27196));
    LocalMux I__6215 (
            .O(N__27205),
            .I(N__27196));
    InMux I__6214 (
            .O(N__27204),
            .I(N__27193));
    Odrv4 I__6213 (
            .O(N__27201),
            .I(N_811_0));
    Odrv4 I__6212 (
            .O(N__27196),
            .I(N_811_0));
    LocalMux I__6211 (
            .O(N__27193),
            .I(N_811_0));
    InMux I__6210 (
            .O(N__27186),
            .I(N__27183));
    LocalMux I__6209 (
            .O(N__27183),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_5 ));
    InMux I__6208 (
            .O(N__27180),
            .I(N__27177));
    LocalMux I__6207 (
            .O(N__27177),
            .I(un1_M_this_sprites_address_q_cry_4_THRU_CO));
    CascadeMux I__6206 (
            .O(N__27174),
            .I(N__27171));
    CascadeBuf I__6205 (
            .O(N__27171),
            .I(N__27168));
    CascadeMux I__6204 (
            .O(N__27168),
            .I(N__27165));
    CascadeBuf I__6203 (
            .O(N__27165),
            .I(N__27162));
    CascadeMux I__6202 (
            .O(N__27162),
            .I(N__27159));
    CascadeBuf I__6201 (
            .O(N__27159),
            .I(N__27156));
    CascadeMux I__6200 (
            .O(N__27156),
            .I(N__27153));
    CascadeBuf I__6199 (
            .O(N__27153),
            .I(N__27150));
    CascadeMux I__6198 (
            .O(N__27150),
            .I(N__27147));
    CascadeBuf I__6197 (
            .O(N__27147),
            .I(N__27144));
    CascadeMux I__6196 (
            .O(N__27144),
            .I(N__27141));
    CascadeBuf I__6195 (
            .O(N__27141),
            .I(N__27138));
    CascadeMux I__6194 (
            .O(N__27138),
            .I(N__27135));
    CascadeBuf I__6193 (
            .O(N__27135),
            .I(N__27132));
    CascadeMux I__6192 (
            .O(N__27132),
            .I(N__27129));
    CascadeBuf I__6191 (
            .O(N__27129),
            .I(N__27126));
    CascadeMux I__6190 (
            .O(N__27126),
            .I(N__27123));
    CascadeBuf I__6189 (
            .O(N__27123),
            .I(N__27120));
    CascadeMux I__6188 (
            .O(N__27120),
            .I(N__27117));
    CascadeBuf I__6187 (
            .O(N__27117),
            .I(N__27114));
    CascadeMux I__6186 (
            .O(N__27114),
            .I(N__27111));
    CascadeBuf I__6185 (
            .O(N__27111),
            .I(N__27108));
    CascadeMux I__6184 (
            .O(N__27108),
            .I(N__27105));
    CascadeBuf I__6183 (
            .O(N__27105),
            .I(N__27102));
    CascadeMux I__6182 (
            .O(N__27102),
            .I(N__27099));
    CascadeBuf I__6181 (
            .O(N__27099),
            .I(N__27096));
    CascadeMux I__6180 (
            .O(N__27096),
            .I(N__27093));
    CascadeBuf I__6179 (
            .O(N__27093),
            .I(N__27090));
    CascadeMux I__6178 (
            .O(N__27090),
            .I(N__27087));
    CascadeBuf I__6177 (
            .O(N__27087),
            .I(N__27084));
    CascadeMux I__6176 (
            .O(N__27084),
            .I(N__27081));
    InMux I__6175 (
            .O(N__27081),
            .I(N__27078));
    LocalMux I__6174 (
            .O(N__27078),
            .I(N__27075));
    Span4Mux_h I__6173 (
            .O(N__27075),
            .I(N__27071));
    CascadeMux I__6172 (
            .O(N__27074),
            .I(N__27066));
    Sp12to4 I__6171 (
            .O(N__27071),
            .I(N__27063));
    InMux I__6170 (
            .O(N__27070),
            .I(N__27060));
    InMux I__6169 (
            .O(N__27069),
            .I(N__27057));
    InMux I__6168 (
            .O(N__27066),
            .I(N__27054));
    Span12Mux_s6_v I__6167 (
            .O(N__27063),
            .I(N__27051));
    LocalMux I__6166 (
            .O(N__27060),
            .I(M_this_sprites_address_qZ0Z_5));
    LocalMux I__6165 (
            .O(N__27057),
            .I(M_this_sprites_address_qZ0Z_5));
    LocalMux I__6164 (
            .O(N__27054),
            .I(M_this_sprites_address_qZ0Z_5));
    Odrv12 I__6163 (
            .O(N__27051),
            .I(M_this_sprites_address_qZ0Z_5));
    CEMux I__6162 (
            .O(N__27042),
            .I(N__27039));
    LocalMux I__6161 (
            .O(N__27039),
            .I(N__27036));
    Span4Mux_v I__6160 (
            .O(N__27036),
            .I(N__27032));
    CEMux I__6159 (
            .O(N__27035),
            .I(N__27029));
    Span4Mux_v I__6158 (
            .O(N__27032),
            .I(N__27024));
    LocalMux I__6157 (
            .O(N__27029),
            .I(N__27024));
    Span4Mux_h I__6156 (
            .O(N__27024),
            .I(N__27021));
    Odrv4 I__6155 (
            .O(N__27021),
            .I(\this_sprites_ram.mem_WE_6 ));
    InMux I__6154 (
            .O(N__27018),
            .I(N__27015));
    LocalMux I__6153 (
            .O(N__27015),
            .I(N__27012));
    Span4Mux_v I__6152 (
            .O(N__27012),
            .I(N__27009));
    Odrv4 I__6151 (
            .O(N__27009),
            .I(\this_sprites_ram.mem_out_bus5_0 ));
    InMux I__6150 (
            .O(N__27006),
            .I(N__27003));
    LocalMux I__6149 (
            .O(N__27003),
            .I(N__27000));
    Span4Mux_v I__6148 (
            .O(N__27000),
            .I(N__26997));
    Span4Mux_v I__6147 (
            .O(N__26997),
            .I(N__26994));
    Odrv4 I__6146 (
            .O(N__26994),
            .I(\this_sprites_ram.mem_out_bus1_0 ));
    InMux I__6145 (
            .O(N__26991),
            .I(N__26988));
    LocalMux I__6144 (
            .O(N__26988),
            .I(N__26985));
    Span12Mux_h I__6143 (
            .O(N__26985),
            .I(N__26982));
    Odrv12 I__6142 (
            .O(N__26982),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ));
    CascadeMux I__6141 (
            .O(N__26979),
            .I(N__26976));
    InMux I__6140 (
            .O(N__26976),
            .I(N__26968));
    InMux I__6139 (
            .O(N__26975),
            .I(N__26964));
    InMux I__6138 (
            .O(N__26974),
            .I(N__26958));
    InMux I__6137 (
            .O(N__26973),
            .I(N__26958));
    InMux I__6136 (
            .O(N__26972),
            .I(N__26955));
    InMux I__6135 (
            .O(N__26971),
            .I(N__26952));
    LocalMux I__6134 (
            .O(N__26968),
            .I(N__26949));
    InMux I__6133 (
            .O(N__26967),
            .I(N__26946));
    LocalMux I__6132 (
            .O(N__26964),
            .I(N__26943));
    InMux I__6131 (
            .O(N__26963),
            .I(N__26940));
    LocalMux I__6130 (
            .O(N__26958),
            .I(N__26937));
    LocalMux I__6129 (
            .O(N__26955),
            .I(N__26934));
    LocalMux I__6128 (
            .O(N__26952),
            .I(N__26931));
    Span4Mux_v I__6127 (
            .O(N__26949),
            .I(N__26928));
    LocalMux I__6126 (
            .O(N__26946),
            .I(N__26925));
    Span4Mux_h I__6125 (
            .O(N__26943),
            .I(N__26922));
    LocalMux I__6124 (
            .O(N__26940),
            .I(N__26917));
    Span4Mux_v I__6123 (
            .O(N__26937),
            .I(N__26917));
    Span4Mux_h I__6122 (
            .O(N__26934),
            .I(N__26912));
    Span4Mux_h I__6121 (
            .O(N__26931),
            .I(N__26912));
    Span4Mux_h I__6120 (
            .O(N__26928),
            .I(N__26907));
    Span4Mux_h I__6119 (
            .O(N__26925),
            .I(N__26907));
    Odrv4 I__6118 (
            .O(N__26922),
            .I(N_10_0));
    Odrv4 I__6117 (
            .O(N__26917),
            .I(N_10_0));
    Odrv4 I__6116 (
            .O(N__26912),
            .I(N_10_0));
    Odrv4 I__6115 (
            .O(N__26907),
            .I(N_10_0));
    InMux I__6114 (
            .O(N__26898),
            .I(N__26895));
    LocalMux I__6113 (
            .O(N__26895),
            .I(\this_start_data_delay.M_this_state_d62Z0Z_11 ));
    InMux I__6112 (
            .O(N__26892),
            .I(N__26889));
    LocalMux I__6111 (
            .O(N__26889),
            .I(\this_start_data_delay.M_this_state_d62Z0Z_10 ));
    CascadeMux I__6110 (
            .O(N__26886),
            .I(\this_start_data_delay.M_this_state_d62Z0Z_9_cascade_ ));
    InMux I__6109 (
            .O(N__26883),
            .I(N__26880));
    LocalMux I__6108 (
            .O(N__26880),
            .I(\this_start_data_delay.M_this_state_d62Z0Z_8 ));
    InMux I__6107 (
            .O(N__26877),
            .I(N__26872));
    InMux I__6106 (
            .O(N__26876),
            .I(N__26868));
    InMux I__6105 (
            .O(N__26875),
            .I(N__26864));
    LocalMux I__6104 (
            .O(N__26872),
            .I(N__26861));
    InMux I__6103 (
            .O(N__26871),
            .I(N__26858));
    LocalMux I__6102 (
            .O(N__26868),
            .I(N__26855));
    InMux I__6101 (
            .O(N__26867),
            .I(N__26852));
    LocalMux I__6100 (
            .O(N__26864),
            .I(N__26848));
    Span4Mux_h I__6099 (
            .O(N__26861),
            .I(N__26845));
    LocalMux I__6098 (
            .O(N__26858),
            .I(N__26840));
    Span4Mux_h I__6097 (
            .O(N__26855),
            .I(N__26840));
    LocalMux I__6096 (
            .O(N__26852),
            .I(N__26837));
    InMux I__6095 (
            .O(N__26851),
            .I(N__26834));
    Span4Mux_v I__6094 (
            .O(N__26848),
            .I(N__26831));
    Span4Mux_v I__6093 (
            .O(N__26845),
            .I(N__26828));
    Span4Mux_v I__6092 (
            .O(N__26840),
            .I(N__26825));
    Span4Mux_h I__6091 (
            .O(N__26837),
            .I(N__26820));
    LocalMux I__6090 (
            .O(N__26834),
            .I(N__26820));
    Odrv4 I__6089 (
            .O(N__26831),
            .I(\this_start_data_delay.M_this_state_dZ0Z62 ));
    Odrv4 I__6088 (
            .O(N__26828),
            .I(\this_start_data_delay.M_this_state_dZ0Z62 ));
    Odrv4 I__6087 (
            .O(N__26825),
            .I(\this_start_data_delay.M_this_state_dZ0Z62 ));
    Odrv4 I__6086 (
            .O(N__26820),
            .I(\this_start_data_delay.M_this_state_dZ0Z62 ));
    CascadeMux I__6085 (
            .O(N__26811),
            .I(N__26808));
    InMux I__6084 (
            .O(N__26808),
            .I(N__26805));
    LocalMux I__6083 (
            .O(N__26805),
            .I(M_this_data_count_q_3_10));
    InMux I__6082 (
            .O(N__26802),
            .I(N__26799));
    LocalMux I__6081 (
            .O(N__26799),
            .I(N__26796));
    Odrv12 I__6080 (
            .O(N__26796),
            .I(this_start_data_delay_M_this_external_address_q_3_i_0_15));
    InMux I__6079 (
            .O(N__26793),
            .I(N__26781));
    InMux I__6078 (
            .O(N__26792),
            .I(N__26781));
    InMux I__6077 (
            .O(N__26791),
            .I(N__26772));
    InMux I__6076 (
            .O(N__26790),
            .I(N__26772));
    InMux I__6075 (
            .O(N__26789),
            .I(N__26772));
    InMux I__6074 (
            .O(N__26788),
            .I(N__26772));
    InMux I__6073 (
            .O(N__26787),
            .I(N__26769));
    CascadeMux I__6072 (
            .O(N__26786),
            .I(N__26766));
    LocalMux I__6071 (
            .O(N__26781),
            .I(N__26762));
    LocalMux I__6070 (
            .O(N__26772),
            .I(N__26759));
    LocalMux I__6069 (
            .O(N__26769),
            .I(N__26756));
    InMux I__6068 (
            .O(N__26766),
            .I(N__26752));
    InMux I__6067 (
            .O(N__26765),
            .I(N__26749));
    Span4Mux_v I__6066 (
            .O(N__26762),
            .I(N__26746));
    Span4Mux_v I__6065 (
            .O(N__26759),
            .I(N__26743));
    Span4Mux_h I__6064 (
            .O(N__26756),
            .I(N__26740));
    InMux I__6063 (
            .O(N__26755),
            .I(N__26737));
    LocalMux I__6062 (
            .O(N__26752),
            .I(N__26734));
    LocalMux I__6061 (
            .O(N__26749),
            .I(N__26731));
    Span4Mux_h I__6060 (
            .O(N__26746),
            .I(N__26726));
    Span4Mux_h I__6059 (
            .O(N__26743),
            .I(N__26726));
    Sp12to4 I__6058 (
            .O(N__26740),
            .I(N__26721));
    LocalMux I__6057 (
            .O(N__26737),
            .I(N__26721));
    Span4Mux_v I__6056 (
            .O(N__26734),
            .I(N__26716));
    Span4Mux_v I__6055 (
            .O(N__26731),
            .I(N__26716));
    Sp12to4 I__6054 (
            .O(N__26726),
            .I(N__26713));
    Span12Mux_s10_v I__6053 (
            .O(N__26721),
            .I(N__26710));
    Odrv4 I__6052 (
            .O(N__26716),
            .I(N_116));
    Odrv12 I__6051 (
            .O(N__26713),
            .I(N_116));
    Odrv12 I__6050 (
            .O(N__26710),
            .I(N_116));
    InMux I__6049 (
            .O(N__26703),
            .I(N__26700));
    LocalMux I__6048 (
            .O(N__26700),
            .I(M_this_external_address_q_3_0_13));
    InMux I__6047 (
            .O(N__26697),
            .I(N__26694));
    LocalMux I__6046 (
            .O(N__26694),
            .I(N__26691));
    Span4Mux_s2_v I__6045 (
            .O(N__26691),
            .I(N__26688));
    Span4Mux_h I__6044 (
            .O(N__26688),
            .I(N__26685));
    Span4Mux_v I__6043 (
            .O(N__26685),
            .I(N__26682));
    Sp12to4 I__6042 (
            .O(N__26682),
            .I(N__26679));
    Odrv12 I__6041 (
            .O(N__26679),
            .I(M_this_map_ram_read_data_0));
    InMux I__6040 (
            .O(N__26676),
            .I(N__26673));
    LocalMux I__6039 (
            .O(N__26673),
            .I(N__26670));
    Span12Mux_h I__6038 (
            .O(N__26670),
            .I(N__26667));
    Span12Mux_v I__6037 (
            .O(N__26667),
            .I(N__26664));
    Odrv12 I__6036 (
            .O(N__26664),
            .I(\this_ppu.un3_sprites_addr_cry_5_c_RNI55GZ0Z8 ));
    CascadeMux I__6035 (
            .O(N__26661),
            .I(N__26658));
    CascadeBuf I__6034 (
            .O(N__26658),
            .I(N__26655));
    CascadeMux I__6033 (
            .O(N__26655),
            .I(N__26652));
    CascadeBuf I__6032 (
            .O(N__26652),
            .I(N__26649));
    CascadeMux I__6031 (
            .O(N__26649),
            .I(N__26646));
    CascadeBuf I__6030 (
            .O(N__26646),
            .I(N__26643));
    CascadeMux I__6029 (
            .O(N__26643),
            .I(N__26640));
    CascadeBuf I__6028 (
            .O(N__26640),
            .I(N__26637));
    CascadeMux I__6027 (
            .O(N__26637),
            .I(N__26634));
    CascadeBuf I__6026 (
            .O(N__26634),
            .I(N__26631));
    CascadeMux I__6025 (
            .O(N__26631),
            .I(N__26628));
    CascadeBuf I__6024 (
            .O(N__26628),
            .I(N__26625));
    CascadeMux I__6023 (
            .O(N__26625),
            .I(N__26622));
    CascadeBuf I__6022 (
            .O(N__26622),
            .I(N__26619));
    CascadeMux I__6021 (
            .O(N__26619),
            .I(N__26616));
    CascadeBuf I__6020 (
            .O(N__26616),
            .I(N__26613));
    CascadeMux I__6019 (
            .O(N__26613),
            .I(N__26610));
    CascadeBuf I__6018 (
            .O(N__26610),
            .I(N__26607));
    CascadeMux I__6017 (
            .O(N__26607),
            .I(N__26604));
    CascadeBuf I__6016 (
            .O(N__26604),
            .I(N__26601));
    CascadeMux I__6015 (
            .O(N__26601),
            .I(N__26598));
    CascadeBuf I__6014 (
            .O(N__26598),
            .I(N__26595));
    CascadeMux I__6013 (
            .O(N__26595),
            .I(N__26592));
    CascadeBuf I__6012 (
            .O(N__26592),
            .I(N__26589));
    CascadeMux I__6011 (
            .O(N__26589),
            .I(N__26586));
    CascadeBuf I__6010 (
            .O(N__26586),
            .I(N__26583));
    CascadeMux I__6009 (
            .O(N__26583),
            .I(N__26580));
    CascadeBuf I__6008 (
            .O(N__26580),
            .I(N__26577));
    CascadeMux I__6007 (
            .O(N__26577),
            .I(N__26574));
    CascadeBuf I__6006 (
            .O(N__26574),
            .I(N__26571));
    CascadeMux I__6005 (
            .O(N__26571),
            .I(N__26568));
    InMux I__6004 (
            .O(N__26568),
            .I(N__26565));
    LocalMux I__6003 (
            .O(N__26565),
            .I(N__26562));
    Odrv4 I__6002 (
            .O(N__26562),
            .I(M_this_ppu_sprites_addr_6));
    CascadeMux I__6001 (
            .O(N__26559),
            .I(N__26556));
    CascadeBuf I__6000 (
            .O(N__26556),
            .I(N__26553));
    CascadeMux I__5999 (
            .O(N__26553),
            .I(N__26550));
    CascadeBuf I__5998 (
            .O(N__26550),
            .I(N__26547));
    CascadeMux I__5997 (
            .O(N__26547),
            .I(N__26544));
    CascadeBuf I__5996 (
            .O(N__26544),
            .I(N__26541));
    CascadeMux I__5995 (
            .O(N__26541),
            .I(N__26538));
    CascadeBuf I__5994 (
            .O(N__26538),
            .I(N__26535));
    CascadeMux I__5993 (
            .O(N__26535),
            .I(N__26532));
    CascadeBuf I__5992 (
            .O(N__26532),
            .I(N__26529));
    CascadeMux I__5991 (
            .O(N__26529),
            .I(N__26526));
    CascadeBuf I__5990 (
            .O(N__26526),
            .I(N__26523));
    CascadeMux I__5989 (
            .O(N__26523),
            .I(N__26520));
    CascadeBuf I__5988 (
            .O(N__26520),
            .I(N__26517));
    CascadeMux I__5987 (
            .O(N__26517),
            .I(N__26514));
    CascadeBuf I__5986 (
            .O(N__26514),
            .I(N__26511));
    CascadeMux I__5985 (
            .O(N__26511),
            .I(N__26508));
    CascadeBuf I__5984 (
            .O(N__26508),
            .I(N__26505));
    CascadeMux I__5983 (
            .O(N__26505),
            .I(N__26502));
    CascadeBuf I__5982 (
            .O(N__26502),
            .I(N__26499));
    CascadeMux I__5981 (
            .O(N__26499),
            .I(N__26496));
    CascadeBuf I__5980 (
            .O(N__26496),
            .I(N__26493));
    CascadeMux I__5979 (
            .O(N__26493),
            .I(N__26490));
    CascadeBuf I__5978 (
            .O(N__26490),
            .I(N__26487));
    CascadeMux I__5977 (
            .O(N__26487),
            .I(N__26484));
    CascadeBuf I__5976 (
            .O(N__26484),
            .I(N__26481));
    CascadeMux I__5975 (
            .O(N__26481),
            .I(N__26478));
    CascadeBuf I__5974 (
            .O(N__26478),
            .I(N__26475));
    CascadeMux I__5973 (
            .O(N__26475),
            .I(N__26472));
    CascadeBuf I__5972 (
            .O(N__26472),
            .I(N__26469));
    CascadeMux I__5971 (
            .O(N__26469),
            .I(N__26466));
    InMux I__5970 (
            .O(N__26466),
            .I(N__26463));
    LocalMux I__5969 (
            .O(N__26463),
            .I(N__26460));
    Span4Mux_h I__5968 (
            .O(N__26460),
            .I(N__26454));
    CascadeMux I__5967 (
            .O(N__26459),
            .I(N__26451));
    CascadeMux I__5966 (
            .O(N__26458),
            .I(N__26448));
    InMux I__5965 (
            .O(N__26457),
            .I(N__26445));
    Sp12to4 I__5964 (
            .O(N__26454),
            .I(N__26442));
    InMux I__5963 (
            .O(N__26451),
            .I(N__26439));
    InMux I__5962 (
            .O(N__26448),
            .I(N__26436));
    LocalMux I__5961 (
            .O(N__26445),
            .I(N__26431));
    Span12Mux_s8_v I__5960 (
            .O(N__26442),
            .I(N__26431));
    LocalMux I__5959 (
            .O(N__26439),
            .I(M_this_sprites_address_qZ0Z_0));
    LocalMux I__5958 (
            .O(N__26436),
            .I(M_this_sprites_address_qZ0Z_0));
    Odrv12 I__5957 (
            .O(N__26431),
            .I(M_this_sprites_address_qZ0Z_0));
    InMux I__5956 (
            .O(N__26424),
            .I(N__26421));
    LocalMux I__5955 (
            .O(N__26421),
            .I(N__26418));
    Odrv4 I__5954 (
            .O(N__26418),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_9 ));
    InMux I__5953 (
            .O(N__26415),
            .I(N__26412));
    LocalMux I__5952 (
            .O(N__26412),
            .I(un1_M_this_sprites_address_q_cry_8_THRU_CO));
    CascadeMux I__5951 (
            .O(N__26409),
            .I(N__26406));
    CascadeBuf I__5950 (
            .O(N__26406),
            .I(N__26403));
    CascadeMux I__5949 (
            .O(N__26403),
            .I(N__26400));
    CascadeBuf I__5948 (
            .O(N__26400),
            .I(N__26397));
    CascadeMux I__5947 (
            .O(N__26397),
            .I(N__26394));
    CascadeBuf I__5946 (
            .O(N__26394),
            .I(N__26391));
    CascadeMux I__5945 (
            .O(N__26391),
            .I(N__26388));
    CascadeBuf I__5944 (
            .O(N__26388),
            .I(N__26385));
    CascadeMux I__5943 (
            .O(N__26385),
            .I(N__26382));
    CascadeBuf I__5942 (
            .O(N__26382),
            .I(N__26379));
    CascadeMux I__5941 (
            .O(N__26379),
            .I(N__26376));
    CascadeBuf I__5940 (
            .O(N__26376),
            .I(N__26373));
    CascadeMux I__5939 (
            .O(N__26373),
            .I(N__26370));
    CascadeBuf I__5938 (
            .O(N__26370),
            .I(N__26367));
    CascadeMux I__5937 (
            .O(N__26367),
            .I(N__26364));
    CascadeBuf I__5936 (
            .O(N__26364),
            .I(N__26361));
    CascadeMux I__5935 (
            .O(N__26361),
            .I(N__26358));
    CascadeBuf I__5934 (
            .O(N__26358),
            .I(N__26355));
    CascadeMux I__5933 (
            .O(N__26355),
            .I(N__26352));
    CascadeBuf I__5932 (
            .O(N__26352),
            .I(N__26349));
    CascadeMux I__5931 (
            .O(N__26349),
            .I(N__26346));
    CascadeBuf I__5930 (
            .O(N__26346),
            .I(N__26343));
    CascadeMux I__5929 (
            .O(N__26343),
            .I(N__26340));
    CascadeBuf I__5928 (
            .O(N__26340),
            .I(N__26337));
    CascadeMux I__5927 (
            .O(N__26337),
            .I(N__26334));
    CascadeBuf I__5926 (
            .O(N__26334),
            .I(N__26331));
    CascadeMux I__5925 (
            .O(N__26331),
            .I(N__26328));
    CascadeBuf I__5924 (
            .O(N__26328),
            .I(N__26325));
    CascadeMux I__5923 (
            .O(N__26325),
            .I(N__26322));
    CascadeBuf I__5922 (
            .O(N__26322),
            .I(N__26319));
    CascadeMux I__5921 (
            .O(N__26319),
            .I(N__26316));
    InMux I__5920 (
            .O(N__26316),
            .I(N__26313));
    LocalMux I__5919 (
            .O(N__26313),
            .I(N__26310));
    Span4Mux_h I__5918 (
            .O(N__26310),
            .I(N__26305));
    CascadeMux I__5917 (
            .O(N__26309),
            .I(N__26302));
    InMux I__5916 (
            .O(N__26308),
            .I(N__26298));
    Sp12to4 I__5915 (
            .O(N__26305),
            .I(N__26295));
    InMux I__5914 (
            .O(N__26302),
            .I(N__26292));
    InMux I__5913 (
            .O(N__26301),
            .I(N__26289));
    LocalMux I__5912 (
            .O(N__26298),
            .I(N__26286));
    Span12Mux_s7_v I__5911 (
            .O(N__26295),
            .I(N__26283));
    LocalMux I__5910 (
            .O(N__26292),
            .I(M_this_sprites_address_qZ0Z_9));
    LocalMux I__5909 (
            .O(N__26289),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv4 I__5908 (
            .O(N__26286),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv12 I__5907 (
            .O(N__26283),
            .I(M_this_sprites_address_qZ0Z_9));
    InMux I__5906 (
            .O(N__26274),
            .I(N__26267));
    InMux I__5905 (
            .O(N__26273),
            .I(N__26264));
    InMux I__5904 (
            .O(N__26272),
            .I(N__26259));
    InMux I__5903 (
            .O(N__26271),
            .I(N__26259));
    InMux I__5902 (
            .O(N__26270),
            .I(N__26256));
    LocalMux I__5901 (
            .O(N__26267),
            .I(N__26252));
    LocalMux I__5900 (
            .O(N__26264),
            .I(N__26245));
    LocalMux I__5899 (
            .O(N__26259),
            .I(N__26245));
    LocalMux I__5898 (
            .O(N__26256),
            .I(N__26245));
    InMux I__5897 (
            .O(N__26255),
            .I(N__26242));
    Span4Mux_h I__5896 (
            .O(N__26252),
            .I(N__26239));
    Span4Mux_v I__5895 (
            .O(N__26245),
            .I(N__26236));
    LocalMux I__5894 (
            .O(N__26242),
            .I(N__26233));
    Odrv4 I__5893 (
            .O(N__26239),
            .I(\this_start_data_delay.N_86_0 ));
    Odrv4 I__5892 (
            .O(N__26236),
            .I(\this_start_data_delay.N_86_0 ));
    Odrv4 I__5891 (
            .O(N__26233),
            .I(\this_start_data_delay.N_86_0 ));
    CascadeMux I__5890 (
            .O(N__26226),
            .I(N__26219));
    CascadeMux I__5889 (
            .O(N__26225),
            .I(N__26215));
    InMux I__5888 (
            .O(N__26224),
            .I(N__26175));
    InMux I__5887 (
            .O(N__26223),
            .I(N__26175));
    InMux I__5886 (
            .O(N__26222),
            .I(N__26172));
    InMux I__5885 (
            .O(N__26219),
            .I(N__26169));
    InMux I__5884 (
            .O(N__26218),
            .I(N__26166));
    InMux I__5883 (
            .O(N__26215),
            .I(N__26161));
    InMux I__5882 (
            .O(N__26214),
            .I(N__26161));
    InMux I__5881 (
            .O(N__26213),
            .I(N__26156));
    InMux I__5880 (
            .O(N__26212),
            .I(N__26156));
    InMux I__5879 (
            .O(N__26211),
            .I(N__26153));
    InMux I__5878 (
            .O(N__26210),
            .I(N__26148));
    InMux I__5877 (
            .O(N__26209),
            .I(N__26148));
    InMux I__5876 (
            .O(N__26208),
            .I(N__26143));
    InMux I__5875 (
            .O(N__26207),
            .I(N__26143));
    InMux I__5874 (
            .O(N__26206),
            .I(N__26140));
    InMux I__5873 (
            .O(N__26205),
            .I(N__26137));
    InMux I__5872 (
            .O(N__26204),
            .I(N__26134));
    InMux I__5871 (
            .O(N__26203),
            .I(N__26131));
    InMux I__5870 (
            .O(N__26202),
            .I(N__26126));
    InMux I__5869 (
            .O(N__26201),
            .I(N__26126));
    InMux I__5868 (
            .O(N__26200),
            .I(N__26123));
    InMux I__5867 (
            .O(N__26199),
            .I(N__26120));
    InMux I__5866 (
            .O(N__26198),
            .I(N__26115));
    InMux I__5865 (
            .O(N__26197),
            .I(N__26115));
    InMux I__5864 (
            .O(N__26196),
            .I(N__26112));
    InMux I__5863 (
            .O(N__26195),
            .I(N__26107));
    InMux I__5862 (
            .O(N__26194),
            .I(N__26107));
    InMux I__5861 (
            .O(N__26193),
            .I(N__26102));
    InMux I__5860 (
            .O(N__26192),
            .I(N__26102));
    InMux I__5859 (
            .O(N__26191),
            .I(N__26097));
    InMux I__5858 (
            .O(N__26190),
            .I(N__26097));
    InMux I__5857 (
            .O(N__26189),
            .I(N__26090));
    InMux I__5856 (
            .O(N__26188),
            .I(N__26090));
    InMux I__5855 (
            .O(N__26187),
            .I(N__26090));
    InMux I__5854 (
            .O(N__26186),
            .I(N__26085));
    InMux I__5853 (
            .O(N__26185),
            .I(N__26085));
    InMux I__5852 (
            .O(N__26184),
            .I(N__26082));
    InMux I__5851 (
            .O(N__26183),
            .I(N__26077));
    InMux I__5850 (
            .O(N__26182),
            .I(N__26077));
    InMux I__5849 (
            .O(N__26181),
            .I(N__26072));
    InMux I__5848 (
            .O(N__26180),
            .I(N__26072));
    LocalMux I__5847 (
            .O(N__26175),
            .I(N__26041));
    LocalMux I__5846 (
            .O(N__26172),
            .I(N__26038));
    LocalMux I__5845 (
            .O(N__26169),
            .I(N__26035));
    LocalMux I__5844 (
            .O(N__26166),
            .I(N__26032));
    LocalMux I__5843 (
            .O(N__26161),
            .I(N__26029));
    LocalMux I__5842 (
            .O(N__26156),
            .I(N__26026));
    LocalMux I__5841 (
            .O(N__26153),
            .I(N__26023));
    LocalMux I__5840 (
            .O(N__26148),
            .I(N__26020));
    LocalMux I__5839 (
            .O(N__26143),
            .I(N__26017));
    LocalMux I__5838 (
            .O(N__26140),
            .I(N__26014));
    LocalMux I__5837 (
            .O(N__26137),
            .I(N__26011));
    LocalMux I__5836 (
            .O(N__26134),
            .I(N__26008));
    LocalMux I__5835 (
            .O(N__26131),
            .I(N__26005));
    LocalMux I__5834 (
            .O(N__26126),
            .I(N__26002));
    LocalMux I__5833 (
            .O(N__26123),
            .I(N__25999));
    LocalMux I__5832 (
            .O(N__26120),
            .I(N__25996));
    LocalMux I__5831 (
            .O(N__26115),
            .I(N__25993));
    LocalMux I__5830 (
            .O(N__26112),
            .I(N__25990));
    LocalMux I__5829 (
            .O(N__26107),
            .I(N__25987));
    LocalMux I__5828 (
            .O(N__26102),
            .I(N__25984));
    LocalMux I__5827 (
            .O(N__26097),
            .I(N__25981));
    LocalMux I__5826 (
            .O(N__26090),
            .I(N__25978));
    LocalMux I__5825 (
            .O(N__26085),
            .I(N__25975));
    LocalMux I__5824 (
            .O(N__26082),
            .I(N__25972));
    LocalMux I__5823 (
            .O(N__26077),
            .I(N__25969));
    LocalMux I__5822 (
            .O(N__26072),
            .I(N__25966));
    SRMux I__5821 (
            .O(N__26071),
            .I(N__25857));
    SRMux I__5820 (
            .O(N__26070),
            .I(N__25857));
    SRMux I__5819 (
            .O(N__26069),
            .I(N__25857));
    SRMux I__5818 (
            .O(N__26068),
            .I(N__25857));
    SRMux I__5817 (
            .O(N__26067),
            .I(N__25857));
    SRMux I__5816 (
            .O(N__26066),
            .I(N__25857));
    SRMux I__5815 (
            .O(N__26065),
            .I(N__25857));
    SRMux I__5814 (
            .O(N__26064),
            .I(N__25857));
    SRMux I__5813 (
            .O(N__26063),
            .I(N__25857));
    SRMux I__5812 (
            .O(N__26062),
            .I(N__25857));
    SRMux I__5811 (
            .O(N__26061),
            .I(N__25857));
    SRMux I__5810 (
            .O(N__26060),
            .I(N__25857));
    SRMux I__5809 (
            .O(N__26059),
            .I(N__25857));
    SRMux I__5808 (
            .O(N__26058),
            .I(N__25857));
    SRMux I__5807 (
            .O(N__26057),
            .I(N__25857));
    SRMux I__5806 (
            .O(N__26056),
            .I(N__25857));
    SRMux I__5805 (
            .O(N__26055),
            .I(N__25857));
    SRMux I__5804 (
            .O(N__26054),
            .I(N__25857));
    SRMux I__5803 (
            .O(N__26053),
            .I(N__25857));
    SRMux I__5802 (
            .O(N__26052),
            .I(N__25857));
    SRMux I__5801 (
            .O(N__26051),
            .I(N__25857));
    SRMux I__5800 (
            .O(N__26050),
            .I(N__25857));
    SRMux I__5799 (
            .O(N__26049),
            .I(N__25857));
    SRMux I__5798 (
            .O(N__26048),
            .I(N__25857));
    SRMux I__5797 (
            .O(N__26047),
            .I(N__25857));
    SRMux I__5796 (
            .O(N__26046),
            .I(N__25857));
    SRMux I__5795 (
            .O(N__26045),
            .I(N__25857));
    SRMux I__5794 (
            .O(N__26044),
            .I(N__25857));
    Glb2LocalMux I__5793 (
            .O(N__26041),
            .I(N__25857));
    Glb2LocalMux I__5792 (
            .O(N__26038),
            .I(N__25857));
    Glb2LocalMux I__5791 (
            .O(N__26035),
            .I(N__25857));
    Glb2LocalMux I__5790 (
            .O(N__26032),
            .I(N__25857));
    Glb2LocalMux I__5789 (
            .O(N__26029),
            .I(N__25857));
    Glb2LocalMux I__5788 (
            .O(N__26026),
            .I(N__25857));
    Glb2LocalMux I__5787 (
            .O(N__26023),
            .I(N__25857));
    Glb2LocalMux I__5786 (
            .O(N__26020),
            .I(N__25857));
    Glb2LocalMux I__5785 (
            .O(N__26017),
            .I(N__25857));
    Glb2LocalMux I__5784 (
            .O(N__26014),
            .I(N__25857));
    Glb2LocalMux I__5783 (
            .O(N__26011),
            .I(N__25857));
    Glb2LocalMux I__5782 (
            .O(N__26008),
            .I(N__25857));
    Glb2LocalMux I__5781 (
            .O(N__26005),
            .I(N__25857));
    Glb2LocalMux I__5780 (
            .O(N__26002),
            .I(N__25857));
    Glb2LocalMux I__5779 (
            .O(N__25999),
            .I(N__25857));
    Glb2LocalMux I__5778 (
            .O(N__25996),
            .I(N__25857));
    Glb2LocalMux I__5777 (
            .O(N__25993),
            .I(N__25857));
    Glb2LocalMux I__5776 (
            .O(N__25990),
            .I(N__25857));
    Glb2LocalMux I__5775 (
            .O(N__25987),
            .I(N__25857));
    Glb2LocalMux I__5774 (
            .O(N__25984),
            .I(N__25857));
    Glb2LocalMux I__5773 (
            .O(N__25981),
            .I(N__25857));
    Glb2LocalMux I__5772 (
            .O(N__25978),
            .I(N__25857));
    Glb2LocalMux I__5771 (
            .O(N__25975),
            .I(N__25857));
    Glb2LocalMux I__5770 (
            .O(N__25972),
            .I(N__25857));
    Glb2LocalMux I__5769 (
            .O(N__25969),
            .I(N__25857));
    Glb2LocalMux I__5768 (
            .O(N__25966),
            .I(N__25857));
    GlobalMux I__5767 (
            .O(N__25857),
            .I(N__25854));
    gio2CtrlBuf I__5766 (
            .O(N__25854),
            .I(M_this_reset_cond_out_g_0));
    InMux I__5765 (
            .O(N__25851),
            .I(N__25848));
    LocalMux I__5764 (
            .O(N__25848),
            .I(N__25845));
    Span4Mux_h I__5763 (
            .O(N__25845),
            .I(N__25842));
    Odrv4 I__5762 (
            .O(N__25842),
            .I(\this_sprites_ram.mem_out_bus5_3 ));
    InMux I__5761 (
            .O(N__25839),
            .I(N__25836));
    LocalMux I__5760 (
            .O(N__25836),
            .I(N__25833));
    Span12Mux_h I__5759 (
            .O(N__25833),
            .I(N__25830));
    Span12Mux_v I__5758 (
            .O(N__25830),
            .I(N__25827));
    Odrv12 I__5757 (
            .O(N__25827),
            .I(\this_sprites_ram.mem_out_bus1_3 ));
    CascadeMux I__5756 (
            .O(N__25824),
            .I(N__25821));
    CascadeBuf I__5755 (
            .O(N__25821),
            .I(N__25818));
    CascadeMux I__5754 (
            .O(N__25818),
            .I(N__25815));
    CascadeBuf I__5753 (
            .O(N__25815),
            .I(N__25812));
    CascadeMux I__5752 (
            .O(N__25812),
            .I(N__25809));
    CascadeBuf I__5751 (
            .O(N__25809),
            .I(N__25806));
    CascadeMux I__5750 (
            .O(N__25806),
            .I(N__25803));
    CascadeBuf I__5749 (
            .O(N__25803),
            .I(N__25800));
    CascadeMux I__5748 (
            .O(N__25800),
            .I(N__25797));
    CascadeBuf I__5747 (
            .O(N__25797),
            .I(N__25794));
    CascadeMux I__5746 (
            .O(N__25794),
            .I(N__25791));
    CascadeBuf I__5745 (
            .O(N__25791),
            .I(N__25788));
    CascadeMux I__5744 (
            .O(N__25788),
            .I(N__25785));
    CascadeBuf I__5743 (
            .O(N__25785),
            .I(N__25782));
    CascadeMux I__5742 (
            .O(N__25782),
            .I(N__25779));
    CascadeBuf I__5741 (
            .O(N__25779),
            .I(N__25776));
    CascadeMux I__5740 (
            .O(N__25776),
            .I(N__25773));
    CascadeBuf I__5739 (
            .O(N__25773),
            .I(N__25770));
    CascadeMux I__5738 (
            .O(N__25770),
            .I(N__25767));
    CascadeBuf I__5737 (
            .O(N__25767),
            .I(N__25764));
    CascadeMux I__5736 (
            .O(N__25764),
            .I(N__25761));
    CascadeBuf I__5735 (
            .O(N__25761),
            .I(N__25758));
    CascadeMux I__5734 (
            .O(N__25758),
            .I(N__25755));
    CascadeBuf I__5733 (
            .O(N__25755),
            .I(N__25752));
    CascadeMux I__5732 (
            .O(N__25752),
            .I(N__25749));
    CascadeBuf I__5731 (
            .O(N__25749),
            .I(N__25746));
    CascadeMux I__5730 (
            .O(N__25746),
            .I(N__25743));
    CascadeBuf I__5729 (
            .O(N__25743),
            .I(N__25740));
    CascadeMux I__5728 (
            .O(N__25740),
            .I(N__25737));
    CascadeBuf I__5727 (
            .O(N__25737),
            .I(N__25734));
    CascadeMux I__5726 (
            .O(N__25734),
            .I(N__25731));
    InMux I__5725 (
            .O(N__25731),
            .I(N__25728));
    LocalMux I__5724 (
            .O(N__25728),
            .I(N__25725));
    Span4Mux_h I__5723 (
            .O(N__25725),
            .I(N__25722));
    Sp12to4 I__5722 (
            .O(N__25722),
            .I(N__25716));
    InMux I__5721 (
            .O(N__25721),
            .I(N__25713));
    InMux I__5720 (
            .O(N__25720),
            .I(N__25708));
    InMux I__5719 (
            .O(N__25719),
            .I(N__25708));
    Span12Mux_s6_v I__5718 (
            .O(N__25716),
            .I(N__25705));
    LocalMux I__5717 (
            .O(N__25713),
            .I(M_this_sprites_address_qZ0Z_6));
    LocalMux I__5716 (
            .O(N__25708),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv12 I__5715 (
            .O(N__25705),
            .I(M_this_sprites_address_qZ0Z_6));
    InMux I__5714 (
            .O(N__25698),
            .I(N__25695));
    LocalMux I__5713 (
            .O(N__25695),
            .I(un1_M_this_sprites_address_q_cry_5_THRU_CO));
    InMux I__5712 (
            .O(N__25692),
            .I(un1_M_this_sprites_address_q_cry_5));
    CascadeMux I__5711 (
            .O(N__25689),
            .I(N__25686));
    CascadeBuf I__5710 (
            .O(N__25686),
            .I(N__25683));
    CascadeMux I__5709 (
            .O(N__25683),
            .I(N__25680));
    CascadeBuf I__5708 (
            .O(N__25680),
            .I(N__25677));
    CascadeMux I__5707 (
            .O(N__25677),
            .I(N__25674));
    CascadeBuf I__5706 (
            .O(N__25674),
            .I(N__25671));
    CascadeMux I__5705 (
            .O(N__25671),
            .I(N__25668));
    CascadeBuf I__5704 (
            .O(N__25668),
            .I(N__25665));
    CascadeMux I__5703 (
            .O(N__25665),
            .I(N__25662));
    CascadeBuf I__5702 (
            .O(N__25662),
            .I(N__25659));
    CascadeMux I__5701 (
            .O(N__25659),
            .I(N__25656));
    CascadeBuf I__5700 (
            .O(N__25656),
            .I(N__25653));
    CascadeMux I__5699 (
            .O(N__25653),
            .I(N__25650));
    CascadeBuf I__5698 (
            .O(N__25650),
            .I(N__25647));
    CascadeMux I__5697 (
            .O(N__25647),
            .I(N__25644));
    CascadeBuf I__5696 (
            .O(N__25644),
            .I(N__25641));
    CascadeMux I__5695 (
            .O(N__25641),
            .I(N__25638));
    CascadeBuf I__5694 (
            .O(N__25638),
            .I(N__25635));
    CascadeMux I__5693 (
            .O(N__25635),
            .I(N__25632));
    CascadeBuf I__5692 (
            .O(N__25632),
            .I(N__25629));
    CascadeMux I__5691 (
            .O(N__25629),
            .I(N__25626));
    CascadeBuf I__5690 (
            .O(N__25626),
            .I(N__25623));
    CascadeMux I__5689 (
            .O(N__25623),
            .I(N__25620));
    CascadeBuf I__5688 (
            .O(N__25620),
            .I(N__25617));
    CascadeMux I__5687 (
            .O(N__25617),
            .I(N__25614));
    CascadeBuf I__5686 (
            .O(N__25614),
            .I(N__25611));
    CascadeMux I__5685 (
            .O(N__25611),
            .I(N__25608));
    CascadeBuf I__5684 (
            .O(N__25608),
            .I(N__25605));
    CascadeMux I__5683 (
            .O(N__25605),
            .I(N__25602));
    CascadeBuf I__5682 (
            .O(N__25602),
            .I(N__25599));
    CascadeMux I__5681 (
            .O(N__25599),
            .I(N__25596));
    InMux I__5680 (
            .O(N__25596),
            .I(N__25593));
    LocalMux I__5679 (
            .O(N__25593),
            .I(N__25590));
    Span4Mux_h I__5678 (
            .O(N__25590),
            .I(N__25585));
    CascadeMux I__5677 (
            .O(N__25589),
            .I(N__25582));
    CascadeMux I__5676 (
            .O(N__25588),
            .I(N__25579));
    Sp12to4 I__5675 (
            .O(N__25585),
            .I(N__25575));
    InMux I__5674 (
            .O(N__25582),
            .I(N__25572));
    InMux I__5673 (
            .O(N__25579),
            .I(N__25569));
    InMux I__5672 (
            .O(N__25578),
            .I(N__25566));
    Span12Mux_s8_v I__5671 (
            .O(N__25575),
            .I(N__25563));
    LocalMux I__5670 (
            .O(N__25572),
            .I(M_this_sprites_address_qZ0Z_7));
    LocalMux I__5669 (
            .O(N__25569),
            .I(M_this_sprites_address_qZ0Z_7));
    LocalMux I__5668 (
            .O(N__25566),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv12 I__5667 (
            .O(N__25563),
            .I(M_this_sprites_address_qZ0Z_7));
    InMux I__5666 (
            .O(N__25554),
            .I(N__25551));
    LocalMux I__5665 (
            .O(N__25551),
            .I(un1_M_this_sprites_address_q_cry_6_THRU_CO));
    InMux I__5664 (
            .O(N__25548),
            .I(un1_M_this_sprites_address_q_cry_6));
    InMux I__5663 (
            .O(N__25545),
            .I(bfn_23_18_0_));
    InMux I__5662 (
            .O(N__25542),
            .I(un1_M_this_sprites_address_q_cry_8));
    CascadeMux I__5661 (
            .O(N__25539),
            .I(N__25536));
    CascadeBuf I__5660 (
            .O(N__25536),
            .I(N__25533));
    CascadeMux I__5659 (
            .O(N__25533),
            .I(N__25530));
    CascadeBuf I__5658 (
            .O(N__25530),
            .I(N__25527));
    CascadeMux I__5657 (
            .O(N__25527),
            .I(N__25524));
    CascadeBuf I__5656 (
            .O(N__25524),
            .I(N__25521));
    CascadeMux I__5655 (
            .O(N__25521),
            .I(N__25518));
    CascadeBuf I__5654 (
            .O(N__25518),
            .I(N__25515));
    CascadeMux I__5653 (
            .O(N__25515),
            .I(N__25512));
    CascadeBuf I__5652 (
            .O(N__25512),
            .I(N__25509));
    CascadeMux I__5651 (
            .O(N__25509),
            .I(N__25506));
    CascadeBuf I__5650 (
            .O(N__25506),
            .I(N__25503));
    CascadeMux I__5649 (
            .O(N__25503),
            .I(N__25500));
    CascadeBuf I__5648 (
            .O(N__25500),
            .I(N__25497));
    CascadeMux I__5647 (
            .O(N__25497),
            .I(N__25494));
    CascadeBuf I__5646 (
            .O(N__25494),
            .I(N__25491));
    CascadeMux I__5645 (
            .O(N__25491),
            .I(N__25488));
    CascadeBuf I__5644 (
            .O(N__25488),
            .I(N__25485));
    CascadeMux I__5643 (
            .O(N__25485),
            .I(N__25482));
    CascadeBuf I__5642 (
            .O(N__25482),
            .I(N__25479));
    CascadeMux I__5641 (
            .O(N__25479),
            .I(N__25476));
    CascadeBuf I__5640 (
            .O(N__25476),
            .I(N__25473));
    CascadeMux I__5639 (
            .O(N__25473),
            .I(N__25470));
    CascadeBuf I__5638 (
            .O(N__25470),
            .I(N__25467));
    CascadeMux I__5637 (
            .O(N__25467),
            .I(N__25464));
    CascadeBuf I__5636 (
            .O(N__25464),
            .I(N__25461));
    CascadeMux I__5635 (
            .O(N__25461),
            .I(N__25458));
    CascadeBuf I__5634 (
            .O(N__25458),
            .I(N__25455));
    CascadeMux I__5633 (
            .O(N__25455),
            .I(N__25452));
    CascadeBuf I__5632 (
            .O(N__25452),
            .I(N__25449));
    CascadeMux I__5631 (
            .O(N__25449),
            .I(N__25446));
    InMux I__5630 (
            .O(N__25446),
            .I(N__25443));
    LocalMux I__5629 (
            .O(N__25443),
            .I(N__25440));
    Span4Mux_h I__5628 (
            .O(N__25440),
            .I(N__25437));
    Sp12to4 I__5627 (
            .O(N__25437),
            .I(N__25431));
    InMux I__5626 (
            .O(N__25436),
            .I(N__25428));
    InMux I__5625 (
            .O(N__25435),
            .I(N__25423));
    InMux I__5624 (
            .O(N__25434),
            .I(N__25423));
    Span12Mux_s5_v I__5623 (
            .O(N__25431),
            .I(N__25420));
    LocalMux I__5622 (
            .O(N__25428),
            .I(M_this_sprites_address_qZ0Z_10));
    LocalMux I__5621 (
            .O(N__25423),
            .I(M_this_sprites_address_qZ0Z_10));
    Odrv12 I__5620 (
            .O(N__25420),
            .I(M_this_sprites_address_qZ0Z_10));
    InMux I__5619 (
            .O(N__25413),
            .I(N__25410));
    LocalMux I__5618 (
            .O(N__25410),
            .I(un1_M_this_sprites_address_q_cry_9_THRU_CO));
    InMux I__5617 (
            .O(N__25407),
            .I(un1_M_this_sprites_address_q_cry_9));
    InMux I__5616 (
            .O(N__25404),
            .I(N__25401));
    LocalMux I__5615 (
            .O(N__25401),
            .I(un1_M_this_sprites_address_q_cry_10_THRU_CO));
    InMux I__5614 (
            .O(N__25398),
            .I(un1_M_this_sprites_address_q_cry_10));
    InMux I__5613 (
            .O(N__25395),
            .I(N__25392));
    LocalMux I__5612 (
            .O(N__25392),
            .I(un1_M_this_sprites_address_q_cry_11_THRU_CO));
    InMux I__5611 (
            .O(N__25389),
            .I(un1_M_this_sprites_address_q_cry_11));
    InMux I__5610 (
            .O(N__25386),
            .I(N__25383));
    LocalMux I__5609 (
            .O(N__25383),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_13 ));
    InMux I__5608 (
            .O(N__25380),
            .I(un1_M_this_sprites_address_q_cry_12));
    InMux I__5607 (
            .O(N__25377),
            .I(N__25374));
    LocalMux I__5606 (
            .O(N__25374),
            .I(N__25371));
    Odrv4 I__5605 (
            .O(N__25371),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_0 ));
    InMux I__5604 (
            .O(N__25368),
            .I(N__25364));
    InMux I__5603 (
            .O(N__25367),
            .I(N__25361));
    LocalMux I__5602 (
            .O(N__25364),
            .I(un30_0));
    LocalMux I__5601 (
            .O(N__25361),
            .I(un30_0));
    CascadeMux I__5600 (
            .O(N__25356),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_1_cascade_ ));
    InMux I__5599 (
            .O(N__25353),
            .I(N__25347));
    InMux I__5598 (
            .O(N__25352),
            .I(N__25347));
    LocalMux I__5597 (
            .O(N__25347),
            .I(N__25340));
    InMux I__5596 (
            .O(N__25346),
            .I(N__25331));
    InMux I__5595 (
            .O(N__25345),
            .I(N__25331));
    InMux I__5594 (
            .O(N__25344),
            .I(N__25331));
    InMux I__5593 (
            .O(N__25343),
            .I(N__25331));
    Span4Mux_v I__5592 (
            .O(N__25340),
            .I(N__25327));
    LocalMux I__5591 (
            .O(N__25331),
            .I(N__25324));
    InMux I__5590 (
            .O(N__25330),
            .I(N__25321));
    Odrv4 I__5589 (
            .O(N__25327),
            .I(\this_start_data_delay.N_993 ));
    Odrv4 I__5588 (
            .O(N__25324),
            .I(\this_start_data_delay.N_993 ));
    LocalMux I__5587 (
            .O(N__25321),
            .I(\this_start_data_delay.N_993 ));
    CascadeMux I__5586 (
            .O(N__25314),
            .I(N__25309));
    CascadeMux I__5585 (
            .O(N__25313),
            .I(N__25306));
    CascadeMux I__5584 (
            .O(N__25312),
            .I(N__25303));
    InMux I__5583 (
            .O(N__25309),
            .I(N__25291));
    InMux I__5582 (
            .O(N__25306),
            .I(N__25291));
    InMux I__5581 (
            .O(N__25303),
            .I(N__25291));
    InMux I__5580 (
            .O(N__25302),
            .I(N__25291));
    InMux I__5579 (
            .O(N__25301),
            .I(N__25286));
    InMux I__5578 (
            .O(N__25300),
            .I(N__25286));
    LocalMux I__5577 (
            .O(N__25291),
            .I(N__25283));
    LocalMux I__5576 (
            .O(N__25286),
            .I(N__25280));
    Span4Mux_v I__5575 (
            .O(N__25283),
            .I(N__25277));
    Odrv4 I__5574 (
            .O(N__25280),
            .I(\this_start_data_delay.N_109 ));
    Odrv4 I__5573 (
            .O(N__25277),
            .I(\this_start_data_delay.N_109 ));
    CascadeMux I__5572 (
            .O(N__25272),
            .I(N__25269));
    CascadeBuf I__5571 (
            .O(N__25269),
            .I(N__25266));
    CascadeMux I__5570 (
            .O(N__25266),
            .I(N__25263));
    CascadeBuf I__5569 (
            .O(N__25263),
            .I(N__25260));
    CascadeMux I__5568 (
            .O(N__25260),
            .I(N__25257));
    CascadeBuf I__5567 (
            .O(N__25257),
            .I(N__25254));
    CascadeMux I__5566 (
            .O(N__25254),
            .I(N__25251));
    CascadeBuf I__5565 (
            .O(N__25251),
            .I(N__25248));
    CascadeMux I__5564 (
            .O(N__25248),
            .I(N__25245));
    CascadeBuf I__5563 (
            .O(N__25245),
            .I(N__25242));
    CascadeMux I__5562 (
            .O(N__25242),
            .I(N__25239));
    CascadeBuf I__5561 (
            .O(N__25239),
            .I(N__25236));
    CascadeMux I__5560 (
            .O(N__25236),
            .I(N__25233));
    CascadeBuf I__5559 (
            .O(N__25233),
            .I(N__25230));
    CascadeMux I__5558 (
            .O(N__25230),
            .I(N__25227));
    CascadeBuf I__5557 (
            .O(N__25227),
            .I(N__25224));
    CascadeMux I__5556 (
            .O(N__25224),
            .I(N__25221));
    CascadeBuf I__5555 (
            .O(N__25221),
            .I(N__25218));
    CascadeMux I__5554 (
            .O(N__25218),
            .I(N__25215));
    CascadeBuf I__5553 (
            .O(N__25215),
            .I(N__25212));
    CascadeMux I__5552 (
            .O(N__25212),
            .I(N__25209));
    CascadeBuf I__5551 (
            .O(N__25209),
            .I(N__25206));
    CascadeMux I__5550 (
            .O(N__25206),
            .I(N__25203));
    CascadeBuf I__5549 (
            .O(N__25203),
            .I(N__25200));
    CascadeMux I__5548 (
            .O(N__25200),
            .I(N__25197));
    CascadeBuf I__5547 (
            .O(N__25197),
            .I(N__25194));
    CascadeMux I__5546 (
            .O(N__25194),
            .I(N__25191));
    CascadeBuf I__5545 (
            .O(N__25191),
            .I(N__25188));
    CascadeMux I__5544 (
            .O(N__25188),
            .I(N__25185));
    CascadeBuf I__5543 (
            .O(N__25185),
            .I(N__25182));
    CascadeMux I__5542 (
            .O(N__25182),
            .I(N__25179));
    InMux I__5541 (
            .O(N__25179),
            .I(N__25176));
    LocalMux I__5540 (
            .O(N__25176),
            .I(N__25172));
    CascadeMux I__5539 (
            .O(N__25175),
            .I(N__25169));
    Span12Mux_s4_v I__5538 (
            .O(N__25172),
            .I(N__25164));
    InMux I__5537 (
            .O(N__25169),
            .I(N__25161));
    InMux I__5536 (
            .O(N__25168),
            .I(N__25156));
    InMux I__5535 (
            .O(N__25167),
            .I(N__25156));
    Span12Mux_v I__5534 (
            .O(N__25164),
            .I(N__25153));
    LocalMux I__5533 (
            .O(N__25161),
            .I(M_this_sprites_address_qZ0Z_1));
    LocalMux I__5532 (
            .O(N__25156),
            .I(M_this_sprites_address_qZ0Z_1));
    Odrv12 I__5531 (
            .O(N__25153),
            .I(M_this_sprites_address_qZ0Z_1));
    InMux I__5530 (
            .O(N__25146),
            .I(N__25143));
    LocalMux I__5529 (
            .O(N__25143),
            .I(un1_M_this_sprites_address_q_cry_0_THRU_CO));
    InMux I__5528 (
            .O(N__25140),
            .I(un1_M_this_sprites_address_q_cry_0));
    CascadeMux I__5527 (
            .O(N__25137),
            .I(N__25134));
    CascadeBuf I__5526 (
            .O(N__25134),
            .I(N__25131));
    CascadeMux I__5525 (
            .O(N__25131),
            .I(N__25128));
    CascadeBuf I__5524 (
            .O(N__25128),
            .I(N__25125));
    CascadeMux I__5523 (
            .O(N__25125),
            .I(N__25122));
    CascadeBuf I__5522 (
            .O(N__25122),
            .I(N__25119));
    CascadeMux I__5521 (
            .O(N__25119),
            .I(N__25116));
    CascadeBuf I__5520 (
            .O(N__25116),
            .I(N__25113));
    CascadeMux I__5519 (
            .O(N__25113),
            .I(N__25110));
    CascadeBuf I__5518 (
            .O(N__25110),
            .I(N__25107));
    CascadeMux I__5517 (
            .O(N__25107),
            .I(N__25104));
    CascadeBuf I__5516 (
            .O(N__25104),
            .I(N__25101));
    CascadeMux I__5515 (
            .O(N__25101),
            .I(N__25098));
    CascadeBuf I__5514 (
            .O(N__25098),
            .I(N__25095));
    CascadeMux I__5513 (
            .O(N__25095),
            .I(N__25092));
    CascadeBuf I__5512 (
            .O(N__25092),
            .I(N__25089));
    CascadeMux I__5511 (
            .O(N__25089),
            .I(N__25086));
    CascadeBuf I__5510 (
            .O(N__25086),
            .I(N__25083));
    CascadeMux I__5509 (
            .O(N__25083),
            .I(N__25080));
    CascadeBuf I__5508 (
            .O(N__25080),
            .I(N__25077));
    CascadeMux I__5507 (
            .O(N__25077),
            .I(N__25074));
    CascadeBuf I__5506 (
            .O(N__25074),
            .I(N__25071));
    CascadeMux I__5505 (
            .O(N__25071),
            .I(N__25068));
    CascadeBuf I__5504 (
            .O(N__25068),
            .I(N__25065));
    CascadeMux I__5503 (
            .O(N__25065),
            .I(N__25062));
    CascadeBuf I__5502 (
            .O(N__25062),
            .I(N__25059));
    CascadeMux I__5501 (
            .O(N__25059),
            .I(N__25056));
    CascadeBuf I__5500 (
            .O(N__25056),
            .I(N__25053));
    CascadeMux I__5499 (
            .O(N__25053),
            .I(N__25050));
    CascadeBuf I__5498 (
            .O(N__25050),
            .I(N__25047));
    CascadeMux I__5497 (
            .O(N__25047),
            .I(N__25044));
    InMux I__5496 (
            .O(N__25044),
            .I(N__25041));
    LocalMux I__5495 (
            .O(N__25041),
            .I(N__25037));
    InMux I__5494 (
            .O(N__25040),
            .I(N__25034));
    Span12Mux_s10_h I__5493 (
            .O(N__25037),
            .I(N__25029));
    LocalMux I__5492 (
            .O(N__25034),
            .I(N__25026));
    InMux I__5491 (
            .O(N__25033),
            .I(N__25023));
    InMux I__5490 (
            .O(N__25032),
            .I(N__25020));
    Span12Mux_v I__5489 (
            .O(N__25029),
            .I(N__25017));
    Odrv4 I__5488 (
            .O(N__25026),
            .I(M_this_sprites_address_qZ0Z_2));
    LocalMux I__5487 (
            .O(N__25023),
            .I(M_this_sprites_address_qZ0Z_2));
    LocalMux I__5486 (
            .O(N__25020),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv12 I__5485 (
            .O(N__25017),
            .I(M_this_sprites_address_qZ0Z_2));
    InMux I__5484 (
            .O(N__25008),
            .I(N__25005));
    LocalMux I__5483 (
            .O(N__25005),
            .I(N__25002));
    Odrv4 I__5482 (
            .O(N__25002),
            .I(un1_M_this_sprites_address_q_cry_1_THRU_CO));
    InMux I__5481 (
            .O(N__24999),
            .I(un1_M_this_sprites_address_q_cry_1));
    CascadeMux I__5480 (
            .O(N__24996),
            .I(N__24993));
    CascadeBuf I__5479 (
            .O(N__24993),
            .I(N__24990));
    CascadeMux I__5478 (
            .O(N__24990),
            .I(N__24987));
    CascadeBuf I__5477 (
            .O(N__24987),
            .I(N__24984));
    CascadeMux I__5476 (
            .O(N__24984),
            .I(N__24981));
    CascadeBuf I__5475 (
            .O(N__24981),
            .I(N__24978));
    CascadeMux I__5474 (
            .O(N__24978),
            .I(N__24975));
    CascadeBuf I__5473 (
            .O(N__24975),
            .I(N__24972));
    CascadeMux I__5472 (
            .O(N__24972),
            .I(N__24969));
    CascadeBuf I__5471 (
            .O(N__24969),
            .I(N__24966));
    CascadeMux I__5470 (
            .O(N__24966),
            .I(N__24963));
    CascadeBuf I__5469 (
            .O(N__24963),
            .I(N__24960));
    CascadeMux I__5468 (
            .O(N__24960),
            .I(N__24957));
    CascadeBuf I__5467 (
            .O(N__24957),
            .I(N__24954));
    CascadeMux I__5466 (
            .O(N__24954),
            .I(N__24951));
    CascadeBuf I__5465 (
            .O(N__24951),
            .I(N__24948));
    CascadeMux I__5464 (
            .O(N__24948),
            .I(N__24945));
    CascadeBuf I__5463 (
            .O(N__24945),
            .I(N__24942));
    CascadeMux I__5462 (
            .O(N__24942),
            .I(N__24939));
    CascadeBuf I__5461 (
            .O(N__24939),
            .I(N__24936));
    CascadeMux I__5460 (
            .O(N__24936),
            .I(N__24933));
    CascadeBuf I__5459 (
            .O(N__24933),
            .I(N__24930));
    CascadeMux I__5458 (
            .O(N__24930),
            .I(N__24927));
    CascadeBuf I__5457 (
            .O(N__24927),
            .I(N__24924));
    CascadeMux I__5456 (
            .O(N__24924),
            .I(N__24921));
    CascadeBuf I__5455 (
            .O(N__24921),
            .I(N__24918));
    CascadeMux I__5454 (
            .O(N__24918),
            .I(N__24915));
    CascadeBuf I__5453 (
            .O(N__24915),
            .I(N__24912));
    CascadeMux I__5452 (
            .O(N__24912),
            .I(N__24909));
    CascadeBuf I__5451 (
            .O(N__24909),
            .I(N__24906));
    CascadeMux I__5450 (
            .O(N__24906),
            .I(N__24903));
    InMux I__5449 (
            .O(N__24903),
            .I(N__24899));
    InMux I__5448 (
            .O(N__24902),
            .I(N__24896));
    LocalMux I__5447 (
            .O(N__24899),
            .I(N__24893));
    LocalMux I__5446 (
            .O(N__24896),
            .I(N__24890));
    Span12Mux_s1_v I__5445 (
            .O(N__24893),
            .I(N__24885));
    Span4Mux_h I__5444 (
            .O(N__24890),
            .I(N__24882));
    InMux I__5443 (
            .O(N__24889),
            .I(N__24879));
    InMux I__5442 (
            .O(N__24888),
            .I(N__24876));
    Span12Mux_v I__5441 (
            .O(N__24885),
            .I(N__24873));
    Odrv4 I__5440 (
            .O(N__24882),
            .I(M_this_sprites_address_qZ0Z_3));
    LocalMux I__5439 (
            .O(N__24879),
            .I(M_this_sprites_address_qZ0Z_3));
    LocalMux I__5438 (
            .O(N__24876),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv12 I__5437 (
            .O(N__24873),
            .I(M_this_sprites_address_qZ0Z_3));
    InMux I__5436 (
            .O(N__24864),
            .I(N__24861));
    LocalMux I__5435 (
            .O(N__24861),
            .I(N__24858));
    Odrv4 I__5434 (
            .O(N__24858),
            .I(un1_M_this_sprites_address_q_cry_2_THRU_CO));
    InMux I__5433 (
            .O(N__24855),
            .I(un1_M_this_sprites_address_q_cry_2));
    CascadeMux I__5432 (
            .O(N__24852),
            .I(N__24849));
    CascadeBuf I__5431 (
            .O(N__24849),
            .I(N__24846));
    CascadeMux I__5430 (
            .O(N__24846),
            .I(N__24843));
    CascadeBuf I__5429 (
            .O(N__24843),
            .I(N__24840));
    CascadeMux I__5428 (
            .O(N__24840),
            .I(N__24837));
    CascadeBuf I__5427 (
            .O(N__24837),
            .I(N__24834));
    CascadeMux I__5426 (
            .O(N__24834),
            .I(N__24831));
    CascadeBuf I__5425 (
            .O(N__24831),
            .I(N__24828));
    CascadeMux I__5424 (
            .O(N__24828),
            .I(N__24825));
    CascadeBuf I__5423 (
            .O(N__24825),
            .I(N__24822));
    CascadeMux I__5422 (
            .O(N__24822),
            .I(N__24819));
    CascadeBuf I__5421 (
            .O(N__24819),
            .I(N__24816));
    CascadeMux I__5420 (
            .O(N__24816),
            .I(N__24813));
    CascadeBuf I__5419 (
            .O(N__24813),
            .I(N__24810));
    CascadeMux I__5418 (
            .O(N__24810),
            .I(N__24807));
    CascadeBuf I__5417 (
            .O(N__24807),
            .I(N__24804));
    CascadeMux I__5416 (
            .O(N__24804),
            .I(N__24801));
    CascadeBuf I__5415 (
            .O(N__24801),
            .I(N__24798));
    CascadeMux I__5414 (
            .O(N__24798),
            .I(N__24795));
    CascadeBuf I__5413 (
            .O(N__24795),
            .I(N__24792));
    CascadeMux I__5412 (
            .O(N__24792),
            .I(N__24789));
    CascadeBuf I__5411 (
            .O(N__24789),
            .I(N__24786));
    CascadeMux I__5410 (
            .O(N__24786),
            .I(N__24783));
    CascadeBuf I__5409 (
            .O(N__24783),
            .I(N__24780));
    CascadeMux I__5408 (
            .O(N__24780),
            .I(N__24777));
    CascadeBuf I__5407 (
            .O(N__24777),
            .I(N__24774));
    CascadeMux I__5406 (
            .O(N__24774),
            .I(N__24771));
    CascadeBuf I__5405 (
            .O(N__24771),
            .I(N__24768));
    CascadeMux I__5404 (
            .O(N__24768),
            .I(N__24765));
    CascadeBuf I__5403 (
            .O(N__24765),
            .I(N__24762));
    CascadeMux I__5402 (
            .O(N__24762),
            .I(N__24759));
    InMux I__5401 (
            .O(N__24759),
            .I(N__24756));
    LocalMux I__5400 (
            .O(N__24756),
            .I(N__24753));
    Span4Mux_s3_v I__5399 (
            .O(N__24753),
            .I(N__24749));
    InMux I__5398 (
            .O(N__24752),
            .I(N__24746));
    Span4Mux_v I__5397 (
            .O(N__24749),
            .I(N__24741));
    LocalMux I__5396 (
            .O(N__24746),
            .I(N__24738));
    InMux I__5395 (
            .O(N__24745),
            .I(N__24735));
    CascadeMux I__5394 (
            .O(N__24744),
            .I(N__24732));
    Sp12to4 I__5393 (
            .O(N__24741),
            .I(N__24729));
    Span4Mux_h I__5392 (
            .O(N__24738),
            .I(N__24726));
    LocalMux I__5391 (
            .O(N__24735),
            .I(N__24723));
    InMux I__5390 (
            .O(N__24732),
            .I(N__24720));
    Span12Mux_v I__5389 (
            .O(N__24729),
            .I(N__24717));
    Odrv4 I__5388 (
            .O(N__24726),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv4 I__5387 (
            .O(N__24723),
            .I(M_this_sprites_address_qZ0Z_4));
    LocalMux I__5386 (
            .O(N__24720),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv12 I__5385 (
            .O(N__24717),
            .I(M_this_sprites_address_qZ0Z_4));
    InMux I__5384 (
            .O(N__24708),
            .I(N__24705));
    LocalMux I__5383 (
            .O(N__24705),
            .I(N__24702));
    Span4Mux_h I__5382 (
            .O(N__24702),
            .I(N__24699));
    Odrv4 I__5381 (
            .O(N__24699),
            .I(un1_M_this_sprites_address_q_cry_3_THRU_CO));
    InMux I__5380 (
            .O(N__24696),
            .I(un1_M_this_sprites_address_q_cry_3));
    InMux I__5379 (
            .O(N__24693),
            .I(un1_M_this_sprites_address_q_cry_4));
    InMux I__5378 (
            .O(N__24690),
            .I(N__24687));
    LocalMux I__5377 (
            .O(N__24687),
            .I(N__24684));
    Span4Mux_h I__5376 (
            .O(N__24684),
            .I(N__24681));
    Span4Mux_v I__5375 (
            .O(N__24681),
            .I(N__24677));
    InMux I__5374 (
            .O(N__24680),
            .I(N__24674));
    Odrv4 I__5373 (
            .O(N__24677),
            .I(\this_start_data_delay.N_93_0 ));
    LocalMux I__5372 (
            .O(N__24674),
            .I(\this_start_data_delay.N_93_0 ));
    InMux I__5371 (
            .O(N__24669),
            .I(N__24666));
    LocalMux I__5370 (
            .O(N__24666),
            .I(N__24663));
    Span4Mux_v I__5369 (
            .O(N__24663),
            .I(N__24660));
    Span4Mux_v I__5368 (
            .O(N__24660),
            .I(N__24657));
    Odrv4 I__5367 (
            .O(N__24657),
            .I(\this_start_data_delay.N_122 ));
    CascadeMux I__5366 (
            .O(N__24654),
            .I(N__24651));
    InMux I__5365 (
            .O(N__24651),
            .I(N__24648));
    LocalMux I__5364 (
            .O(N__24648),
            .I(N__24644));
    InMux I__5363 (
            .O(N__24647),
            .I(N__24641));
    Odrv12 I__5362 (
            .O(N__24644),
            .I(\this_start_data_delay.N_149 ));
    LocalMux I__5361 (
            .O(N__24641),
            .I(\this_start_data_delay.N_149 ));
    InMux I__5360 (
            .O(N__24636),
            .I(N__24633));
    LocalMux I__5359 (
            .O(N__24633),
            .I(N__24630));
    Span4Mux_v I__5358 (
            .O(N__24630),
            .I(N__24627));
    Odrv4 I__5357 (
            .O(N__24627),
            .I(\this_start_data_delay.N_121 ));
    InMux I__5356 (
            .O(N__24624),
            .I(N__24619));
    InMux I__5355 (
            .O(N__24623),
            .I(N__24616));
    InMux I__5354 (
            .O(N__24622),
            .I(N__24613));
    LocalMux I__5353 (
            .O(N__24619),
            .I(N__24610));
    LocalMux I__5352 (
            .O(N__24616),
            .I(N__24605));
    LocalMux I__5351 (
            .O(N__24613),
            .I(N__24600));
    Span4Mux_h I__5350 (
            .O(N__24610),
            .I(N__24600));
    InMux I__5349 (
            .O(N__24609),
            .I(N__24597));
    InMux I__5348 (
            .O(N__24608),
            .I(N__24594));
    Odrv12 I__5347 (
            .O(N__24605),
            .I(\this_start_data_delay.N_938_0 ));
    Odrv4 I__5346 (
            .O(N__24600),
            .I(\this_start_data_delay.N_938_0 ));
    LocalMux I__5345 (
            .O(N__24597),
            .I(\this_start_data_delay.N_938_0 ));
    LocalMux I__5344 (
            .O(N__24594),
            .I(\this_start_data_delay.N_938_0 ));
    InMux I__5343 (
            .O(N__24585),
            .I(N__24581));
    InMux I__5342 (
            .O(N__24584),
            .I(N__24577));
    LocalMux I__5341 (
            .O(N__24581),
            .I(N__24573));
    InMux I__5340 (
            .O(N__24580),
            .I(N__24570));
    LocalMux I__5339 (
            .O(N__24577),
            .I(N__24566));
    InMux I__5338 (
            .O(N__24576),
            .I(N__24563));
    Span4Mux_v I__5337 (
            .O(N__24573),
            .I(N__24557));
    LocalMux I__5336 (
            .O(N__24570),
            .I(N__24557));
    InMux I__5335 (
            .O(N__24569),
            .I(N__24554));
    Span4Mux_s2_v I__5334 (
            .O(N__24566),
            .I(N__24548));
    LocalMux I__5333 (
            .O(N__24563),
            .I(N__24548));
    InMux I__5332 (
            .O(N__24562),
            .I(N__24545));
    Span4Mux_v I__5331 (
            .O(N__24557),
            .I(N__24541));
    LocalMux I__5330 (
            .O(N__24554),
            .I(N__24538));
    InMux I__5329 (
            .O(N__24553),
            .I(N__24535));
    Span4Mux_v I__5328 (
            .O(N__24548),
            .I(N__24530));
    LocalMux I__5327 (
            .O(N__24545),
            .I(N__24530));
    InMux I__5326 (
            .O(N__24544),
            .I(N__24527));
    Span4Mux_v I__5325 (
            .O(N__24541),
            .I(N__24520));
    Span4Mux_v I__5324 (
            .O(N__24538),
            .I(N__24520));
    LocalMux I__5323 (
            .O(N__24535),
            .I(N__24520));
    Span4Mux_v I__5322 (
            .O(N__24530),
            .I(N__24515));
    LocalMux I__5321 (
            .O(N__24527),
            .I(N__24515));
    Span4Mux_v I__5320 (
            .O(N__24520),
            .I(N__24510));
    Span4Mux_v I__5319 (
            .O(N__24515),
            .I(N__24510));
    Odrv4 I__5318 (
            .O(N__24510),
            .I(N_813_0));
    InMux I__5317 (
            .O(N__24507),
            .I(N__24504));
    LocalMux I__5316 (
            .O(N__24504),
            .I(N__24499));
    InMux I__5315 (
            .O(N__24503),
            .I(N__24494));
    InMux I__5314 (
            .O(N__24502),
            .I(N__24491));
    Span4Mux_v I__5313 (
            .O(N__24499),
            .I(N__24484));
    CascadeMux I__5312 (
            .O(N__24498),
            .I(N__24481));
    CascadeMux I__5311 (
            .O(N__24497),
            .I(N__24478));
    LocalMux I__5310 (
            .O(N__24494),
            .I(N__24475));
    LocalMux I__5309 (
            .O(N__24491),
            .I(N__24470));
    InMux I__5308 (
            .O(N__24490),
            .I(N__24467));
    InMux I__5307 (
            .O(N__24489),
            .I(N__24464));
    InMux I__5306 (
            .O(N__24488),
            .I(N__24459));
    CascadeMux I__5305 (
            .O(N__24487),
            .I(N__24455));
    Span4Mux_h I__5304 (
            .O(N__24484),
            .I(N__24452));
    InMux I__5303 (
            .O(N__24481),
            .I(N__24449));
    InMux I__5302 (
            .O(N__24478),
            .I(N__24446));
    Span4Mux_v I__5301 (
            .O(N__24475),
            .I(N__24442));
    InMux I__5300 (
            .O(N__24474),
            .I(N__24439));
    CascadeMux I__5299 (
            .O(N__24473),
            .I(N__24436));
    Span4Mux_h I__5298 (
            .O(N__24470),
            .I(N__24429));
    LocalMux I__5297 (
            .O(N__24467),
            .I(N__24429));
    LocalMux I__5296 (
            .O(N__24464),
            .I(N__24429));
    InMux I__5295 (
            .O(N__24463),
            .I(N__24426));
    CascadeMux I__5294 (
            .O(N__24462),
            .I(N__24423));
    LocalMux I__5293 (
            .O(N__24459),
            .I(N__24420));
    InMux I__5292 (
            .O(N__24458),
            .I(N__24415));
    InMux I__5291 (
            .O(N__24455),
            .I(N__24415));
    Span4Mux_h I__5290 (
            .O(N__24452),
            .I(N__24412));
    LocalMux I__5289 (
            .O(N__24449),
            .I(N__24409));
    LocalMux I__5288 (
            .O(N__24446),
            .I(N__24406));
    InMux I__5287 (
            .O(N__24445),
            .I(N__24403));
    Span4Mux_v I__5286 (
            .O(N__24442),
            .I(N__24398));
    LocalMux I__5285 (
            .O(N__24439),
            .I(N__24398));
    InMux I__5284 (
            .O(N__24436),
            .I(N__24395));
    Span4Mux_v I__5283 (
            .O(N__24429),
            .I(N__24392));
    LocalMux I__5282 (
            .O(N__24426),
            .I(N__24389));
    InMux I__5281 (
            .O(N__24423),
            .I(N__24386));
    Span4Mux_h I__5280 (
            .O(N__24420),
            .I(N__24381));
    LocalMux I__5279 (
            .O(N__24415),
            .I(N__24381));
    Span4Mux_h I__5278 (
            .O(N__24412),
            .I(N__24372));
    Span4Mux_v I__5277 (
            .O(N__24409),
            .I(N__24372));
    Span4Mux_v I__5276 (
            .O(N__24406),
            .I(N__24372));
    LocalMux I__5275 (
            .O(N__24403),
            .I(N__24372));
    Span4Mux_v I__5274 (
            .O(N__24398),
            .I(N__24367));
    LocalMux I__5273 (
            .O(N__24395),
            .I(N__24367));
    Sp12to4 I__5272 (
            .O(N__24392),
            .I(N__24364));
    Span12Mux_h I__5271 (
            .O(N__24389),
            .I(N__24359));
    LocalMux I__5270 (
            .O(N__24386),
            .I(N__24359));
    Span4Mux_v I__5269 (
            .O(N__24381),
            .I(N__24354));
    Span4Mux_v I__5268 (
            .O(N__24372),
            .I(N__24354));
    Span4Mux_h I__5267 (
            .O(N__24367),
            .I(N__24351));
    Span12Mux_h I__5266 (
            .O(N__24364),
            .I(N__24348));
    Span12Mux_h I__5265 (
            .O(N__24359),
            .I(N__24345));
    Sp12to4 I__5264 (
            .O(N__24354),
            .I(N__24342));
    Span4Mux_h I__5263 (
            .O(N__24351),
            .I(N__24339));
    Odrv12 I__5262 (
            .O(N__24348),
            .I(port_data_c_5));
    Odrv12 I__5261 (
            .O(N__24345),
            .I(port_data_c_5));
    Odrv12 I__5260 (
            .O(N__24342),
            .I(port_data_c_5));
    Odrv4 I__5259 (
            .O(N__24339),
            .I(port_data_c_5));
    CascadeMux I__5258 (
            .O(N__24330),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_6_cascade_ ));
    InMux I__5257 (
            .O(N__24327),
            .I(N__24324));
    LocalMux I__5256 (
            .O(N__24324),
            .I(N__24321));
    Odrv12 I__5255 (
            .O(N__24321),
            .I(\this_start_data_delay.N_68 ));
    CascadeMux I__5254 (
            .O(N__24318),
            .I(N__24314));
    CascadeMux I__5253 (
            .O(N__24317),
            .I(N__24310));
    InMux I__5252 (
            .O(N__24314),
            .I(N__24305));
    CascadeMux I__5251 (
            .O(N__24313),
            .I(N__24302));
    InMux I__5250 (
            .O(N__24310),
            .I(N__24298));
    InMux I__5249 (
            .O(N__24309),
            .I(N__24295));
    InMux I__5248 (
            .O(N__24308),
            .I(N__24292));
    LocalMux I__5247 (
            .O(N__24305),
            .I(N__24289));
    InMux I__5246 (
            .O(N__24302),
            .I(N__24286));
    CascadeMux I__5245 (
            .O(N__24301),
            .I(N__24282));
    LocalMux I__5244 (
            .O(N__24298),
            .I(N__24278));
    LocalMux I__5243 (
            .O(N__24295),
            .I(N__24275));
    LocalMux I__5242 (
            .O(N__24292),
            .I(N__24268));
    Span4Mux_h I__5241 (
            .O(N__24289),
            .I(N__24268));
    LocalMux I__5240 (
            .O(N__24286),
            .I(N__24268));
    InMux I__5239 (
            .O(N__24285),
            .I(N__24265));
    InMux I__5238 (
            .O(N__24282),
            .I(N__24260));
    InMux I__5237 (
            .O(N__24281),
            .I(N__24260));
    Span4Mux_h I__5236 (
            .O(N__24278),
            .I(N__24257));
    Span4Mux_v I__5235 (
            .O(N__24275),
            .I(N__24252));
    Span4Mux_h I__5234 (
            .O(N__24268),
            .I(N__24252));
    LocalMux I__5233 (
            .O(N__24265),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__5232 (
            .O(N__24260),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__5231 (
            .O(N__24257),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__5230 (
            .O(N__24252),
            .I(M_this_state_qZ0Z_5));
    InMux I__5229 (
            .O(N__24243),
            .I(N__24236));
    InMux I__5228 (
            .O(N__24242),
            .I(N__24232));
    InMux I__5227 (
            .O(N__24241),
            .I(N__24228));
    InMux I__5226 (
            .O(N__24240),
            .I(N__24218));
    InMux I__5225 (
            .O(N__24239),
            .I(N__24214));
    LocalMux I__5224 (
            .O(N__24236),
            .I(N__24211));
    InMux I__5223 (
            .O(N__24235),
            .I(N__24208));
    LocalMux I__5222 (
            .O(N__24232),
            .I(N__24205));
    InMux I__5221 (
            .O(N__24231),
            .I(N__24201));
    LocalMux I__5220 (
            .O(N__24228),
            .I(N__24198));
    InMux I__5219 (
            .O(N__24227),
            .I(N__24195));
    InMux I__5218 (
            .O(N__24226),
            .I(N__24192));
    InMux I__5217 (
            .O(N__24225),
            .I(N__24187));
    InMux I__5216 (
            .O(N__24224),
            .I(N__24187));
    InMux I__5215 (
            .O(N__24223),
            .I(N__24180));
    InMux I__5214 (
            .O(N__24222),
            .I(N__24180));
    InMux I__5213 (
            .O(N__24221),
            .I(N__24180));
    LocalMux I__5212 (
            .O(N__24218),
            .I(N__24175));
    InMux I__5211 (
            .O(N__24217),
            .I(N__24172));
    LocalMux I__5210 (
            .O(N__24214),
            .I(N__24165));
    Span4Mux_v I__5209 (
            .O(N__24211),
            .I(N__24165));
    LocalMux I__5208 (
            .O(N__24208),
            .I(N__24165));
    Span4Mux_h I__5207 (
            .O(N__24205),
            .I(N__24154));
    InMux I__5206 (
            .O(N__24204),
            .I(N__24151));
    LocalMux I__5205 (
            .O(N__24201),
            .I(N__24144));
    Span4Mux_h I__5204 (
            .O(N__24198),
            .I(N__24144));
    LocalMux I__5203 (
            .O(N__24195),
            .I(N__24144));
    LocalMux I__5202 (
            .O(N__24192),
            .I(N__24141));
    LocalMux I__5201 (
            .O(N__24187),
            .I(N__24136));
    LocalMux I__5200 (
            .O(N__24180),
            .I(N__24136));
    InMux I__5199 (
            .O(N__24179),
            .I(N__24131));
    InMux I__5198 (
            .O(N__24178),
            .I(N__24131));
    Span4Mux_v I__5197 (
            .O(N__24175),
            .I(N__24118));
    LocalMux I__5196 (
            .O(N__24172),
            .I(N__24118));
    Span4Mux_h I__5195 (
            .O(N__24165),
            .I(N__24118));
    InMux I__5194 (
            .O(N__24164),
            .I(N__24115));
    InMux I__5193 (
            .O(N__24163),
            .I(N__24110));
    InMux I__5192 (
            .O(N__24162),
            .I(N__24110));
    InMux I__5191 (
            .O(N__24161),
            .I(N__24107));
    InMux I__5190 (
            .O(N__24160),
            .I(N__24098));
    InMux I__5189 (
            .O(N__24159),
            .I(N__24098));
    InMux I__5188 (
            .O(N__24158),
            .I(N__24098));
    InMux I__5187 (
            .O(N__24157),
            .I(N__24098));
    Span4Mux_h I__5186 (
            .O(N__24154),
            .I(N__24093));
    LocalMux I__5185 (
            .O(N__24151),
            .I(N__24093));
    Span4Mux_h I__5184 (
            .O(N__24144),
            .I(N__24084));
    Span4Mux_v I__5183 (
            .O(N__24141),
            .I(N__24084));
    Span4Mux_h I__5182 (
            .O(N__24136),
            .I(N__24084));
    LocalMux I__5181 (
            .O(N__24131),
            .I(N__24084));
    InMux I__5180 (
            .O(N__24130),
            .I(N__24077));
    InMux I__5179 (
            .O(N__24129),
            .I(N__24077));
    InMux I__5178 (
            .O(N__24128),
            .I(N__24077));
    InMux I__5177 (
            .O(N__24127),
            .I(N__24070));
    InMux I__5176 (
            .O(N__24126),
            .I(N__24070));
    InMux I__5175 (
            .O(N__24125),
            .I(N__24070));
    Odrv4 I__5174 (
            .O(N__24118),
            .I(N_554_0));
    LocalMux I__5173 (
            .O(N__24115),
            .I(N_554_0));
    LocalMux I__5172 (
            .O(N__24110),
            .I(N_554_0));
    LocalMux I__5171 (
            .O(N__24107),
            .I(N_554_0));
    LocalMux I__5170 (
            .O(N__24098),
            .I(N_554_0));
    Odrv4 I__5169 (
            .O(N__24093),
            .I(N_554_0));
    Odrv4 I__5168 (
            .O(N__24084),
            .I(N_554_0));
    LocalMux I__5167 (
            .O(N__24077),
            .I(N_554_0));
    LocalMux I__5166 (
            .O(N__24070),
            .I(N_554_0));
    CascadeMux I__5165 (
            .O(N__24051),
            .I(this_start_data_delay_M_this_data_count_q_3_0_a3_0_6_cascade_));
    InMux I__5164 (
            .O(N__24048),
            .I(N__24029));
    InMux I__5163 (
            .O(N__24047),
            .I(N__24029));
    InMux I__5162 (
            .O(N__24046),
            .I(N__24029));
    InMux I__5161 (
            .O(N__24045),
            .I(N__24029));
    InMux I__5160 (
            .O(N__24044),
            .I(N__24020));
    InMux I__5159 (
            .O(N__24043),
            .I(N__24020));
    InMux I__5158 (
            .O(N__24042),
            .I(N__24020));
    InMux I__5157 (
            .O(N__24041),
            .I(N__24020));
    InMux I__5156 (
            .O(N__24040),
            .I(N__24016));
    InMux I__5155 (
            .O(N__24039),
            .I(N__24011));
    InMux I__5154 (
            .O(N__24038),
            .I(N__24011));
    LocalMux I__5153 (
            .O(N__24029),
            .I(N__24006));
    LocalMux I__5152 (
            .O(N__24020),
            .I(N__24006));
    InMux I__5151 (
            .O(N__24019),
            .I(N__24003));
    LocalMux I__5150 (
            .O(N__24016),
            .I(N__24000));
    LocalMux I__5149 (
            .O(N__24011),
            .I(N__23994));
    Span12Mux_v I__5148 (
            .O(N__24006),
            .I(N__23994));
    LocalMux I__5147 (
            .O(N__24003),
            .I(N__23991));
    Span4Mux_v I__5146 (
            .O(N__24000),
            .I(N__23988));
    InMux I__5145 (
            .O(N__23999),
            .I(N__23985));
    Span12Mux_h I__5144 (
            .O(N__23994),
            .I(N__23982));
    Span4Mux_h I__5143 (
            .O(N__23991),
            .I(N__23979));
    Odrv4 I__5142 (
            .O(N__23988),
            .I(N_911));
    LocalMux I__5141 (
            .O(N__23985),
            .I(N_911));
    Odrv12 I__5140 (
            .O(N__23982),
            .I(N_911));
    Odrv4 I__5139 (
            .O(N__23979),
            .I(N_911));
    InMux I__5138 (
            .O(N__23970),
            .I(N__23967));
    LocalMux I__5137 (
            .O(N__23967),
            .I(N__23964));
    Span4Mux_h I__5136 (
            .O(N__23964),
            .I(N__23961));
    Odrv4 I__5135 (
            .O(N__23961),
            .I(M_this_data_count_q_3_0_13));
    InMux I__5134 (
            .O(N__23958),
            .I(N__23951));
    InMux I__5133 (
            .O(N__23957),
            .I(N__23948));
    InMux I__5132 (
            .O(N__23956),
            .I(N__23942));
    InMux I__5131 (
            .O(N__23955),
            .I(N__23942));
    InMux I__5130 (
            .O(N__23954),
            .I(N__23939));
    LocalMux I__5129 (
            .O(N__23951),
            .I(N__23936));
    LocalMux I__5128 (
            .O(N__23948),
            .I(N__23933));
    InMux I__5127 (
            .O(N__23947),
            .I(N__23930));
    LocalMux I__5126 (
            .O(N__23942),
            .I(N__23927));
    LocalMux I__5125 (
            .O(N__23939),
            .I(N__23922));
    Span4Mux_h I__5124 (
            .O(N__23936),
            .I(N__23922));
    Odrv4 I__5123 (
            .O(N__23933),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__5122 (
            .O(N__23930),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__5121 (
            .O(N__23927),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__5120 (
            .O(N__23922),
            .I(M_this_state_qZ0Z_9));
    InMux I__5119 (
            .O(N__23913),
            .I(N__23910));
    LocalMux I__5118 (
            .O(N__23910),
            .I(N__23907));
    Span4Mux_h I__5117 (
            .O(N__23907),
            .I(N__23902));
    InMux I__5116 (
            .O(N__23906),
            .I(N__23896));
    InMux I__5115 (
            .O(N__23905),
            .I(N__23896));
    Span4Mux_h I__5114 (
            .O(N__23902),
            .I(N__23893));
    InMux I__5113 (
            .O(N__23901),
            .I(N__23890));
    LocalMux I__5112 (
            .O(N__23896),
            .I(N__23886));
    Sp12to4 I__5111 (
            .O(N__23893),
            .I(N__23881));
    LocalMux I__5110 (
            .O(N__23890),
            .I(N__23881));
    InMux I__5109 (
            .O(N__23889),
            .I(N__23878));
    Span4Mux_v I__5108 (
            .O(N__23886),
            .I(N__23875));
    Odrv12 I__5107 (
            .O(N__23881),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__5106 (
            .O(N__23878),
            .I(M_this_state_qZ0Z_7));
    Odrv4 I__5105 (
            .O(N__23875),
            .I(M_this_state_qZ0Z_7));
    CascadeMux I__5104 (
            .O(N__23868),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_3_cascade_ ));
    CascadeMux I__5103 (
            .O(N__23865),
            .I(N__23862));
    InMux I__5102 (
            .O(N__23862),
            .I(N__23859));
    LocalMux I__5101 (
            .O(N__23859),
            .I(N__23856));
    Span4Mux_h I__5100 (
            .O(N__23856),
            .I(N__23853));
    Sp12to4 I__5099 (
            .O(N__23853),
            .I(N__23850));
    Span12Mux_v I__5098 (
            .O(N__23850),
            .I(N__23847));
    Span12Mux_h I__5097 (
            .O(N__23847),
            .I(N__23844));
    Odrv12 I__5096 (
            .O(N__23844),
            .I(M_this_map_ram_read_data_7));
    InMux I__5095 (
            .O(N__23841),
            .I(N__23838));
    LocalMux I__5094 (
            .O(N__23838),
            .I(N__23835));
    Odrv12 I__5093 (
            .O(N__23835),
            .I(\this_ppu.un10_sprites_addr_cry_4_c_RNIUV9BZ0 ));
    InMux I__5092 (
            .O(N__23832),
            .I(N__23829));
    LocalMux I__5091 (
            .O(N__23829),
            .I(N__23824));
    InMux I__5090 (
            .O(N__23828),
            .I(N__23821));
    InMux I__5089 (
            .O(N__23827),
            .I(N__23817));
    Span4Mux_v I__5088 (
            .O(N__23824),
            .I(N__23812));
    LocalMux I__5087 (
            .O(N__23821),
            .I(N__23812));
    InMux I__5086 (
            .O(N__23820),
            .I(N__23809));
    LocalMux I__5085 (
            .O(N__23817),
            .I(\this_start_data_delay.N_91_0 ));
    Odrv4 I__5084 (
            .O(N__23812),
            .I(\this_start_data_delay.N_91_0 ));
    LocalMux I__5083 (
            .O(N__23809),
            .I(\this_start_data_delay.N_91_0 ));
    CascadeMux I__5082 (
            .O(N__23802),
            .I(\this_start_data_delay.N_149_cascade_ ));
    InMux I__5081 (
            .O(N__23799),
            .I(N__23792));
    CascadeMux I__5080 (
            .O(N__23798),
            .I(N__23788));
    InMux I__5079 (
            .O(N__23797),
            .I(N__23785));
    InMux I__5078 (
            .O(N__23796),
            .I(N__23782));
    CascadeMux I__5077 (
            .O(N__23795),
            .I(N__23777));
    LocalMux I__5076 (
            .O(N__23792),
            .I(N__23773));
    InMux I__5075 (
            .O(N__23791),
            .I(N__23770));
    InMux I__5074 (
            .O(N__23788),
            .I(N__23767));
    LocalMux I__5073 (
            .O(N__23785),
            .I(N__23762));
    LocalMux I__5072 (
            .O(N__23782),
            .I(N__23762));
    InMux I__5071 (
            .O(N__23781),
            .I(N__23757));
    InMux I__5070 (
            .O(N__23780),
            .I(N__23757));
    InMux I__5069 (
            .O(N__23777),
            .I(N__23752));
    InMux I__5068 (
            .O(N__23776),
            .I(N__23752));
    Span4Mux_v I__5067 (
            .O(N__23773),
            .I(N__23745));
    LocalMux I__5066 (
            .O(N__23770),
            .I(N__23745));
    LocalMux I__5065 (
            .O(N__23767),
            .I(N__23745));
    Span4Mux_v I__5064 (
            .O(N__23762),
            .I(N__23740));
    LocalMux I__5063 (
            .O(N__23757),
            .I(N__23740));
    LocalMux I__5062 (
            .O(N__23752),
            .I(M_this_state_qZ0Z_6));
    Odrv4 I__5061 (
            .O(N__23745),
            .I(M_this_state_qZ0Z_6));
    Odrv4 I__5060 (
            .O(N__23740),
            .I(M_this_state_qZ0Z_6));
    InMux I__5059 (
            .O(N__23733),
            .I(N__23728));
    InMux I__5058 (
            .O(N__23732),
            .I(N__23723));
    InMux I__5057 (
            .O(N__23731),
            .I(N__23720));
    LocalMux I__5056 (
            .O(N__23728),
            .I(N__23717));
    InMux I__5055 (
            .O(N__23727),
            .I(N__23714));
    InMux I__5054 (
            .O(N__23726),
            .I(N__23711));
    LocalMux I__5053 (
            .O(N__23723),
            .I(N__23708));
    LocalMux I__5052 (
            .O(N__23720),
            .I(N__23703));
    Span4Mux_h I__5051 (
            .O(N__23717),
            .I(N__23703));
    LocalMux I__5050 (
            .O(N__23714),
            .I(\this_start_data_delay.N_555_0 ));
    LocalMux I__5049 (
            .O(N__23711),
            .I(\this_start_data_delay.N_555_0 ));
    Odrv4 I__5048 (
            .O(N__23708),
            .I(\this_start_data_delay.N_555_0 ));
    Odrv4 I__5047 (
            .O(N__23703),
            .I(\this_start_data_delay.N_555_0 ));
    InMux I__5046 (
            .O(N__23694),
            .I(N__23691));
    LocalMux I__5045 (
            .O(N__23691),
            .I(N__23688));
    Odrv4 I__5044 (
            .O(N__23688),
            .I(\this_start_data_delay.M_this_data_count_qlde_i_a3_0 ));
    InMux I__5043 (
            .O(N__23685),
            .I(N__23682));
    LocalMux I__5042 (
            .O(N__23682),
            .I(\this_start_data_delay.M_this_data_count_qlde_i_2_tz_0 ));
    CascadeMux I__5041 (
            .O(N__23679),
            .I(\this_start_data_delay.N_820_0_cascade_ ));
    InMux I__5040 (
            .O(N__23676),
            .I(N__23673));
    LocalMux I__5039 (
            .O(N__23673),
            .I(N__23670));
    Span4Mux_h I__5038 (
            .O(N__23670),
            .I(N__23667));
    Odrv4 I__5037 (
            .O(N__23667),
            .I(\this_start_data_delay.N_151 ));
    InMux I__5036 (
            .O(N__23664),
            .I(N__23660));
    InMux I__5035 (
            .O(N__23663),
            .I(N__23657));
    LocalMux I__5034 (
            .O(N__23660),
            .I(N__23653));
    LocalMux I__5033 (
            .O(N__23657),
            .I(N__23649));
    InMux I__5032 (
            .O(N__23656),
            .I(N__23646));
    Span4Mux_h I__5031 (
            .O(N__23653),
            .I(N__23643));
    InMux I__5030 (
            .O(N__23652),
            .I(N__23640));
    Span4Mux_v I__5029 (
            .O(N__23649),
            .I(N__23637));
    LocalMux I__5028 (
            .O(N__23646),
            .I(\this_start_data_delay.N_820_0 ));
    Odrv4 I__5027 (
            .O(N__23643),
            .I(\this_start_data_delay.N_820_0 ));
    LocalMux I__5026 (
            .O(N__23640),
            .I(\this_start_data_delay.N_820_0 ));
    Odrv4 I__5025 (
            .O(N__23637),
            .I(\this_start_data_delay.N_820_0 ));
    CascadeMux I__5024 (
            .O(N__23628),
            .I(\this_start_data_delay.M_this_data_count_qlde_i_1_cascade_ ));
    InMux I__5023 (
            .O(N__23625),
            .I(N__23622));
    LocalMux I__5022 (
            .O(N__23622),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_11 ));
    CascadeMux I__5021 (
            .O(N__23619),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_10_cascade_ ));
    InMux I__5020 (
            .O(N__23616),
            .I(N__23613));
    LocalMux I__5019 (
            .O(N__23613),
            .I(N__23610));
    Span4Mux_v I__5018 (
            .O(N__23610),
            .I(N__23607));
    Span4Mux_v I__5017 (
            .O(N__23607),
            .I(N__23604));
    Span4Mux_h I__5016 (
            .O(N__23604),
            .I(N__23601));
    Odrv4 I__5015 (
            .O(N__23601),
            .I(\this_sprites_ram.mem_out_bus7_1 ));
    InMux I__5014 (
            .O(N__23598),
            .I(N__23595));
    LocalMux I__5013 (
            .O(N__23595),
            .I(N__23592));
    Span4Mux_v I__5012 (
            .O(N__23592),
            .I(N__23589));
    Span4Mux_h I__5011 (
            .O(N__23589),
            .I(N__23586));
    Odrv4 I__5010 (
            .O(N__23586),
            .I(\this_sprites_ram.mem_out_bus3_1 ));
    InMux I__5009 (
            .O(N__23583),
            .I(N__23580));
    LocalMux I__5008 (
            .O(N__23580),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ));
    CascadeMux I__5007 (
            .O(N__23577),
            .I(N__23573));
    InMux I__5006 (
            .O(N__23576),
            .I(N__23568));
    InMux I__5005 (
            .O(N__23573),
            .I(N__23565));
    CascadeMux I__5004 (
            .O(N__23572),
            .I(N__23562));
    InMux I__5003 (
            .O(N__23571),
            .I(N__23559));
    LocalMux I__5002 (
            .O(N__23568),
            .I(N__23556));
    LocalMux I__5001 (
            .O(N__23565),
            .I(N__23553));
    InMux I__5000 (
            .O(N__23562),
            .I(N__23550));
    LocalMux I__4999 (
            .O(N__23559),
            .I(N__23547));
    Span4Mux_v I__4998 (
            .O(N__23556),
            .I(N__23542));
    Span4Mux_v I__4997 (
            .O(N__23553),
            .I(N__23542));
    LocalMux I__4996 (
            .O(N__23550),
            .I(N__23539));
    Odrv4 I__4995 (
            .O(N__23547),
            .I(\this_start_data_delay.N_55_0 ));
    Odrv4 I__4994 (
            .O(N__23542),
            .I(\this_start_data_delay.N_55_0 ));
    Odrv4 I__4993 (
            .O(N__23539),
            .I(\this_start_data_delay.N_55_0 ));
    InMux I__4992 (
            .O(N__23532),
            .I(N__23528));
    InMux I__4991 (
            .O(N__23531),
            .I(N__23525));
    LocalMux I__4990 (
            .O(N__23528),
            .I(N__23522));
    LocalMux I__4989 (
            .O(N__23525),
            .I(N__23519));
    Odrv4 I__4988 (
            .O(N__23522),
            .I(\this_start_data_delay.N_84 ));
    Odrv4 I__4987 (
            .O(N__23519),
            .I(\this_start_data_delay.N_84 ));
    CascadeMux I__4986 (
            .O(N__23514),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_2_cascade_ ));
    CascadeMux I__4985 (
            .O(N__23511),
            .I(\this_start_data_delay.N_913_cascade_ ));
    InMux I__4984 (
            .O(N__23508),
            .I(N__23505));
    LocalMux I__4983 (
            .O(N__23505),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_7 ));
    CascadeMux I__4982 (
            .O(N__23502),
            .I(\this_start_data_delay.N_129_cascade_ ));
    CascadeMux I__4981 (
            .O(N__23499),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_12_cascade_ ));
    CascadeMux I__4980 (
            .O(N__23496),
            .I(N__23492));
    CascadeMux I__4979 (
            .O(N__23495),
            .I(N__23486));
    InMux I__4978 (
            .O(N__23492),
            .I(N__23483));
    InMux I__4977 (
            .O(N__23491),
            .I(N__23478));
    InMux I__4976 (
            .O(N__23490),
            .I(N__23478));
    InMux I__4975 (
            .O(N__23489),
            .I(N__23475));
    InMux I__4974 (
            .O(N__23486),
            .I(N__23469));
    LocalMux I__4973 (
            .O(N__23483),
            .I(N__23464));
    LocalMux I__4972 (
            .O(N__23478),
            .I(N__23464));
    LocalMux I__4971 (
            .O(N__23475),
            .I(N__23461));
    InMux I__4970 (
            .O(N__23474),
            .I(N__23458));
    InMux I__4969 (
            .O(N__23473),
            .I(N__23455));
    InMux I__4968 (
            .O(N__23472),
            .I(N__23452));
    LocalMux I__4967 (
            .O(N__23469),
            .I(N__23447));
    Span4Mux_h I__4966 (
            .O(N__23464),
            .I(N__23447));
    Odrv4 I__4965 (
            .O(N__23461),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__4964 (
            .O(N__23458),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__4963 (
            .O(N__23455),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__4962 (
            .O(N__23452),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__4961 (
            .O(N__23447),
            .I(M_this_state_qZ0Z_8));
    CascadeMux I__4960 (
            .O(N__23436),
            .I(\this_start_data_delay.N_821_0_cascade_ ));
    InMux I__4959 (
            .O(N__23433),
            .I(N__23430));
    LocalMux I__4958 (
            .O(N__23430),
            .I(N__23425));
    InMux I__4957 (
            .O(N__23429),
            .I(N__23420));
    InMux I__4956 (
            .O(N__23428),
            .I(N__23420));
    Odrv4 I__4955 (
            .O(N__23425),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    LocalMux I__4954 (
            .O(N__23420),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    InMux I__4953 (
            .O(N__23415),
            .I(N__23412));
    LocalMux I__4952 (
            .O(N__23412),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    CEMux I__4951 (
            .O(N__23409),
            .I(N__23403));
    CEMux I__4950 (
            .O(N__23408),
            .I(N__23398));
    CEMux I__4949 (
            .O(N__23407),
            .I(N__23394));
    CEMux I__4948 (
            .O(N__23406),
            .I(N__23391));
    LocalMux I__4947 (
            .O(N__23403),
            .I(N__23388));
    CEMux I__4946 (
            .O(N__23402),
            .I(N__23385));
    CEMux I__4945 (
            .O(N__23401),
            .I(N__23382));
    LocalMux I__4944 (
            .O(N__23398),
            .I(N__23379));
    CEMux I__4943 (
            .O(N__23397),
            .I(N__23376));
    LocalMux I__4942 (
            .O(N__23394),
            .I(N__23373));
    LocalMux I__4941 (
            .O(N__23391),
            .I(N__23370));
    Span4Mux_h I__4940 (
            .O(N__23388),
            .I(N__23367));
    LocalMux I__4939 (
            .O(N__23385),
            .I(N__23364));
    LocalMux I__4938 (
            .O(N__23382),
            .I(N__23361));
    Span4Mux_h I__4937 (
            .O(N__23379),
            .I(N__23355));
    LocalMux I__4936 (
            .O(N__23376),
            .I(N__23355));
    Span4Mux_h I__4935 (
            .O(N__23373),
            .I(N__23352));
    Span4Mux_v I__4934 (
            .O(N__23370),
            .I(N__23349));
    Span4Mux_v I__4933 (
            .O(N__23367),
            .I(N__23342));
    Span4Mux_h I__4932 (
            .O(N__23364),
            .I(N__23342));
    Span4Mux_h I__4931 (
            .O(N__23361),
            .I(N__23342));
    CEMux I__4930 (
            .O(N__23360),
            .I(N__23339));
    Span4Mux_h I__4929 (
            .O(N__23355),
            .I(N__23336));
    Span4Mux_h I__4928 (
            .O(N__23352),
            .I(N__23333));
    Sp12to4 I__4927 (
            .O(N__23349),
            .I(N__23326));
    Sp12to4 I__4926 (
            .O(N__23342),
            .I(N__23326));
    LocalMux I__4925 (
            .O(N__23339),
            .I(N__23326));
    Odrv4 I__4924 (
            .O(N__23336),
            .I(\this_vga_signals.N_1090_0 ));
    Odrv4 I__4923 (
            .O(N__23333),
            .I(\this_vga_signals.N_1090_0 ));
    Odrv12 I__4922 (
            .O(N__23326),
            .I(\this_vga_signals.N_1090_0 ));
    SRMux I__4921 (
            .O(N__23319),
            .I(N__23292));
    SRMux I__4920 (
            .O(N__23318),
            .I(N__23292));
    SRMux I__4919 (
            .O(N__23317),
            .I(N__23292));
    SRMux I__4918 (
            .O(N__23316),
            .I(N__23292));
    SRMux I__4917 (
            .O(N__23315),
            .I(N__23292));
    SRMux I__4916 (
            .O(N__23314),
            .I(N__23292));
    SRMux I__4915 (
            .O(N__23313),
            .I(N__23292));
    SRMux I__4914 (
            .O(N__23312),
            .I(N__23292));
    SRMux I__4913 (
            .O(N__23311),
            .I(N__23292));
    GlobalMux I__4912 (
            .O(N__23292),
            .I(N__23289));
    gio2CtrlBuf I__4911 (
            .O(N__23289),
            .I(\this_vga_signals.N_1358_g ));
    CascadeMux I__4910 (
            .O(N__23286),
            .I(N__23279));
    InMux I__4909 (
            .O(N__23285),
            .I(N__23273));
    CascadeMux I__4908 (
            .O(N__23284),
            .I(N__23269));
    CascadeMux I__4907 (
            .O(N__23283),
            .I(N__23263));
    CascadeMux I__4906 (
            .O(N__23282),
            .I(N__23260));
    InMux I__4905 (
            .O(N__23279),
            .I(N__23254));
    InMux I__4904 (
            .O(N__23278),
            .I(N__23254));
    CascadeMux I__4903 (
            .O(N__23277),
            .I(N__23251));
    InMux I__4902 (
            .O(N__23276),
            .I(N__23245));
    LocalMux I__4901 (
            .O(N__23273),
            .I(N__23242));
    InMux I__4900 (
            .O(N__23272),
            .I(N__23237));
    InMux I__4899 (
            .O(N__23269),
            .I(N__23237));
    InMux I__4898 (
            .O(N__23268),
            .I(N__23234));
    InMux I__4897 (
            .O(N__23267),
            .I(N__23229));
    InMux I__4896 (
            .O(N__23266),
            .I(N__23229));
    InMux I__4895 (
            .O(N__23263),
            .I(N__23222));
    InMux I__4894 (
            .O(N__23260),
            .I(N__23222));
    InMux I__4893 (
            .O(N__23259),
            .I(N__23222));
    LocalMux I__4892 (
            .O(N__23254),
            .I(N__23218));
    InMux I__4891 (
            .O(N__23251),
            .I(N__23215));
    CascadeMux I__4890 (
            .O(N__23250),
            .I(N__23210));
    CascadeMux I__4889 (
            .O(N__23249),
            .I(N__23207));
    InMux I__4888 (
            .O(N__23248),
            .I(N__23204));
    LocalMux I__4887 (
            .O(N__23245),
            .I(N__23194));
    Span4Mux_v I__4886 (
            .O(N__23242),
            .I(N__23194));
    LocalMux I__4885 (
            .O(N__23237),
            .I(N__23191));
    LocalMux I__4884 (
            .O(N__23234),
            .I(N__23184));
    LocalMux I__4883 (
            .O(N__23229),
            .I(N__23184));
    LocalMux I__4882 (
            .O(N__23222),
            .I(N__23184));
    InMux I__4881 (
            .O(N__23221),
            .I(N__23180));
    Span4Mux_v I__4880 (
            .O(N__23218),
            .I(N__23175));
    LocalMux I__4879 (
            .O(N__23215),
            .I(N__23175));
    InMux I__4878 (
            .O(N__23214),
            .I(N__23166));
    InMux I__4877 (
            .O(N__23213),
            .I(N__23166));
    InMux I__4876 (
            .O(N__23210),
            .I(N__23166));
    InMux I__4875 (
            .O(N__23207),
            .I(N__23166));
    LocalMux I__4874 (
            .O(N__23204),
            .I(N__23163));
    CascadeMux I__4873 (
            .O(N__23203),
            .I(N__23160));
    InMux I__4872 (
            .O(N__23202),
            .I(N__23155));
    InMux I__4871 (
            .O(N__23201),
            .I(N__23152));
    InMux I__4870 (
            .O(N__23200),
            .I(N__23147));
    InMux I__4869 (
            .O(N__23199),
            .I(N__23147));
    Span4Mux_v I__4868 (
            .O(N__23194),
            .I(N__23140));
    Span4Mux_v I__4867 (
            .O(N__23191),
            .I(N__23140));
    Span4Mux_v I__4866 (
            .O(N__23184),
            .I(N__23140));
    InMux I__4865 (
            .O(N__23183),
            .I(N__23137));
    LocalMux I__4864 (
            .O(N__23180),
            .I(N__23134));
    Span4Mux_h I__4863 (
            .O(N__23175),
            .I(N__23127));
    LocalMux I__4862 (
            .O(N__23166),
            .I(N__23127));
    Span4Mux_h I__4861 (
            .O(N__23163),
            .I(N__23127));
    InMux I__4860 (
            .O(N__23160),
            .I(N__23120));
    InMux I__4859 (
            .O(N__23159),
            .I(N__23120));
    InMux I__4858 (
            .O(N__23158),
            .I(N__23120));
    LocalMux I__4857 (
            .O(N__23155),
            .I(N__23115));
    LocalMux I__4856 (
            .O(N__23152),
            .I(N__23115));
    LocalMux I__4855 (
            .O(N__23147),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__4854 (
            .O(N__23140),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__4853 (
            .O(N__23137),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv12 I__4852 (
            .O(N__23134),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__4851 (
            .O(N__23127),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__4850 (
            .O(N__23120),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__4849 (
            .O(N__23115),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    CascadeMux I__4848 (
            .O(N__23100),
            .I(N__23094));
    CascadeMux I__4847 (
            .O(N__23099),
            .I(N__23084));
    CascadeMux I__4846 (
            .O(N__23098),
            .I(N__23081));
    CascadeMux I__4845 (
            .O(N__23097),
            .I(N__23078));
    InMux I__4844 (
            .O(N__23094),
            .I(N__23074));
    CascadeMux I__4843 (
            .O(N__23093),
            .I(N__23070));
    CascadeMux I__4842 (
            .O(N__23092),
            .I(N__23066));
    InMux I__4841 (
            .O(N__23091),
            .I(N__23060));
    InMux I__4840 (
            .O(N__23090),
            .I(N__23060));
    InMux I__4839 (
            .O(N__23089),
            .I(N__23057));
    InMux I__4838 (
            .O(N__23088),
            .I(N__23054));
    InMux I__4837 (
            .O(N__23087),
            .I(N__23051));
    InMux I__4836 (
            .O(N__23084),
            .I(N__23048));
    InMux I__4835 (
            .O(N__23081),
            .I(N__23045));
    InMux I__4834 (
            .O(N__23078),
            .I(N__23040));
    InMux I__4833 (
            .O(N__23077),
            .I(N__23040));
    LocalMux I__4832 (
            .O(N__23074),
            .I(N__23036));
    InMux I__4831 (
            .O(N__23073),
            .I(N__23031));
    InMux I__4830 (
            .O(N__23070),
            .I(N__23031));
    InMux I__4829 (
            .O(N__23069),
            .I(N__23026));
    InMux I__4828 (
            .O(N__23066),
            .I(N__23026));
    InMux I__4827 (
            .O(N__23065),
            .I(N__23023));
    LocalMux I__4826 (
            .O(N__23060),
            .I(N__23020));
    LocalMux I__4825 (
            .O(N__23057),
            .I(N__23017));
    LocalMux I__4824 (
            .O(N__23054),
            .I(N__23014));
    LocalMux I__4823 (
            .O(N__23051),
            .I(N__23011));
    LocalMux I__4822 (
            .O(N__23048),
            .I(N__23004));
    LocalMux I__4821 (
            .O(N__23045),
            .I(N__23004));
    LocalMux I__4820 (
            .O(N__23040),
            .I(N__23004));
    CascadeMux I__4819 (
            .O(N__23039),
            .I(N__23001));
    Span4Mux_v I__4818 (
            .O(N__23036),
            .I(N__22991));
    LocalMux I__4817 (
            .O(N__23031),
            .I(N__22988));
    LocalMux I__4816 (
            .O(N__23026),
            .I(N__22983));
    LocalMux I__4815 (
            .O(N__23023),
            .I(N__22983));
    Span4Mux_h I__4814 (
            .O(N__23020),
            .I(N__22980));
    Span4Mux_v I__4813 (
            .O(N__23017),
            .I(N__22971));
    Span4Mux_v I__4812 (
            .O(N__23014),
            .I(N__22971));
    Span4Mux_h I__4811 (
            .O(N__23011),
            .I(N__22971));
    Span4Mux_v I__4810 (
            .O(N__23004),
            .I(N__22971));
    InMux I__4809 (
            .O(N__23001),
            .I(N__22966));
    InMux I__4808 (
            .O(N__23000),
            .I(N__22966));
    InMux I__4807 (
            .O(N__22999),
            .I(N__22957));
    InMux I__4806 (
            .O(N__22998),
            .I(N__22957));
    InMux I__4805 (
            .O(N__22997),
            .I(N__22957));
    InMux I__4804 (
            .O(N__22996),
            .I(N__22957));
    InMux I__4803 (
            .O(N__22995),
            .I(N__22952));
    InMux I__4802 (
            .O(N__22994),
            .I(N__22952));
    Odrv4 I__4801 (
            .O(N__22991),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__4800 (
            .O(N__22988),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__4799 (
            .O(N__22983),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__4798 (
            .O(N__22980),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__4797 (
            .O(N__22971),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__4796 (
            .O(N__22966),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__4795 (
            .O(N__22957),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__4794 (
            .O(N__22952),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    InMux I__4793 (
            .O(N__22935),
            .I(N__22930));
    InMux I__4792 (
            .O(N__22934),
            .I(N__22925));
    InMux I__4791 (
            .O(N__22933),
            .I(N__22922));
    LocalMux I__4790 (
            .O(N__22930),
            .I(N__22919));
    InMux I__4789 (
            .O(N__22929),
            .I(N__22916));
    InMux I__4788 (
            .O(N__22928),
            .I(N__22912));
    LocalMux I__4787 (
            .O(N__22925),
            .I(N__22907));
    LocalMux I__4786 (
            .O(N__22922),
            .I(N__22907));
    Span4Mux_v I__4785 (
            .O(N__22919),
            .I(N__22902));
    LocalMux I__4784 (
            .O(N__22916),
            .I(N__22902));
    InMux I__4783 (
            .O(N__22915),
            .I(N__22899));
    LocalMux I__4782 (
            .O(N__22912),
            .I(N__22895));
    Span4Mux_v I__4781 (
            .O(N__22907),
            .I(N__22890));
    Span4Mux_h I__4780 (
            .O(N__22902),
            .I(N__22890));
    LocalMux I__4779 (
            .O(N__22899),
            .I(N__22887));
    InMux I__4778 (
            .O(N__22898),
            .I(N__22884));
    Span12Mux_h I__4777 (
            .O(N__22895),
            .I(N__22881));
    Span4Mux_h I__4776 (
            .O(N__22890),
            .I(N__22878));
    Odrv12 I__4775 (
            .O(N__22887),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__4774 (
            .O(N__22884),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv12 I__4773 (
            .O(N__22881),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__4772 (
            .O(N__22878),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    CascadeMux I__4771 (
            .O(N__22869),
            .I(N__22862));
    CascadeMux I__4770 (
            .O(N__22868),
            .I(N__22851));
    InMux I__4769 (
            .O(N__22867),
            .I(N__22844));
    InMux I__4768 (
            .O(N__22866),
            .I(N__22844));
    CascadeMux I__4767 (
            .O(N__22865),
            .I(N__22836));
    InMux I__4766 (
            .O(N__22862),
            .I(N__22833));
    InMux I__4765 (
            .O(N__22861),
            .I(N__22830));
    CascadeMux I__4764 (
            .O(N__22860),
            .I(N__22827));
    InMux I__4763 (
            .O(N__22859),
            .I(N__22824));
    InMux I__4762 (
            .O(N__22858),
            .I(N__22821));
    InMux I__4761 (
            .O(N__22857),
            .I(N__22816));
    InMux I__4760 (
            .O(N__22856),
            .I(N__22816));
    InMux I__4759 (
            .O(N__22855),
            .I(N__22813));
    InMux I__4758 (
            .O(N__22854),
            .I(N__22808));
    InMux I__4757 (
            .O(N__22851),
            .I(N__22808));
    InMux I__4756 (
            .O(N__22850),
            .I(N__22803));
    InMux I__4755 (
            .O(N__22849),
            .I(N__22803));
    LocalMux I__4754 (
            .O(N__22844),
            .I(N__22800));
    InMux I__4753 (
            .O(N__22843),
            .I(N__22797));
    InMux I__4752 (
            .O(N__22842),
            .I(N__22794));
    InMux I__4751 (
            .O(N__22841),
            .I(N__22791));
    InMux I__4750 (
            .O(N__22840),
            .I(N__22788));
    InMux I__4749 (
            .O(N__22839),
            .I(N__22783));
    InMux I__4748 (
            .O(N__22836),
            .I(N__22783));
    LocalMux I__4747 (
            .O(N__22833),
            .I(N__22778));
    LocalMux I__4746 (
            .O(N__22830),
            .I(N__22778));
    InMux I__4745 (
            .O(N__22827),
            .I(N__22775));
    LocalMux I__4744 (
            .O(N__22824),
            .I(N__22772));
    LocalMux I__4743 (
            .O(N__22821),
            .I(N__22760));
    LocalMux I__4742 (
            .O(N__22816),
            .I(N__22760));
    LocalMux I__4741 (
            .O(N__22813),
            .I(N__22760));
    LocalMux I__4740 (
            .O(N__22808),
            .I(N__22760));
    LocalMux I__4739 (
            .O(N__22803),
            .I(N__22760));
    Span4Mux_h I__4738 (
            .O(N__22800),
            .I(N__22755));
    LocalMux I__4737 (
            .O(N__22797),
            .I(N__22755));
    LocalMux I__4736 (
            .O(N__22794),
            .I(N__22750));
    LocalMux I__4735 (
            .O(N__22791),
            .I(N__22750));
    LocalMux I__4734 (
            .O(N__22788),
            .I(N__22739));
    LocalMux I__4733 (
            .O(N__22783),
            .I(N__22739));
    Span4Mux_v I__4732 (
            .O(N__22778),
            .I(N__22739));
    LocalMux I__4731 (
            .O(N__22775),
            .I(N__22739));
    Span4Mux_h I__4730 (
            .O(N__22772),
            .I(N__22739));
    InMux I__4729 (
            .O(N__22771),
            .I(N__22736));
    Span4Mux_v I__4728 (
            .O(N__22760),
            .I(N__22733));
    Span4Mux_v I__4727 (
            .O(N__22755),
            .I(N__22730));
    Span4Mux_v I__4726 (
            .O(N__22750),
            .I(N__22725));
    Span4Mux_h I__4725 (
            .O(N__22739),
            .I(N__22725));
    LocalMux I__4724 (
            .O(N__22736),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__4723 (
            .O(N__22733),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__4722 (
            .O(N__22730),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__4721 (
            .O(N__22725),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    CascadeMux I__4720 (
            .O(N__22716),
            .I(N__22710));
    InMux I__4719 (
            .O(N__22715),
            .I(N__22697));
    InMux I__4718 (
            .O(N__22714),
            .I(N__22697));
    InMux I__4717 (
            .O(N__22713),
            .I(N__22694));
    InMux I__4716 (
            .O(N__22710),
            .I(N__22691));
    CascadeMux I__4715 (
            .O(N__22709),
            .I(N__22688));
    InMux I__4714 (
            .O(N__22708),
            .I(N__22685));
    InMux I__4713 (
            .O(N__22707),
            .I(N__22682));
    InMux I__4712 (
            .O(N__22706),
            .I(N__22677));
    InMux I__4711 (
            .O(N__22705),
            .I(N__22677));
    InMux I__4710 (
            .O(N__22704),
            .I(N__22674));
    InMux I__4709 (
            .O(N__22703),
            .I(N__22669));
    InMux I__4708 (
            .O(N__22702),
            .I(N__22666));
    LocalMux I__4707 (
            .O(N__22697),
            .I(N__22659));
    LocalMux I__4706 (
            .O(N__22694),
            .I(N__22659));
    LocalMux I__4705 (
            .O(N__22691),
            .I(N__22659));
    InMux I__4704 (
            .O(N__22688),
            .I(N__22656));
    LocalMux I__4703 (
            .O(N__22685),
            .I(N__22649));
    LocalMux I__4702 (
            .O(N__22682),
            .I(N__22649));
    LocalMux I__4701 (
            .O(N__22677),
            .I(N__22649));
    LocalMux I__4700 (
            .O(N__22674),
            .I(N__22645));
    InMux I__4699 (
            .O(N__22673),
            .I(N__22642));
    InMux I__4698 (
            .O(N__22672),
            .I(N__22639));
    LocalMux I__4697 (
            .O(N__22669),
            .I(N__22636));
    LocalMux I__4696 (
            .O(N__22666),
            .I(N__22633));
    Span4Mux_v I__4695 (
            .O(N__22659),
            .I(N__22630));
    LocalMux I__4694 (
            .O(N__22656),
            .I(N__22627));
    Span4Mux_v I__4693 (
            .O(N__22649),
            .I(N__22624));
    InMux I__4692 (
            .O(N__22648),
            .I(N__22621));
    Span4Mux_v I__4691 (
            .O(N__22645),
            .I(N__22618));
    LocalMux I__4690 (
            .O(N__22642),
            .I(N__22613));
    LocalMux I__4689 (
            .O(N__22639),
            .I(N__22613));
    Span4Mux_h I__4688 (
            .O(N__22636),
            .I(N__22610));
    Span4Mux_h I__4687 (
            .O(N__22633),
            .I(N__22605));
    Span4Mux_h I__4686 (
            .O(N__22630),
            .I(N__22605));
    Span4Mux_v I__4685 (
            .O(N__22627),
            .I(N__22600));
    Span4Mux_h I__4684 (
            .O(N__22624),
            .I(N__22600));
    LocalMux I__4683 (
            .O(N__22621),
            .I(N__22593));
    Span4Mux_h I__4682 (
            .O(N__22618),
            .I(N__22593));
    Span4Mux_v I__4681 (
            .O(N__22613),
            .I(N__22593));
    Odrv4 I__4680 (
            .O(N__22610),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__4679 (
            .O(N__22605),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__4678 (
            .O(N__22600),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__4677 (
            .O(N__22593),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    InMux I__4676 (
            .O(N__22584),
            .I(N__22575));
    InMux I__4675 (
            .O(N__22583),
            .I(N__22572));
    InMux I__4674 (
            .O(N__22582),
            .I(N__22566));
    InMux I__4673 (
            .O(N__22581),
            .I(N__22559));
    InMux I__4672 (
            .O(N__22580),
            .I(N__22559));
    InMux I__4671 (
            .O(N__22579),
            .I(N__22559));
    InMux I__4670 (
            .O(N__22578),
            .I(N__22556));
    LocalMux I__4669 (
            .O(N__22575),
            .I(N__22551));
    LocalMux I__4668 (
            .O(N__22572),
            .I(N__22551));
    InMux I__4667 (
            .O(N__22571),
            .I(N__22546));
    InMux I__4666 (
            .O(N__22570),
            .I(N__22546));
    InMux I__4665 (
            .O(N__22569),
            .I(N__22541));
    LocalMux I__4664 (
            .O(N__22566),
            .I(N__22538));
    LocalMux I__4663 (
            .O(N__22559),
            .I(N__22527));
    LocalMux I__4662 (
            .O(N__22556),
            .I(N__22524));
    Span4Mux_v I__4661 (
            .O(N__22551),
            .I(N__22521));
    LocalMux I__4660 (
            .O(N__22546),
            .I(N__22518));
    InMux I__4659 (
            .O(N__22545),
            .I(N__22513));
    InMux I__4658 (
            .O(N__22544),
            .I(N__22513));
    LocalMux I__4657 (
            .O(N__22541),
            .I(N__22510));
    Span4Mux_h I__4656 (
            .O(N__22538),
            .I(N__22507));
    InMux I__4655 (
            .O(N__22537),
            .I(N__22504));
    CascadeMux I__4654 (
            .O(N__22536),
            .I(N__22498));
    CascadeMux I__4653 (
            .O(N__22535),
            .I(N__22495));
    InMux I__4652 (
            .O(N__22534),
            .I(N__22492));
    InMux I__4651 (
            .O(N__22533),
            .I(N__22489));
    InMux I__4650 (
            .O(N__22532),
            .I(N__22482));
    InMux I__4649 (
            .O(N__22531),
            .I(N__22482));
    InMux I__4648 (
            .O(N__22530),
            .I(N__22482));
    Span4Mux_h I__4647 (
            .O(N__22527),
            .I(N__22471));
    Span4Mux_v I__4646 (
            .O(N__22524),
            .I(N__22471));
    Span4Mux_h I__4645 (
            .O(N__22521),
            .I(N__22471));
    Span4Mux_v I__4644 (
            .O(N__22518),
            .I(N__22471));
    LocalMux I__4643 (
            .O(N__22513),
            .I(N__22471));
    Span4Mux_v I__4642 (
            .O(N__22510),
            .I(N__22464));
    Span4Mux_h I__4641 (
            .O(N__22507),
            .I(N__22464));
    LocalMux I__4640 (
            .O(N__22504),
            .I(N__22464));
    InMux I__4639 (
            .O(N__22503),
            .I(N__22459));
    InMux I__4638 (
            .O(N__22502),
            .I(N__22459));
    InMux I__4637 (
            .O(N__22501),
            .I(N__22452));
    InMux I__4636 (
            .O(N__22498),
            .I(N__22452));
    InMux I__4635 (
            .O(N__22495),
            .I(N__22452));
    LocalMux I__4634 (
            .O(N__22492),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__4633 (
            .O(N__22489),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__4632 (
            .O(N__22482),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__4631 (
            .O(N__22471),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__4630 (
            .O(N__22464),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__4629 (
            .O(N__22459),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__4628 (
            .O(N__22452),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    CascadeMux I__4627 (
            .O(N__22437),
            .I(N__22434));
    InMux I__4626 (
            .O(N__22434),
            .I(N__22430));
    InMux I__4625 (
            .O(N__22433),
            .I(N__22427));
    LocalMux I__4624 (
            .O(N__22430),
            .I(N__22424));
    LocalMux I__4623 (
            .O(N__22427),
            .I(N__22421));
    Span4Mux_h I__4622 (
            .O(N__22424),
            .I(N__22418));
    Odrv4 I__4621 (
            .O(N__22421),
            .I(\this_vga_signals.m58_1 ));
    Odrv4 I__4620 (
            .O(N__22418),
            .I(\this_vga_signals.m58_1 ));
    InMux I__4619 (
            .O(N__22413),
            .I(N__22410));
    LocalMux I__4618 (
            .O(N__22410),
            .I(\this_vga_signals.m58_0 ));
    CascadeMux I__4617 (
            .O(N__22407),
            .I(\this_vga_signals.m58_4_cascade_ ));
    CascadeMux I__4616 (
            .O(N__22404),
            .I(N__22397));
    InMux I__4615 (
            .O(N__22403),
            .I(N__22394));
    CascadeMux I__4614 (
            .O(N__22402),
            .I(N__22388));
    InMux I__4613 (
            .O(N__22401),
            .I(N__22383));
    InMux I__4612 (
            .O(N__22400),
            .I(N__22380));
    InMux I__4611 (
            .O(N__22397),
            .I(N__22377));
    LocalMux I__4610 (
            .O(N__22394),
            .I(N__22374));
    InMux I__4609 (
            .O(N__22393),
            .I(N__22367));
    InMux I__4608 (
            .O(N__22392),
            .I(N__22367));
    InMux I__4607 (
            .O(N__22391),
            .I(N__22367));
    InMux I__4606 (
            .O(N__22388),
            .I(N__22364));
    InMux I__4605 (
            .O(N__22387),
            .I(N__22357));
    InMux I__4604 (
            .O(N__22386),
            .I(N__22353));
    LocalMux I__4603 (
            .O(N__22383),
            .I(N__22348));
    LocalMux I__4602 (
            .O(N__22380),
            .I(N__22345));
    LocalMux I__4601 (
            .O(N__22377),
            .I(N__22342));
    Span4Mux_v I__4600 (
            .O(N__22374),
            .I(N__22335));
    LocalMux I__4599 (
            .O(N__22367),
            .I(N__22335));
    LocalMux I__4598 (
            .O(N__22364),
            .I(N__22335));
    CascadeMux I__4597 (
            .O(N__22363),
            .I(N__22331));
    InMux I__4596 (
            .O(N__22362),
            .I(N__22328));
    InMux I__4595 (
            .O(N__22361),
            .I(N__22324));
    InMux I__4594 (
            .O(N__22360),
            .I(N__22321));
    LocalMux I__4593 (
            .O(N__22357),
            .I(N__22317));
    InMux I__4592 (
            .O(N__22356),
            .I(N__22313));
    LocalMux I__4591 (
            .O(N__22353),
            .I(N__22310));
    InMux I__4590 (
            .O(N__22352),
            .I(N__22305));
    InMux I__4589 (
            .O(N__22351),
            .I(N__22305));
    Span4Mux_v I__4588 (
            .O(N__22348),
            .I(N__22296));
    Span4Mux_h I__4587 (
            .O(N__22345),
            .I(N__22296));
    Span4Mux_v I__4586 (
            .O(N__22342),
            .I(N__22296));
    Span4Mux_v I__4585 (
            .O(N__22335),
            .I(N__22296));
    InMux I__4584 (
            .O(N__22334),
            .I(N__22291));
    InMux I__4583 (
            .O(N__22331),
            .I(N__22291));
    LocalMux I__4582 (
            .O(N__22328),
            .I(N__22288));
    CascadeMux I__4581 (
            .O(N__22327),
            .I(N__22285));
    LocalMux I__4580 (
            .O(N__22324),
            .I(N__22282));
    LocalMux I__4579 (
            .O(N__22321),
            .I(N__22279));
    InMux I__4578 (
            .O(N__22320),
            .I(N__22276));
    Span4Mux_h I__4577 (
            .O(N__22317),
            .I(N__22273));
    CascadeMux I__4576 (
            .O(N__22316),
            .I(N__22266));
    LocalMux I__4575 (
            .O(N__22313),
            .I(N__22257));
    Span4Mux_h I__4574 (
            .O(N__22310),
            .I(N__22257));
    LocalMux I__4573 (
            .O(N__22305),
            .I(N__22257));
    Span4Mux_h I__4572 (
            .O(N__22296),
            .I(N__22250));
    LocalMux I__4571 (
            .O(N__22291),
            .I(N__22250));
    Span4Mux_h I__4570 (
            .O(N__22288),
            .I(N__22250));
    InMux I__4569 (
            .O(N__22285),
            .I(N__22247));
    Span4Mux_v I__4568 (
            .O(N__22282),
            .I(N__22244));
    Span4Mux_v I__4567 (
            .O(N__22279),
            .I(N__22237));
    LocalMux I__4566 (
            .O(N__22276),
            .I(N__22237));
    Span4Mux_v I__4565 (
            .O(N__22273),
            .I(N__22237));
    InMux I__4564 (
            .O(N__22272),
            .I(N__22228));
    InMux I__4563 (
            .O(N__22271),
            .I(N__22228));
    InMux I__4562 (
            .O(N__22270),
            .I(N__22228));
    InMux I__4561 (
            .O(N__22269),
            .I(N__22228));
    InMux I__4560 (
            .O(N__22266),
            .I(N__22225));
    InMux I__4559 (
            .O(N__22265),
            .I(N__22220));
    InMux I__4558 (
            .O(N__22264),
            .I(N__22220));
    Span4Mux_v I__4557 (
            .O(N__22257),
            .I(N__22213));
    Span4Mux_v I__4556 (
            .O(N__22250),
            .I(N__22213));
    LocalMux I__4555 (
            .O(N__22247),
            .I(N__22213));
    Odrv4 I__4554 (
            .O(N__22244),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__4553 (
            .O(N__22237),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__4552 (
            .O(N__22228),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__4551 (
            .O(N__22225),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__4550 (
            .O(N__22220),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__4549 (
            .O(N__22213),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    IoInMux I__4548 (
            .O(N__22200),
            .I(N__22197));
    LocalMux I__4547 (
            .O(N__22197),
            .I(N__22194));
    Span4Mux_s1_v I__4546 (
            .O(N__22194),
            .I(N__22191));
    Sp12to4 I__4545 (
            .O(N__22191),
            .I(N__22188));
    Span12Mux_s8_h I__4544 (
            .O(N__22188),
            .I(N__22185));
    Span12Mux_h I__4543 (
            .O(N__22185),
            .I(N__22182));
    Odrv12 I__4542 (
            .O(N__22182),
            .I(this_vga_signals_vsync_1_i));
    InMux I__4541 (
            .O(N__22179),
            .I(N__22175));
    InMux I__4540 (
            .O(N__22178),
            .I(N__22172));
    LocalMux I__4539 (
            .O(N__22175),
            .I(N__22168));
    LocalMux I__4538 (
            .O(N__22172),
            .I(N__22164));
    InMux I__4537 (
            .O(N__22171),
            .I(N__22160));
    Span4Mux_h I__4536 (
            .O(N__22168),
            .I(N__22157));
    InMux I__4535 (
            .O(N__22167),
            .I(N__22154));
    Span4Mux_h I__4534 (
            .O(N__22164),
            .I(N__22151));
    InMux I__4533 (
            .O(N__22163),
            .I(N__22148));
    LocalMux I__4532 (
            .O(N__22160),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__4531 (
            .O(N__22157),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__4530 (
            .O(N__22154),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__4529 (
            .O(N__22151),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__4528 (
            .O(N__22148),
            .I(M_this_state_qZ0Z_3));
    CascadeMux I__4527 (
            .O(N__22137),
            .I(\this_start_data_delay.N_123_cascade_ ));
    InMux I__4526 (
            .O(N__22134),
            .I(N__22130));
    InMux I__4525 (
            .O(N__22133),
            .I(N__22126));
    LocalMux I__4524 (
            .O(N__22130),
            .I(N__22122));
    InMux I__4523 (
            .O(N__22129),
            .I(N__22119));
    LocalMux I__4522 (
            .O(N__22126),
            .I(N__22115));
    InMux I__4521 (
            .O(N__22125),
            .I(N__22112));
    Span4Mux_h I__4520 (
            .O(N__22122),
            .I(N__22108));
    LocalMux I__4519 (
            .O(N__22119),
            .I(N__22105));
    InMux I__4518 (
            .O(N__22118),
            .I(N__22102));
    Span4Mux_v I__4517 (
            .O(N__22115),
            .I(N__22097));
    LocalMux I__4516 (
            .O(N__22112),
            .I(N__22097));
    InMux I__4515 (
            .O(N__22111),
            .I(N__22094));
    Span4Mux_v I__4514 (
            .O(N__22108),
            .I(N__22087));
    Span4Mux_h I__4513 (
            .O(N__22105),
            .I(N__22087));
    LocalMux I__4512 (
            .O(N__22102),
            .I(N__22084));
    Span4Mux_v I__4511 (
            .O(N__22097),
            .I(N__22079));
    LocalMux I__4510 (
            .O(N__22094),
            .I(N__22079));
    InMux I__4509 (
            .O(N__22093),
            .I(N__22076));
    InMux I__4508 (
            .O(N__22092),
            .I(N__22073));
    Span4Mux_v I__4507 (
            .O(N__22087),
            .I(N__22068));
    Span4Mux_h I__4506 (
            .O(N__22084),
            .I(N__22068));
    Span4Mux_v I__4505 (
            .O(N__22079),
            .I(N__22063));
    LocalMux I__4504 (
            .O(N__22076),
            .I(N__22063));
    LocalMux I__4503 (
            .O(N__22073),
            .I(N__22060));
    Span4Mux_v I__4502 (
            .O(N__22068),
            .I(N__22053));
    Span4Mux_h I__4501 (
            .O(N__22063),
            .I(N__22053));
    Span4Mux_h I__4500 (
            .O(N__22060),
            .I(N__22053));
    Odrv4 I__4499 (
            .O(N__22053),
            .I(N_812_0));
    InMux I__4498 (
            .O(N__22050),
            .I(bfn_21_21_0_));
    InMux I__4497 (
            .O(N__22047),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    CascadeMux I__4496 (
            .O(N__22044),
            .I(N__22041));
    InMux I__4495 (
            .O(N__22041),
            .I(N__22038));
    LocalMux I__4494 (
            .O(N__22038),
            .I(N__22035));
    Odrv4 I__4493 (
            .O(N__22035),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    InMux I__4492 (
            .O(N__22032),
            .I(N__22023));
    InMux I__4491 (
            .O(N__22031),
            .I(N__22023));
    InMux I__4490 (
            .O(N__22030),
            .I(N__22023));
    LocalMux I__4489 (
            .O(N__22023),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    CascadeMux I__4488 (
            .O(N__22020),
            .I(N__22017));
    InMux I__4487 (
            .O(N__22017),
            .I(N__22014));
    LocalMux I__4486 (
            .O(N__22014),
            .I(N__22011));
    Span4Mux_v I__4485 (
            .O(N__22011),
            .I(N__22008));
    Span4Mux_h I__4484 (
            .O(N__22008),
            .I(N__22005));
    Odrv4 I__4483 (
            .O(N__22005),
            .I(\this_vga_signals.N_4557_0 ));
    InMux I__4482 (
            .O(N__22002),
            .I(N__21994));
    InMux I__4481 (
            .O(N__22001),
            .I(N__21994));
    InMux I__4480 (
            .O(N__22000),
            .I(N__21991));
    InMux I__4479 (
            .O(N__21999),
            .I(N__21986));
    LocalMux I__4478 (
            .O(N__21994),
            .I(N__21982));
    LocalMux I__4477 (
            .O(N__21991),
            .I(N__21979));
    InMux I__4476 (
            .O(N__21990),
            .I(N__21974));
    InMux I__4475 (
            .O(N__21989),
            .I(N__21974));
    LocalMux I__4474 (
            .O(N__21986),
            .I(N__21971));
    InMux I__4473 (
            .O(N__21985),
            .I(N__21968));
    Span4Mux_h I__4472 (
            .O(N__21982),
            .I(N__21964));
    Span4Mux_v I__4471 (
            .O(N__21979),
            .I(N__21957));
    LocalMux I__4470 (
            .O(N__21974),
            .I(N__21957));
    Span4Mux_v I__4469 (
            .O(N__21971),
            .I(N__21952));
    LocalMux I__4468 (
            .O(N__21968),
            .I(N__21952));
    InMux I__4467 (
            .O(N__21967),
            .I(N__21943));
    Span4Mux_h I__4466 (
            .O(N__21964),
            .I(N__21940));
    InMux I__4465 (
            .O(N__21963),
            .I(N__21935));
    InMux I__4464 (
            .O(N__21962),
            .I(N__21935));
    Span4Mux_h I__4463 (
            .O(N__21957),
            .I(N__21930));
    Span4Mux_v I__4462 (
            .O(N__21952),
            .I(N__21930));
    InMux I__4461 (
            .O(N__21951),
            .I(N__21923));
    InMux I__4460 (
            .O(N__21950),
            .I(N__21923));
    InMux I__4459 (
            .O(N__21949),
            .I(N__21923));
    InMux I__4458 (
            .O(N__21948),
            .I(N__21916));
    InMux I__4457 (
            .O(N__21947),
            .I(N__21916));
    InMux I__4456 (
            .O(N__21946),
            .I(N__21916));
    LocalMux I__4455 (
            .O(N__21943),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__4454 (
            .O(N__21940),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__4453 (
            .O(N__21935),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__4452 (
            .O(N__21930),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__4451 (
            .O(N__21923),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__4450 (
            .O(N__21916),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    InMux I__4449 (
            .O(N__21903),
            .I(N__21898));
    InMux I__4448 (
            .O(N__21902),
            .I(N__21894));
    InMux I__4447 (
            .O(N__21901),
            .I(N__21889));
    LocalMux I__4446 (
            .O(N__21898),
            .I(N__21886));
    InMux I__4445 (
            .O(N__21897),
            .I(N__21883));
    LocalMux I__4444 (
            .O(N__21894),
            .I(N__21879));
    InMux I__4443 (
            .O(N__21893),
            .I(N__21874));
    InMux I__4442 (
            .O(N__21892),
            .I(N__21874));
    LocalMux I__4441 (
            .O(N__21889),
            .I(N__21868));
    Span4Mux_v I__4440 (
            .O(N__21886),
            .I(N__21863));
    LocalMux I__4439 (
            .O(N__21883),
            .I(N__21863));
    InMux I__4438 (
            .O(N__21882),
            .I(N__21857));
    Span12Mux_s11_v I__4437 (
            .O(N__21879),
            .I(N__21852));
    LocalMux I__4436 (
            .O(N__21874),
            .I(N__21852));
    InMux I__4435 (
            .O(N__21873),
            .I(N__21847));
    InMux I__4434 (
            .O(N__21872),
            .I(N__21847));
    InMux I__4433 (
            .O(N__21871),
            .I(N__21844));
    Span4Mux_h I__4432 (
            .O(N__21868),
            .I(N__21839));
    Span4Mux_h I__4431 (
            .O(N__21863),
            .I(N__21839));
    InMux I__4430 (
            .O(N__21862),
            .I(N__21832));
    InMux I__4429 (
            .O(N__21861),
            .I(N__21832));
    InMux I__4428 (
            .O(N__21860),
            .I(N__21832));
    LocalMux I__4427 (
            .O(N__21857),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv12 I__4426 (
            .O(N__21852),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__4425 (
            .O(N__21847),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__4424 (
            .O(N__21844),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__4423 (
            .O(N__21839),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__4422 (
            .O(N__21832),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    InMux I__4421 (
            .O(N__21819),
            .I(N__21815));
    CascadeMux I__4420 (
            .O(N__21818),
            .I(N__21807));
    LocalMux I__4419 (
            .O(N__21815),
            .I(N__21803));
    InMux I__4418 (
            .O(N__21814),
            .I(N__21800));
    InMux I__4417 (
            .O(N__21813),
            .I(N__21795));
    InMux I__4416 (
            .O(N__21812),
            .I(N__21795));
    InMux I__4415 (
            .O(N__21811),
            .I(N__21786));
    InMux I__4414 (
            .O(N__21810),
            .I(N__21786));
    InMux I__4413 (
            .O(N__21807),
            .I(N__21786));
    InMux I__4412 (
            .O(N__21806),
            .I(N__21786));
    Odrv4 I__4411 (
            .O(N__21803),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__4410 (
            .O(N__21800),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__4409 (
            .O(N__21795),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__4408 (
            .O(N__21786),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    CascadeMux I__4407 (
            .O(N__21777),
            .I(N__21771));
    InMux I__4406 (
            .O(N__21776),
            .I(N__21765));
    InMux I__4405 (
            .O(N__21775),
            .I(N__21762));
    InMux I__4404 (
            .O(N__21774),
            .I(N__21759));
    InMux I__4403 (
            .O(N__21771),
            .I(N__21756));
    InMux I__4402 (
            .O(N__21770),
            .I(N__21751));
    InMux I__4401 (
            .O(N__21769),
            .I(N__21751));
    InMux I__4400 (
            .O(N__21768),
            .I(N__21748));
    LocalMux I__4399 (
            .O(N__21765),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__4398 (
            .O(N__21762),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__4397 (
            .O(N__21759),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__4396 (
            .O(N__21756),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__4395 (
            .O(N__21751),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__4394 (
            .O(N__21748),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    InMux I__4393 (
            .O(N__21735),
            .I(N__21729));
    InMux I__4392 (
            .O(N__21734),
            .I(N__21729));
    LocalMux I__4391 (
            .O(N__21729),
            .I(N__21726));
    Span4Mux_h I__4390 (
            .O(N__21726),
            .I(N__21723));
    Odrv4 I__4389 (
            .O(N__21723),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_601 ));
    InMux I__4388 (
            .O(N__21720),
            .I(N__21716));
    InMux I__4387 (
            .O(N__21719),
            .I(N__21712));
    LocalMux I__4386 (
            .O(N__21716),
            .I(N__21709));
    InMux I__4385 (
            .O(N__21715),
            .I(N__21706));
    LocalMux I__4384 (
            .O(N__21712),
            .I(N__21703));
    Span4Mux_v I__4383 (
            .O(N__21709),
            .I(N__21698));
    LocalMux I__4382 (
            .O(N__21706),
            .I(N__21698));
    Odrv4 I__4381 (
            .O(N__21703),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    Odrv4 I__4380 (
            .O(N__21698),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    InMux I__4379 (
            .O(N__21693),
            .I(N__21687));
    InMux I__4378 (
            .O(N__21692),
            .I(N__21680));
    InMux I__4377 (
            .O(N__21691),
            .I(N__21680));
    InMux I__4376 (
            .O(N__21690),
            .I(N__21680));
    LocalMux I__4375 (
            .O(N__21687),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__4374 (
            .O(N__21680),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    CascadeMux I__4373 (
            .O(N__21675),
            .I(N__21671));
    InMux I__4372 (
            .O(N__21674),
            .I(N__21667));
    InMux I__4371 (
            .O(N__21671),
            .I(N__21664));
    InMux I__4370 (
            .O(N__21670),
            .I(N__21657));
    LocalMux I__4369 (
            .O(N__21667),
            .I(N__21654));
    LocalMux I__4368 (
            .O(N__21664),
            .I(N__21651));
    InMux I__4367 (
            .O(N__21663),
            .I(N__21648));
    InMux I__4366 (
            .O(N__21662),
            .I(N__21643));
    InMux I__4365 (
            .O(N__21661),
            .I(N__21643));
    InMux I__4364 (
            .O(N__21660),
            .I(N__21640));
    LocalMux I__4363 (
            .O(N__21657),
            .I(N__21634));
    Span4Mux_v I__4362 (
            .O(N__21654),
            .I(N__21631));
    Span4Mux_v I__4361 (
            .O(N__21651),
            .I(N__21628));
    LocalMux I__4360 (
            .O(N__21648),
            .I(N__21623));
    LocalMux I__4359 (
            .O(N__21643),
            .I(N__21623));
    LocalMux I__4358 (
            .O(N__21640),
            .I(N__21619));
    InMux I__4357 (
            .O(N__21639),
            .I(N__21616));
    InMux I__4356 (
            .O(N__21638),
            .I(N__21613));
    InMux I__4355 (
            .O(N__21637),
            .I(N__21610));
    Span4Mux_h I__4354 (
            .O(N__21634),
            .I(N__21607));
    Span4Mux_h I__4353 (
            .O(N__21631),
            .I(N__21602));
    Span4Mux_h I__4352 (
            .O(N__21628),
            .I(N__21602));
    Span4Mux_h I__4351 (
            .O(N__21623),
            .I(N__21599));
    InMux I__4350 (
            .O(N__21622),
            .I(N__21596));
    Odrv4 I__4349 (
            .O(N__21619),
            .I(this_vga_signals_M_hcounter_d7_0));
    LocalMux I__4348 (
            .O(N__21616),
            .I(this_vga_signals_M_hcounter_d7_0));
    LocalMux I__4347 (
            .O(N__21613),
            .I(this_vga_signals_M_hcounter_d7_0));
    LocalMux I__4346 (
            .O(N__21610),
            .I(this_vga_signals_M_hcounter_d7_0));
    Odrv4 I__4345 (
            .O(N__21607),
            .I(this_vga_signals_M_hcounter_d7_0));
    Odrv4 I__4344 (
            .O(N__21602),
            .I(this_vga_signals_M_hcounter_d7_0));
    Odrv4 I__4343 (
            .O(N__21599),
            .I(this_vga_signals_M_hcounter_d7_0));
    LocalMux I__4342 (
            .O(N__21596),
            .I(this_vga_signals_M_hcounter_d7_0));
    InMux I__4341 (
            .O(N__21579),
            .I(N__21575));
    InMux I__4340 (
            .O(N__21578),
            .I(N__21572));
    LocalMux I__4339 (
            .O(N__21575),
            .I(N__21569));
    LocalMux I__4338 (
            .O(N__21572),
            .I(N__21565));
    Span4Mux_h I__4337 (
            .O(N__21569),
            .I(N__21562));
    InMux I__4336 (
            .O(N__21568),
            .I(N__21559));
    Span12Mux_h I__4335 (
            .O(N__21565),
            .I(N__21556));
    Span4Mux_h I__4334 (
            .O(N__21562),
            .I(N__21553));
    LocalMux I__4333 (
            .O(N__21559),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv12 I__4332 (
            .O(N__21556),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv4 I__4331 (
            .O(N__21553),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    InMux I__4330 (
            .O(N__21546),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    InMux I__4329 (
            .O(N__21543),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__4328 (
            .O(N__21540),
            .I(N__21531));
    InMux I__4327 (
            .O(N__21539),
            .I(N__21531));
    InMux I__4326 (
            .O(N__21538),
            .I(N__21526));
    InMux I__4325 (
            .O(N__21537),
            .I(N__21526));
    InMux I__4324 (
            .O(N__21536),
            .I(N__21518));
    LocalMux I__4323 (
            .O(N__21531),
            .I(N__21515));
    LocalMux I__4322 (
            .O(N__21526),
            .I(N__21512));
    InMux I__4321 (
            .O(N__21525),
            .I(N__21509));
    CEMux I__4320 (
            .O(N__21524),
            .I(N__21506));
    InMux I__4319 (
            .O(N__21523),
            .I(N__21501));
    InMux I__4318 (
            .O(N__21522),
            .I(N__21501));
    InMux I__4317 (
            .O(N__21521),
            .I(N__21498));
    LocalMux I__4316 (
            .O(N__21518),
            .I(N__21485));
    Span4Mux_v I__4315 (
            .O(N__21515),
            .I(N__21482));
    Span4Mux_v I__4314 (
            .O(N__21512),
            .I(N__21479));
    LocalMux I__4313 (
            .O(N__21509),
            .I(N__21473));
    LocalMux I__4312 (
            .O(N__21506),
            .I(N__21466));
    LocalMux I__4311 (
            .O(N__21501),
            .I(N__21466));
    LocalMux I__4310 (
            .O(N__21498),
            .I(N__21466));
    InMux I__4309 (
            .O(N__21497),
            .I(N__21461));
    InMux I__4308 (
            .O(N__21496),
            .I(N__21461));
    InMux I__4307 (
            .O(N__21495),
            .I(N__21458));
    InMux I__4306 (
            .O(N__21494),
            .I(N__21449));
    InMux I__4305 (
            .O(N__21493),
            .I(N__21449));
    InMux I__4304 (
            .O(N__21492),
            .I(N__21449));
    InMux I__4303 (
            .O(N__21491),
            .I(N__21449));
    InMux I__4302 (
            .O(N__21490),
            .I(N__21442));
    InMux I__4301 (
            .O(N__21489),
            .I(N__21442));
    InMux I__4300 (
            .O(N__21488),
            .I(N__21442));
    Span4Mux_v I__4299 (
            .O(N__21485),
            .I(N__21435));
    Span4Mux_h I__4298 (
            .O(N__21482),
            .I(N__21435));
    Span4Mux_h I__4297 (
            .O(N__21479),
            .I(N__21435));
    InMux I__4296 (
            .O(N__21478),
            .I(N__21432));
    InMux I__4295 (
            .O(N__21477),
            .I(N__21429));
    InMux I__4294 (
            .O(N__21476),
            .I(N__21426));
    Span4Mux_h I__4293 (
            .O(N__21473),
            .I(N__21423));
    Span4Mux_v I__4292 (
            .O(N__21466),
            .I(N__21420));
    LocalMux I__4291 (
            .O(N__21461),
            .I(N__21417));
    LocalMux I__4290 (
            .O(N__21458),
            .I(N__21402));
    LocalMux I__4289 (
            .O(N__21449),
            .I(N__21402));
    LocalMux I__4288 (
            .O(N__21442),
            .I(N__21402));
    Sp12to4 I__4287 (
            .O(N__21435),
            .I(N__21402));
    LocalMux I__4286 (
            .O(N__21432),
            .I(N__21402));
    LocalMux I__4285 (
            .O(N__21429),
            .I(N__21402));
    LocalMux I__4284 (
            .O(N__21426),
            .I(N__21402));
    Odrv4 I__4283 (
            .O(N__21423),
            .I(G_442));
    Odrv4 I__4282 (
            .O(N__21420),
            .I(G_442));
    Odrv4 I__4281 (
            .O(N__21417),
            .I(G_442));
    Odrv12 I__4280 (
            .O(N__21402),
            .I(G_442));
    InMux I__4279 (
            .O(N__21393),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__4278 (
            .O(N__21390),
            .I(N__21386));
    InMux I__4277 (
            .O(N__21389),
            .I(N__21382));
    LocalMux I__4276 (
            .O(N__21386),
            .I(N__21379));
    InMux I__4275 (
            .O(N__21385),
            .I(N__21376));
    LocalMux I__4274 (
            .O(N__21382),
            .I(N__21373));
    Span4Mux_v I__4273 (
            .O(N__21379),
            .I(N__21368));
    LocalMux I__4272 (
            .O(N__21376),
            .I(N__21368));
    Span4Mux_h I__4271 (
            .O(N__21373),
            .I(N__21365));
    Span4Mux_v I__4270 (
            .O(N__21368),
            .I(N__21362));
    Odrv4 I__4269 (
            .O(N__21365),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    Odrv4 I__4268 (
            .O(N__21362),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    InMux I__4267 (
            .O(N__21357),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__4266 (
            .O(N__21354),
            .I(N__21345));
    InMux I__4265 (
            .O(N__21353),
            .I(N__21345));
    InMux I__4264 (
            .O(N__21352),
            .I(N__21345));
    LocalMux I__4263 (
            .O(N__21345),
            .I(N__21342));
    Span4Mux_h I__4262 (
            .O(N__21342),
            .I(N__21339));
    Odrv4 I__4261 (
            .O(N__21339),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    InMux I__4260 (
            .O(N__21336),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__4259 (
            .O(N__21333),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__4258 (
            .O(N__21330),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    CascadeMux I__4257 (
            .O(N__21327),
            .I(\this_start_data_delay.N_91_0_cascade_ ));
    InMux I__4256 (
            .O(N__21324),
            .I(N__21313));
    InMux I__4255 (
            .O(N__21323),
            .I(N__21313));
    InMux I__4254 (
            .O(N__21322),
            .I(N__21310));
    InMux I__4253 (
            .O(N__21321),
            .I(N__21307));
    InMux I__4252 (
            .O(N__21320),
            .I(N__21304));
    InMux I__4251 (
            .O(N__21319),
            .I(N__21299));
    InMux I__4250 (
            .O(N__21318),
            .I(N__21299));
    LocalMux I__4249 (
            .O(N__21313),
            .I(N__21292));
    LocalMux I__4248 (
            .O(N__21310),
            .I(N__21292));
    LocalMux I__4247 (
            .O(N__21307),
            .I(N__21292));
    LocalMux I__4246 (
            .O(N__21304),
            .I(N__21289));
    LocalMux I__4245 (
            .O(N__21299),
            .I(N__21284));
    Span4Mux_v I__4244 (
            .O(N__21292),
            .I(N__21284));
    Odrv4 I__4243 (
            .O(N__21289),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__4242 (
            .O(N__21284),
            .I(M_this_state_qZ0Z_1));
    CascadeMux I__4241 (
            .O(N__21279),
            .I(\this_start_data_delay.N_110_cascade_ ));
    CascadeMux I__4240 (
            .O(N__21276),
            .I(N__21273));
    InMux I__4239 (
            .O(N__21273),
            .I(N__21267));
    InMux I__4238 (
            .O(N__21272),
            .I(N__21267));
    LocalMux I__4237 (
            .O(N__21267),
            .I(N__21264));
    Span4Mux_h I__4236 (
            .O(N__21264),
            .I(N__21259));
    InMux I__4235 (
            .O(N__21263),
            .I(N__21254));
    InMux I__4234 (
            .O(N__21262),
            .I(N__21254));
    Odrv4 I__4233 (
            .O(N__21259),
            .I(M_this_state_qZ0Z_4));
    LocalMux I__4232 (
            .O(N__21254),
            .I(M_this_state_qZ0Z_4));
    InMux I__4231 (
            .O(N__21249),
            .I(N__21246));
    LocalMux I__4230 (
            .O(N__21246),
            .I(N__21243));
    Span4Mux_h I__4229 (
            .O(N__21243),
            .I(N__21240));
    Odrv4 I__4228 (
            .O(N__21240),
            .I(\this_sprites_ram.mem_out_bus5_1 ));
    InMux I__4227 (
            .O(N__21237),
            .I(N__21234));
    LocalMux I__4226 (
            .O(N__21234),
            .I(N__21231));
    Span4Mux_h I__4225 (
            .O(N__21231),
            .I(N__21228));
    Sp12to4 I__4224 (
            .O(N__21228),
            .I(N__21225));
    Span12Mux_v I__4223 (
            .O(N__21225),
            .I(N__21222));
    Odrv12 I__4222 (
            .O(N__21222),
            .I(\this_sprites_ram.mem_out_bus1_1 ));
    InMux I__4221 (
            .O(N__21219),
            .I(N__21216));
    LocalMux I__4220 (
            .O(N__21216),
            .I(N__21213));
    Span4Mux_h I__4219 (
            .O(N__21213),
            .I(N__21210));
    Span4Mux_v I__4218 (
            .O(N__21210),
            .I(N__21207));
    Odrv4 I__4217 (
            .O(N__21207),
            .I(\this_sprites_ram.mem_out_bus6_1 ));
    InMux I__4216 (
            .O(N__21204),
            .I(N__21201));
    LocalMux I__4215 (
            .O(N__21201),
            .I(N__21198));
    Span4Mux_v I__4214 (
            .O(N__21198),
            .I(N__21195));
    Span4Mux_h I__4213 (
            .O(N__21195),
            .I(N__21192));
    Span4Mux_v I__4212 (
            .O(N__21192),
            .I(N__21189));
    Odrv4 I__4211 (
            .O(N__21189),
            .I(\this_sprites_ram.mem_out_bus2_1 ));
    CascadeMux I__4210 (
            .O(N__21186),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0_cascade_ ));
    InMux I__4209 (
            .O(N__21183),
            .I(N__21180));
    LocalMux I__4208 (
            .O(N__21180),
            .I(N__21177));
    Span12Mux_v I__4207 (
            .O(N__21177),
            .I(N__21174));
    Odrv12 I__4206 (
            .O(N__21174),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ));
    CascadeMux I__4205 (
            .O(N__21171),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ));
    InMux I__4204 (
            .O(N__21168),
            .I(N__21165));
    LocalMux I__4203 (
            .O(N__21165),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ));
    InMux I__4202 (
            .O(N__21162),
            .I(N__21157));
    InMux I__4201 (
            .O(N__21161),
            .I(N__21154));
    InMux I__4200 (
            .O(N__21160),
            .I(N__21151));
    LocalMux I__4199 (
            .O(N__21157),
            .I(N__21148));
    LocalMux I__4198 (
            .O(N__21154),
            .I(N__21145));
    LocalMux I__4197 (
            .O(N__21151),
            .I(N__21142));
    Span12Mux_s8_h I__4196 (
            .O(N__21148),
            .I(N__21139));
    Span4Mux_h I__4195 (
            .O(N__21145),
            .I(N__21136));
    Span4Mux_h I__4194 (
            .O(N__21142),
            .I(N__21133));
    Span12Mux_h I__4193 (
            .O(N__21139),
            .I(N__21130));
    Span4Mux_h I__4192 (
            .O(N__21136),
            .I(N__21127));
    Span4Mux_h I__4191 (
            .O(N__21133),
            .I(N__21124));
    Odrv12 I__4190 (
            .O(N__21130),
            .I(M_this_ppu_vram_data_1));
    Odrv4 I__4189 (
            .O(N__21127),
            .I(M_this_ppu_vram_data_1));
    Odrv4 I__4188 (
            .O(N__21124),
            .I(M_this_ppu_vram_data_1));
    CascadeMux I__4187 (
            .O(N__21117),
            .I(N__21114));
    InMux I__4186 (
            .O(N__21114),
            .I(N__21111));
    LocalMux I__4185 (
            .O(N__21111),
            .I(\this_start_data_delay.M_this_state_q_ns_0_i_2_0 ));
    CascadeMux I__4184 (
            .O(N__21108),
            .I(N_554_0_cascade_));
    CascadeMux I__4183 (
            .O(N__21105),
            .I(N__21102));
    InMux I__4182 (
            .O(N__21102),
            .I(N__21094));
    InMux I__4181 (
            .O(N__21101),
            .I(N__21094));
    InMux I__4180 (
            .O(N__21100),
            .I(N__21090));
    InMux I__4179 (
            .O(N__21099),
            .I(N__21085));
    LocalMux I__4178 (
            .O(N__21094),
            .I(N__21082));
    InMux I__4177 (
            .O(N__21093),
            .I(N__21079));
    LocalMux I__4176 (
            .O(N__21090),
            .I(N__21076));
    InMux I__4175 (
            .O(N__21089),
            .I(N__21073));
    InMux I__4174 (
            .O(N__21088),
            .I(N__21070));
    LocalMux I__4173 (
            .O(N__21085),
            .I(N__21067));
    Span4Mux_v I__4172 (
            .O(N__21082),
            .I(N__21064));
    LocalMux I__4171 (
            .O(N__21079),
            .I(N__21057));
    Span4Mux_h I__4170 (
            .O(N__21076),
            .I(N__21057));
    LocalMux I__4169 (
            .O(N__21073),
            .I(N__21057));
    LocalMux I__4168 (
            .O(N__21070),
            .I(M_this_state_qZ0Z_2));
    Odrv12 I__4167 (
            .O(N__21067),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__4166 (
            .O(N__21064),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__4165 (
            .O(N__21057),
            .I(M_this_state_qZ0Z_2));
    CascadeMux I__4164 (
            .O(N__21048),
            .I(\this_start_data_delay.N_109_cascade_ ));
    InMux I__4163 (
            .O(N__21045),
            .I(N__21042));
    LocalMux I__4162 (
            .O(N__21042),
            .I(N__21039));
    Odrv4 I__4161 (
            .O(N__21039),
            .I(\this_start_data_delay.M_this_sprites_address_q_0_0_0_4 ));
    InMux I__4160 (
            .O(N__21036),
            .I(N__21033));
    LocalMux I__4159 (
            .O(N__21033),
            .I(N__21030));
    Odrv12 I__4158 (
            .O(N__21030),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    InMux I__4157 (
            .O(N__21027),
            .I(N__21020));
    InMux I__4156 (
            .O(N__21026),
            .I(N__21020));
    InMux I__4155 (
            .O(N__21025),
            .I(N__21017));
    LocalMux I__4154 (
            .O(N__21020),
            .I(\this_start_data_delay.M_last_qZ0 ));
    LocalMux I__4153 (
            .O(N__21017),
            .I(\this_start_data_delay.M_last_qZ0 ));
    InMux I__4152 (
            .O(N__21012),
            .I(N__21004));
    InMux I__4151 (
            .O(N__21011),
            .I(N__21004));
    InMux I__4150 (
            .O(N__21010),
            .I(N__20999));
    InMux I__4149 (
            .O(N__21009),
            .I(N__20999));
    LocalMux I__4148 (
            .O(N__21004),
            .I(N__20994));
    LocalMux I__4147 (
            .O(N__20999),
            .I(N__20994));
    Span4Mux_v I__4146 (
            .O(N__20994),
            .I(N__20991));
    Span4Mux_h I__4145 (
            .O(N__20991),
            .I(N__20988));
    Sp12to4 I__4144 (
            .O(N__20988),
            .I(N__20985));
    Span12Mux_h I__4143 (
            .O(N__20985),
            .I(N__20982));
    Odrv12 I__4142 (
            .O(N__20982),
            .I(port_enb_c));
    InMux I__4141 (
            .O(N__20979),
            .I(N__20971));
    InMux I__4140 (
            .O(N__20978),
            .I(N__20971));
    InMux I__4139 (
            .O(N__20977),
            .I(N__20966));
    InMux I__4138 (
            .O(N__20976),
            .I(N__20966));
    LocalMux I__4137 (
            .O(N__20971),
            .I(M_this_delay_clk_out_0));
    LocalMux I__4136 (
            .O(N__20966),
            .I(M_this_delay_clk_out_0));
    InMux I__4135 (
            .O(N__20961),
            .I(N__20958));
    LocalMux I__4134 (
            .O(N__20958),
            .I(\this_vga_signals.vaddress_1_6 ));
    InMux I__4133 (
            .O(N__20955),
            .I(N__20952));
    LocalMux I__4132 (
            .O(N__20952),
            .I(N__20949));
    Span12Mux_h I__4131 (
            .O(N__20949),
            .I(N__20946));
    Span12Mux_v I__4130 (
            .O(N__20946),
            .I(N__20943));
    Odrv12 I__4129 (
            .O(N__20943),
            .I(\this_ppu.un3_sprites_addr_cry_0_c_RNIRLAZ0Z8 ));
    CascadeMux I__4128 (
            .O(N__20940),
            .I(N__20937));
    InMux I__4127 (
            .O(N__20937),
            .I(N__20934));
    LocalMux I__4126 (
            .O(N__20934),
            .I(N__20930));
    InMux I__4125 (
            .O(N__20933),
            .I(N__20927));
    Span4Mux_v I__4124 (
            .O(N__20930),
            .I(N__20923));
    LocalMux I__4123 (
            .O(N__20927),
            .I(N__20920));
    CascadeMux I__4122 (
            .O(N__20926),
            .I(N__20917));
    Span4Mux_h I__4121 (
            .O(N__20923),
            .I(N__20914));
    Span12Mux_h I__4120 (
            .O(N__20920),
            .I(N__20907));
    InMux I__4119 (
            .O(N__20917),
            .I(N__20904));
    Span4Mux_v I__4118 (
            .O(N__20914),
            .I(N__20901));
    InMux I__4117 (
            .O(N__20913),
            .I(N__20894));
    InMux I__4116 (
            .O(N__20912),
            .I(N__20894));
    InMux I__4115 (
            .O(N__20911),
            .I(N__20894));
    InMux I__4114 (
            .O(N__20910),
            .I(N__20891));
    Span12Mux_v I__4113 (
            .O(N__20907),
            .I(N__20886));
    LocalMux I__4112 (
            .O(N__20904),
            .I(N__20886));
    Odrv4 I__4111 (
            .O(N__20901),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__4110 (
            .O(N__20894),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__4109 (
            .O(N__20891),
            .I(M_this_ppu_vram_addr_1));
    Odrv12 I__4108 (
            .O(N__20886),
            .I(M_this_ppu_vram_addr_1));
    CascadeMux I__4107 (
            .O(N__20877),
            .I(N__20874));
    CascadeBuf I__4106 (
            .O(N__20874),
            .I(N__20871));
    CascadeMux I__4105 (
            .O(N__20871),
            .I(N__20868));
    CascadeBuf I__4104 (
            .O(N__20868),
            .I(N__20865));
    CascadeMux I__4103 (
            .O(N__20865),
            .I(N__20862));
    CascadeBuf I__4102 (
            .O(N__20862),
            .I(N__20859));
    CascadeMux I__4101 (
            .O(N__20859),
            .I(N__20856));
    CascadeBuf I__4100 (
            .O(N__20856),
            .I(N__20853));
    CascadeMux I__4099 (
            .O(N__20853),
            .I(N__20850));
    CascadeBuf I__4098 (
            .O(N__20850),
            .I(N__20847));
    CascadeMux I__4097 (
            .O(N__20847),
            .I(N__20844));
    CascadeBuf I__4096 (
            .O(N__20844),
            .I(N__20841));
    CascadeMux I__4095 (
            .O(N__20841),
            .I(N__20838));
    CascadeBuf I__4094 (
            .O(N__20838),
            .I(N__20835));
    CascadeMux I__4093 (
            .O(N__20835),
            .I(N__20832));
    CascadeBuf I__4092 (
            .O(N__20832),
            .I(N__20829));
    CascadeMux I__4091 (
            .O(N__20829),
            .I(N__20826));
    CascadeBuf I__4090 (
            .O(N__20826),
            .I(N__20823));
    CascadeMux I__4089 (
            .O(N__20823),
            .I(N__20820));
    CascadeBuf I__4088 (
            .O(N__20820),
            .I(N__20817));
    CascadeMux I__4087 (
            .O(N__20817),
            .I(N__20814));
    CascadeBuf I__4086 (
            .O(N__20814),
            .I(N__20811));
    CascadeMux I__4085 (
            .O(N__20811),
            .I(N__20808));
    CascadeBuf I__4084 (
            .O(N__20808),
            .I(N__20805));
    CascadeMux I__4083 (
            .O(N__20805),
            .I(N__20802));
    CascadeBuf I__4082 (
            .O(N__20802),
            .I(N__20799));
    CascadeMux I__4081 (
            .O(N__20799),
            .I(N__20796));
    CascadeBuf I__4080 (
            .O(N__20796),
            .I(N__20793));
    CascadeMux I__4079 (
            .O(N__20793),
            .I(N__20790));
    CascadeBuf I__4078 (
            .O(N__20790),
            .I(N__20787));
    CascadeMux I__4077 (
            .O(N__20787),
            .I(N__20784));
    InMux I__4076 (
            .O(N__20784),
            .I(N__20781));
    LocalMux I__4075 (
            .O(N__20781),
            .I(N__20778));
    Odrv12 I__4074 (
            .O(N__20778),
            .I(M_this_ppu_sprites_addr_1));
    InMux I__4073 (
            .O(N__20775),
            .I(N__20772));
    LocalMux I__4072 (
            .O(N__20772),
            .I(N__20769));
    Span4Mux_h I__4071 (
            .O(N__20769),
            .I(N__20766));
    Span4Mux_v I__4070 (
            .O(N__20766),
            .I(N__20763));
    Odrv4 I__4069 (
            .O(N__20763),
            .I(\this_sprites_ram.mem_out_bus4_1 ));
    InMux I__4068 (
            .O(N__20760),
            .I(N__20757));
    LocalMux I__4067 (
            .O(N__20757),
            .I(N__20754));
    Span4Mux_v I__4066 (
            .O(N__20754),
            .I(N__20751));
    Span4Mux_h I__4065 (
            .O(N__20751),
            .I(N__20748));
    Span4Mux_v I__4064 (
            .O(N__20748),
            .I(N__20745));
    Odrv4 I__4063 (
            .O(N__20745),
            .I(\this_sprites_ram.mem_out_bus0_1 ));
    InMux I__4062 (
            .O(N__20742),
            .I(N__20738));
    CascadeMux I__4061 (
            .O(N__20741),
            .I(N__20735));
    LocalMux I__4060 (
            .O(N__20738),
            .I(N__20732));
    InMux I__4059 (
            .O(N__20735),
            .I(N__20726));
    Span4Mux_h I__4058 (
            .O(N__20732),
            .I(N__20723));
    InMux I__4057 (
            .O(N__20731),
            .I(N__20716));
    InMux I__4056 (
            .O(N__20730),
            .I(N__20716));
    InMux I__4055 (
            .O(N__20729),
            .I(N__20716));
    LocalMux I__4054 (
            .O(N__20726),
            .I(M_this_state_qZ0Z_12));
    Odrv4 I__4053 (
            .O(N__20723),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__4052 (
            .O(N__20716),
            .I(M_this_state_qZ0Z_12));
    CascadeMux I__4051 (
            .O(N__20709),
            .I(N__20706));
    InMux I__4050 (
            .O(N__20706),
            .I(N__20703));
    LocalMux I__4049 (
            .O(N__20703),
            .I(\this_start_data_delay.N_125 ));
    CascadeMux I__4048 (
            .O(N__20700),
            .I(\this_start_data_delay.un30_0_0_cascade_ ));
    InMux I__4047 (
            .O(N__20697),
            .I(N__20694));
    LocalMux I__4046 (
            .O(N__20694),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_3_x1 ));
    InMux I__4045 (
            .O(N__20691),
            .I(N__20688));
    LocalMux I__4044 (
            .O(N__20688),
            .I(N__20684));
    InMux I__4043 (
            .O(N__20687),
            .I(N__20681));
    Span4Mux_h I__4042 (
            .O(N__20684),
            .I(N__20678));
    LocalMux I__4041 (
            .O(N__20681),
            .I(N__20675));
    Odrv4 I__4040 (
            .O(N__20678),
            .I(\this_vga_signals.N_4_0 ));
    Odrv4 I__4039 (
            .O(N__20675),
            .I(\this_vga_signals.N_4_0 ));
    CascadeMux I__4038 (
            .O(N__20670),
            .I(\this_vga_signals.g0_6_1_cascade_ ));
    InMux I__4037 (
            .O(N__20667),
            .I(N__20663));
    InMux I__4036 (
            .O(N__20666),
            .I(N__20657));
    LocalMux I__4035 (
            .O(N__20663),
            .I(N__20648));
    InMux I__4034 (
            .O(N__20662),
            .I(N__20645));
    InMux I__4033 (
            .O(N__20661),
            .I(N__20640));
    InMux I__4032 (
            .O(N__20660),
            .I(N__20640));
    LocalMux I__4031 (
            .O(N__20657),
            .I(N__20637));
    InMux I__4030 (
            .O(N__20656),
            .I(N__20632));
    InMux I__4029 (
            .O(N__20655),
            .I(N__20632));
    InMux I__4028 (
            .O(N__20654),
            .I(N__20623));
    InMux I__4027 (
            .O(N__20653),
            .I(N__20623));
    InMux I__4026 (
            .O(N__20652),
            .I(N__20623));
    InMux I__4025 (
            .O(N__20651),
            .I(N__20623));
    Odrv4 I__4024 (
            .O(N__20648),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__4023 (
            .O(N__20645),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__4022 (
            .O(N__20640),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    Odrv12 I__4021 (
            .O(N__20637),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__4020 (
            .O(N__20632),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__4019 (
            .O(N__20623),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    InMux I__4018 (
            .O(N__20610),
            .I(N__20607));
    LocalMux I__4017 (
            .O(N__20607),
            .I(N__20604));
    Odrv4 I__4016 (
            .O(N__20604),
            .I(\this_vga_signals.N_4_0_0_1 ));
    InMux I__4015 (
            .O(N__20601),
            .I(N__20598));
    LocalMux I__4014 (
            .O(N__20598),
            .I(N__20595));
    Odrv4 I__4013 (
            .O(N__20595),
            .I(\this_vga_signals.vaddress_0_5 ));
    CascadeMux I__4012 (
            .O(N__20592),
            .I(\this_vga_signals.vaddress_0_6_cascade_ ));
    InMux I__4011 (
            .O(N__20589),
            .I(N__20586));
    LocalMux I__4010 (
            .O(N__20586),
            .I(N__20583));
    Odrv4 I__4009 (
            .O(N__20583),
            .I(\this_vga_signals.mult1_un47_sum_c3_0 ));
    InMux I__4008 (
            .O(N__20580),
            .I(N__20576));
    CascadeMux I__4007 (
            .O(N__20579),
            .I(N__20573));
    LocalMux I__4006 (
            .O(N__20576),
            .I(N__20566));
    InMux I__4005 (
            .O(N__20573),
            .I(N__20560));
    InMux I__4004 (
            .O(N__20572),
            .I(N__20560));
    InMux I__4003 (
            .O(N__20571),
            .I(N__20553));
    InMux I__4002 (
            .O(N__20570),
            .I(N__20553));
    InMux I__4001 (
            .O(N__20569),
            .I(N__20553));
    Span4Mux_h I__4000 (
            .O(N__20566),
            .I(N__20548));
    InMux I__3999 (
            .O(N__20565),
            .I(N__20545));
    LocalMux I__3998 (
            .O(N__20560),
            .I(N__20542));
    LocalMux I__3997 (
            .O(N__20553),
            .I(N__20539));
    InMux I__3996 (
            .O(N__20552),
            .I(N__20536));
    InMux I__3995 (
            .O(N__20551),
            .I(N__20533));
    Odrv4 I__3994 (
            .O(N__20548),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__3993 (
            .O(N__20545),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__3992 (
            .O(N__20542),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__3991 (
            .O(N__20539),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__3990 (
            .O(N__20536),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__3989 (
            .O(N__20533),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    InMux I__3988 (
            .O(N__20520),
            .I(N__20515));
    CascadeMux I__3987 (
            .O(N__20519),
            .I(N__20510));
    InMux I__3986 (
            .O(N__20518),
            .I(N__20505));
    LocalMux I__3985 (
            .O(N__20515),
            .I(N__20499));
    InMux I__3984 (
            .O(N__20514),
            .I(N__20496));
    InMux I__3983 (
            .O(N__20513),
            .I(N__20489));
    InMux I__3982 (
            .O(N__20510),
            .I(N__20489));
    InMux I__3981 (
            .O(N__20509),
            .I(N__20489));
    InMux I__3980 (
            .O(N__20508),
            .I(N__20486));
    LocalMux I__3979 (
            .O(N__20505),
            .I(N__20483));
    InMux I__3978 (
            .O(N__20504),
            .I(N__20478));
    InMux I__3977 (
            .O(N__20503),
            .I(N__20478));
    InMux I__3976 (
            .O(N__20502),
            .I(N__20475));
    Span4Mux_h I__3975 (
            .O(N__20499),
            .I(N__20466));
    LocalMux I__3974 (
            .O(N__20496),
            .I(N__20466));
    LocalMux I__3973 (
            .O(N__20489),
            .I(N__20466));
    LocalMux I__3972 (
            .O(N__20486),
            .I(N__20466));
    Odrv12 I__3971 (
            .O(N__20483),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__3970 (
            .O(N__20478),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__3969 (
            .O(N__20475),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__3968 (
            .O(N__20466),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    CascadeMux I__3967 (
            .O(N__20457),
            .I(N__20451));
    CascadeMux I__3966 (
            .O(N__20456),
            .I(N__20447));
    CascadeMux I__3965 (
            .O(N__20455),
            .I(N__20444));
    InMux I__3964 (
            .O(N__20454),
            .I(N__20439));
    InMux I__3963 (
            .O(N__20451),
            .I(N__20439));
    InMux I__3962 (
            .O(N__20450),
            .I(N__20436));
    InMux I__3961 (
            .O(N__20447),
            .I(N__20431));
    InMux I__3960 (
            .O(N__20444),
            .I(N__20431));
    LocalMux I__3959 (
            .O(N__20439),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__3958 (
            .O(N__20436),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__3957 (
            .O(N__20431),
            .I(\this_vga_signals.vaddress_5 ));
    InMux I__3956 (
            .O(N__20424),
            .I(N__20420));
    InMux I__3955 (
            .O(N__20423),
            .I(N__20415));
    LocalMux I__3954 (
            .O(N__20420),
            .I(N__20406));
    InMux I__3953 (
            .O(N__20419),
            .I(N__20401));
    InMux I__3952 (
            .O(N__20418),
            .I(N__20401));
    LocalMux I__3951 (
            .O(N__20415),
            .I(N__20398));
    InMux I__3950 (
            .O(N__20414),
            .I(N__20393));
    InMux I__3949 (
            .O(N__20413),
            .I(N__20393));
    InMux I__3948 (
            .O(N__20412),
            .I(N__20384));
    InMux I__3947 (
            .O(N__20411),
            .I(N__20384));
    InMux I__3946 (
            .O(N__20410),
            .I(N__20384));
    InMux I__3945 (
            .O(N__20409),
            .I(N__20384));
    Odrv4 I__3944 (
            .O(N__20406),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__3943 (
            .O(N__20401),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__3942 (
            .O(N__20398),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__3941 (
            .O(N__20393),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__3940 (
            .O(N__20384),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    CascadeMux I__3939 (
            .O(N__20373),
            .I(N__20367));
    InMux I__3938 (
            .O(N__20372),
            .I(N__20363));
    InMux I__3937 (
            .O(N__20371),
            .I(N__20360));
    InMux I__3936 (
            .O(N__20370),
            .I(N__20355));
    InMux I__3935 (
            .O(N__20367),
            .I(N__20355));
    InMux I__3934 (
            .O(N__20366),
            .I(N__20352));
    LocalMux I__3933 (
            .O(N__20363),
            .I(N__20348));
    LocalMux I__3932 (
            .O(N__20360),
            .I(N__20343));
    LocalMux I__3931 (
            .O(N__20355),
            .I(N__20343));
    LocalMux I__3930 (
            .O(N__20352),
            .I(N__20338));
    InMux I__3929 (
            .O(N__20351),
            .I(N__20335));
    Span4Mux_v I__3928 (
            .O(N__20348),
            .I(N__20328));
    Span4Mux_v I__3927 (
            .O(N__20343),
            .I(N__20328));
    InMux I__3926 (
            .O(N__20342),
            .I(N__20323));
    InMux I__3925 (
            .O(N__20341),
            .I(N__20323));
    Span4Mux_h I__3924 (
            .O(N__20338),
            .I(N__20320));
    LocalMux I__3923 (
            .O(N__20335),
            .I(N__20317));
    InMux I__3922 (
            .O(N__20334),
            .I(N__20312));
    InMux I__3921 (
            .O(N__20333),
            .I(N__20312));
    Odrv4 I__3920 (
            .O(N__20328),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__3919 (
            .O(N__20323),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__3918 (
            .O(N__20320),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__3917 (
            .O(N__20317),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__3916 (
            .O(N__20312),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    CascadeMux I__3915 (
            .O(N__20301),
            .I(\this_vga_signals.g2_1_cascade_ ));
    InMux I__3914 (
            .O(N__20298),
            .I(N__20294));
    InMux I__3913 (
            .O(N__20297),
            .I(N__20291));
    LocalMux I__3912 (
            .O(N__20294),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_2 ));
    LocalMux I__3911 (
            .O(N__20291),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_2 ));
    InMux I__3910 (
            .O(N__20286),
            .I(N__20283));
    LocalMux I__3909 (
            .O(N__20283),
            .I(N__20280));
    Span4Mux_h I__3908 (
            .O(N__20280),
            .I(N__20277));
    Odrv4 I__3907 (
            .O(N__20277),
            .I(\this_vga_signals.g0_i_x4_0_0 ));
    CascadeMux I__3906 (
            .O(N__20274),
            .I(N__20271));
    InMux I__3905 (
            .O(N__20271),
            .I(N__20268));
    LocalMux I__3904 (
            .O(N__20268),
            .I(N__20265));
    Odrv12 I__3903 (
            .O(N__20265),
            .I(\this_vga_signals.g0_3_0_a3_1 ));
    InMux I__3902 (
            .O(N__20262),
            .I(N__20259));
    LocalMux I__3901 (
            .O(N__20259),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_602_x0 ));
    InMux I__3900 (
            .O(N__20256),
            .I(N__20252));
    InMux I__3899 (
            .O(N__20255),
            .I(N__20249));
    LocalMux I__3898 (
            .O(N__20252),
            .I(N__20240));
    LocalMux I__3897 (
            .O(N__20249),
            .I(N__20240));
    InMux I__3896 (
            .O(N__20248),
            .I(N__20234));
    CascadeMux I__3895 (
            .O(N__20247),
            .I(N__20230));
    InMux I__3894 (
            .O(N__20246),
            .I(N__20227));
    InMux I__3893 (
            .O(N__20245),
            .I(N__20224));
    Span4Mux_v I__3892 (
            .O(N__20240),
            .I(N__20221));
    InMux I__3891 (
            .O(N__20239),
            .I(N__20216));
    InMux I__3890 (
            .O(N__20238),
            .I(N__20216));
    InMux I__3889 (
            .O(N__20237),
            .I(N__20213));
    LocalMux I__3888 (
            .O(N__20234),
            .I(N__20210));
    InMux I__3887 (
            .O(N__20233),
            .I(N__20205));
    InMux I__3886 (
            .O(N__20230),
            .I(N__20205));
    LocalMux I__3885 (
            .O(N__20227),
            .I(N__20202));
    LocalMux I__3884 (
            .O(N__20224),
            .I(\this_vga_signals.vaddress_c2 ));
    Odrv4 I__3883 (
            .O(N__20221),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__3882 (
            .O(N__20216),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__3881 (
            .O(N__20213),
            .I(\this_vga_signals.vaddress_c2 ));
    Odrv4 I__3880 (
            .O(N__20210),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__3879 (
            .O(N__20205),
            .I(\this_vga_signals.vaddress_c2 ));
    Odrv4 I__3878 (
            .O(N__20202),
            .I(\this_vga_signals.vaddress_c2 ));
    CascadeMux I__3877 (
            .O(N__20187),
            .I(N__20184));
    InMux I__3876 (
            .O(N__20184),
            .I(N__20180));
    CascadeMux I__3875 (
            .O(N__20183),
            .I(N__20177));
    LocalMux I__3874 (
            .O(N__20180),
            .I(N__20174));
    InMux I__3873 (
            .O(N__20177),
            .I(N__20171));
    Span4Mux_v I__3872 (
            .O(N__20174),
            .I(N__20168));
    LocalMux I__3871 (
            .O(N__20171),
            .I(N__20165));
    Span4Mux_h I__3870 (
            .O(N__20168),
            .I(N__20162));
    Span4Mux_v I__3869 (
            .O(N__20165),
            .I(N__20159));
    Odrv4 I__3868 (
            .O(N__20162),
            .I(\this_vga_signals.r_N_4_mux ));
    Odrv4 I__3867 (
            .O(N__20159),
            .I(\this_vga_signals.r_N_4_mux ));
    CascadeMux I__3866 (
            .O(N__20154),
            .I(\this_vga_signals.r_N_4_mux_cascade_ ));
    InMux I__3865 (
            .O(N__20151),
            .I(N__20148));
    LocalMux I__3864 (
            .O(N__20148),
            .I(N__20144));
    CascadeMux I__3863 (
            .O(N__20147),
            .I(N__20141));
    Span4Mux_v I__3862 (
            .O(N__20144),
            .I(N__20138));
    InMux I__3861 (
            .O(N__20141),
            .I(N__20135));
    Odrv4 I__3860 (
            .O(N__20138),
            .I(\this_vga_signals.SUM_2 ));
    LocalMux I__3859 (
            .O(N__20135),
            .I(\this_vga_signals.SUM_2 ));
    CascadeMux I__3858 (
            .O(N__20130),
            .I(N__20127));
    InMux I__3857 (
            .O(N__20127),
            .I(N__20121));
    InMux I__3856 (
            .O(N__20126),
            .I(N__20118));
    InMux I__3855 (
            .O(N__20125),
            .I(N__20113));
    InMux I__3854 (
            .O(N__20124),
            .I(N__20113));
    LocalMux I__3853 (
            .O(N__20121),
            .I(N__20110));
    LocalMux I__3852 (
            .O(N__20118),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__3851 (
            .O(N__20113),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    Odrv4 I__3850 (
            .O(N__20110),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    CascadeMux I__3849 (
            .O(N__20103),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x1_cascade_ ));
    InMux I__3848 (
            .O(N__20100),
            .I(N__20097));
    LocalMux I__3847 (
            .O(N__20097),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a1_ns ));
    InMux I__3846 (
            .O(N__20094),
            .I(N__20091));
    LocalMux I__3845 (
            .O(N__20091),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x0 ));
    CascadeMux I__3844 (
            .O(N__20088),
            .I(N__20080));
    InMux I__3843 (
            .O(N__20087),
            .I(N__20077));
    CascadeMux I__3842 (
            .O(N__20086),
            .I(N__20074));
    CascadeMux I__3841 (
            .O(N__20085),
            .I(N__20067));
    InMux I__3840 (
            .O(N__20084),
            .I(N__20064));
    InMux I__3839 (
            .O(N__20083),
            .I(N__20059));
    InMux I__3838 (
            .O(N__20080),
            .I(N__20059));
    LocalMux I__3837 (
            .O(N__20077),
            .I(N__20056));
    InMux I__3836 (
            .O(N__20074),
            .I(N__20049));
    InMux I__3835 (
            .O(N__20073),
            .I(N__20049));
    InMux I__3834 (
            .O(N__20072),
            .I(N__20049));
    InMux I__3833 (
            .O(N__20071),
            .I(N__20044));
    InMux I__3832 (
            .O(N__20070),
            .I(N__20044));
    InMux I__3831 (
            .O(N__20067),
            .I(N__20041));
    LocalMux I__3830 (
            .O(N__20064),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__3829 (
            .O(N__20059),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    Odrv4 I__3828 (
            .O(N__20056),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__3827 (
            .O(N__20049),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__3826 (
            .O(N__20044),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__3825 (
            .O(N__20041),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    InMux I__3824 (
            .O(N__20028),
            .I(N__20022));
    InMux I__3823 (
            .O(N__20027),
            .I(N__20015));
    InMux I__3822 (
            .O(N__20026),
            .I(N__20015));
    InMux I__3821 (
            .O(N__20025),
            .I(N__20015));
    LocalMux I__3820 (
            .O(N__20022),
            .I(N__20012));
    LocalMux I__3819 (
            .O(N__20015),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    Odrv4 I__3818 (
            .O(N__20012),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    CascadeMux I__3817 (
            .O(N__20007),
            .I(N__20004));
    InMux I__3816 (
            .O(N__20004),
            .I(N__20001));
    LocalMux I__3815 (
            .O(N__20001),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_602_x1 ));
    InMux I__3814 (
            .O(N__19998),
            .I(N__19995));
    LocalMux I__3813 (
            .O(N__19995),
            .I(\this_start_data_delay.N_67 ));
    InMux I__3812 (
            .O(N__19992),
            .I(N__19989));
    LocalMux I__3811 (
            .O(N__19989),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_2_1_0 ));
    InMux I__3810 (
            .O(N__19986),
            .I(N__19983));
    LocalMux I__3809 (
            .O(N__19983),
            .I(\this_vga_signals.N_4558_0 ));
    CascadeMux I__3808 (
            .O(N__19980),
            .I(\this_vga_signals.g0_4_i_a3_1_cascade_ ));
    CascadeMux I__3807 (
            .O(N__19977),
            .I(\this_vga_signals.g0_4_i_1_cascade_ ));
    InMux I__3806 (
            .O(N__19974),
            .I(N__19971));
    LocalMux I__3805 (
            .O(N__19971),
            .I(\this_vga_signals.N_6_2 ));
    InMux I__3804 (
            .O(N__19968),
            .I(N__19964));
    InMux I__3803 (
            .O(N__19967),
            .I(N__19961));
    LocalMux I__3802 (
            .O(N__19964),
            .I(\this_start_data_delay.N_47_0 ));
    LocalMux I__3801 (
            .O(N__19961),
            .I(\this_start_data_delay.N_47_0 ));
    CascadeMux I__3800 (
            .O(N__19956),
            .I(\this_start_data_delay.N_909_0_cascade_ ));
    IoInMux I__3799 (
            .O(N__19953),
            .I(N__19950));
    LocalMux I__3798 (
            .O(N__19950),
            .I(N__19947));
    IoSpan4Mux I__3797 (
            .O(N__19947),
            .I(N__19944));
    Span4Mux_s0_h I__3796 (
            .O(N__19944),
            .I(N__19941));
    Span4Mux_v I__3795 (
            .O(N__19941),
            .I(N__19938));
    Sp12to4 I__3794 (
            .O(N__19938),
            .I(N__19935));
    Span12Mux_h I__3793 (
            .O(N__19935),
            .I(N__19929));
    InMux I__3792 (
            .O(N__19934),
            .I(N__19926));
    InMux I__3791 (
            .O(N__19933),
            .I(N__19921));
    InMux I__3790 (
            .O(N__19932),
            .I(N__19921));
    Odrv12 I__3789 (
            .O(N__19929),
            .I(led_c_1));
    LocalMux I__3788 (
            .O(N__19926),
            .I(led_c_1));
    LocalMux I__3787 (
            .O(N__19921),
            .I(led_c_1));
    InMux I__3786 (
            .O(N__19914),
            .I(N__19911));
    LocalMux I__3785 (
            .O(N__19911),
            .I(N__19908));
    Odrv4 I__3784 (
            .O(N__19908),
            .I(\this_start_data_delay.M_this_state_q_ns_0_i_0_0 ));
    InMux I__3783 (
            .O(N__19905),
            .I(N__19902));
    LocalMux I__3782 (
            .O(N__19902),
            .I(\this_start_data_delay.M_this_state_q_ns_0_i_2_0_0 ));
    CEMux I__3781 (
            .O(N__19899),
            .I(N__19893));
    CEMux I__3780 (
            .O(N__19898),
            .I(N__19888));
    InMux I__3779 (
            .O(N__19897),
            .I(N__19884));
    CascadeMux I__3778 (
            .O(N__19896),
            .I(N__19880));
    LocalMux I__3777 (
            .O(N__19893),
            .I(N__19877));
    InMux I__3776 (
            .O(N__19892),
            .I(N__19873));
    InMux I__3775 (
            .O(N__19891),
            .I(N__19869));
    LocalMux I__3774 (
            .O(N__19888),
            .I(N__19865));
    InMux I__3773 (
            .O(N__19887),
            .I(N__19862));
    LocalMux I__3772 (
            .O(N__19884),
            .I(N__19859));
    InMux I__3771 (
            .O(N__19883),
            .I(N__19856));
    InMux I__3770 (
            .O(N__19880),
            .I(N__19853));
    Span4Mux_h I__3769 (
            .O(N__19877),
            .I(N__19850));
    InMux I__3768 (
            .O(N__19876),
            .I(N__19847));
    LocalMux I__3767 (
            .O(N__19873),
            .I(N__19844));
    InMux I__3766 (
            .O(N__19872),
            .I(N__19841));
    LocalMux I__3765 (
            .O(N__19869),
            .I(N__19838));
    InMux I__3764 (
            .O(N__19868),
            .I(N__19835));
    Span4Mux_h I__3763 (
            .O(N__19865),
            .I(N__19824));
    LocalMux I__3762 (
            .O(N__19862),
            .I(N__19824));
    Span4Mux_v I__3761 (
            .O(N__19859),
            .I(N__19824));
    LocalMux I__3760 (
            .O(N__19856),
            .I(N__19824));
    LocalMux I__3759 (
            .O(N__19853),
            .I(N__19824));
    Span4Mux_v I__3758 (
            .O(N__19850),
            .I(N__19818));
    LocalMux I__3757 (
            .O(N__19847),
            .I(N__19818));
    Span4Mux_h I__3756 (
            .O(N__19844),
            .I(N__19813));
    LocalMux I__3755 (
            .O(N__19841),
            .I(N__19813));
    Span4Mux_h I__3754 (
            .O(N__19838),
            .I(N__19806));
    LocalMux I__3753 (
            .O(N__19835),
            .I(N__19806));
    Span4Mux_v I__3752 (
            .O(N__19824),
            .I(N__19806));
    InMux I__3751 (
            .O(N__19823),
            .I(N__19803));
    Span4Mux_h I__3750 (
            .O(N__19818),
            .I(N__19800));
    Span4Mux_v I__3749 (
            .O(N__19813),
            .I(N__19795));
    Span4Mux_h I__3748 (
            .O(N__19806),
            .I(N__19795));
    LocalMux I__3747 (
            .O(N__19803),
            .I(N__19791));
    Span4Mux_h I__3746 (
            .O(N__19800),
            .I(N__19788));
    Span4Mux_h I__3745 (
            .O(N__19795),
            .I(N__19785));
    InMux I__3744 (
            .O(N__19794),
            .I(N__19782));
    Span12Mux_h I__3743 (
            .O(N__19791),
            .I(N__19777));
    Sp12to4 I__3742 (
            .O(N__19788),
            .I(N__19777));
    Span4Mux_v I__3741 (
            .O(N__19785),
            .I(N__19774));
    LocalMux I__3740 (
            .O(N__19782),
            .I(N_822_0));
    Odrv12 I__3739 (
            .O(N__19777),
            .I(N_822_0));
    Odrv4 I__3738 (
            .O(N__19774),
            .I(N_822_0));
    CascadeMux I__3737 (
            .O(N__19767),
            .I(\this_start_data_delay.N_910_cascade_ ));
    InMux I__3736 (
            .O(N__19764),
            .I(N__19760));
    InMux I__3735 (
            .O(N__19763),
            .I(N__19757));
    LocalMux I__3734 (
            .O(N__19760),
            .I(N__19749));
    LocalMux I__3733 (
            .O(N__19757),
            .I(N__19749));
    InMux I__3732 (
            .O(N__19756),
            .I(N__19746));
    InMux I__3731 (
            .O(N__19755),
            .I(N__19743));
    InMux I__3730 (
            .O(N__19754),
            .I(N__19740));
    Odrv4 I__3729 (
            .O(N__19749),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__3728 (
            .O(N__19746),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__3727 (
            .O(N__19743),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__3726 (
            .O(N__19740),
            .I(M_this_state_qZ0Z_10));
    CascadeMux I__3725 (
            .O(N__19731),
            .I(N__19728));
    InMux I__3724 (
            .O(N__19728),
            .I(N__19724));
    InMux I__3723 (
            .O(N__19727),
            .I(N__19720));
    LocalMux I__3722 (
            .O(N__19724),
            .I(N__19717));
    InMux I__3721 (
            .O(N__19723),
            .I(N__19714));
    LocalMux I__3720 (
            .O(N__19720),
            .I(\this_start_data_delay.N_90_0 ));
    Odrv4 I__3719 (
            .O(N__19717),
            .I(\this_start_data_delay.N_90_0 ));
    LocalMux I__3718 (
            .O(N__19714),
            .I(\this_start_data_delay.N_90_0 ));
    CascadeMux I__3717 (
            .O(N__19707),
            .I(N__19700));
    CascadeMux I__3716 (
            .O(N__19706),
            .I(N__19697));
    CascadeMux I__3715 (
            .O(N__19705),
            .I(N__19693));
    InMux I__3714 (
            .O(N__19704),
            .I(N__19688));
    InMux I__3713 (
            .O(N__19703),
            .I(N__19688));
    InMux I__3712 (
            .O(N__19700),
            .I(N__19681));
    InMux I__3711 (
            .O(N__19697),
            .I(N__19681));
    InMux I__3710 (
            .O(N__19696),
            .I(N__19678));
    InMux I__3709 (
            .O(N__19693),
            .I(N__19675));
    LocalMux I__3708 (
            .O(N__19688),
            .I(N__19672));
    InMux I__3707 (
            .O(N__19687),
            .I(N__19667));
    InMux I__3706 (
            .O(N__19686),
            .I(N__19667));
    LocalMux I__3705 (
            .O(N__19681),
            .I(N__19662));
    LocalMux I__3704 (
            .O(N__19678),
            .I(N__19662));
    LocalMux I__3703 (
            .O(N__19675),
            .I(N__19655));
    Span4Mux_v I__3702 (
            .O(N__19672),
            .I(N__19655));
    LocalMux I__3701 (
            .O(N__19667),
            .I(N__19655));
    Span4Mux_v I__3700 (
            .O(N__19662),
            .I(N__19652));
    Span4Mux_h I__3699 (
            .O(N__19655),
            .I(N__19649));
    Span4Mux_v I__3698 (
            .O(N__19652),
            .I(N__19646));
    Span4Mux_h I__3697 (
            .O(N__19649),
            .I(N__19643));
    Sp12to4 I__3696 (
            .O(N__19646),
            .I(N__19640));
    Sp12to4 I__3695 (
            .O(N__19643),
            .I(N__19637));
    Span12Mux_h I__3694 (
            .O(N__19640),
            .I(N__19634));
    Odrv12 I__3693 (
            .O(N__19637),
            .I(port_address_in_1));
    Odrv12 I__3692 (
            .O(N__19634),
            .I(port_address_in_1));
    InMux I__3691 (
            .O(N__19629),
            .I(N__19621));
    InMux I__3690 (
            .O(N__19628),
            .I(N__19616));
    InMux I__3689 (
            .O(N__19627),
            .I(N__19611));
    InMux I__3688 (
            .O(N__19626),
            .I(N__19611));
    InMux I__3687 (
            .O(N__19625),
            .I(N__19606));
    InMux I__3686 (
            .O(N__19624),
            .I(N__19606));
    LocalMux I__3685 (
            .O(N__19621),
            .I(N__19603));
    InMux I__3684 (
            .O(N__19620),
            .I(N__19598));
    InMux I__3683 (
            .O(N__19619),
            .I(N__19598));
    LocalMux I__3682 (
            .O(N__19616),
            .I(N__19593));
    LocalMux I__3681 (
            .O(N__19611),
            .I(N__19593));
    LocalMux I__3680 (
            .O(N__19606),
            .I(N__19586));
    Span4Mux_v I__3679 (
            .O(N__19603),
            .I(N__19586));
    LocalMux I__3678 (
            .O(N__19598),
            .I(N__19586));
    Span4Mux_v I__3677 (
            .O(N__19593),
            .I(N__19583));
    Span4Mux_h I__3676 (
            .O(N__19586),
            .I(N__19580));
    Sp12to4 I__3675 (
            .O(N__19583),
            .I(N__19577));
    Sp12to4 I__3674 (
            .O(N__19580),
            .I(N__19572));
    Span12Mux_h I__3673 (
            .O(N__19577),
            .I(N__19572));
    Odrv12 I__3672 (
            .O(N__19572),
            .I(port_address_in_0));
    CascadeMux I__3671 (
            .O(N__19569),
            .I(N__19564));
    CascadeMux I__3670 (
            .O(N__19568),
            .I(N__19561));
    CascadeMux I__3669 (
            .O(N__19567),
            .I(N__19556));
    InMux I__3668 (
            .O(N__19564),
            .I(N__19551));
    InMux I__3667 (
            .O(N__19561),
            .I(N__19551));
    InMux I__3666 (
            .O(N__19560),
            .I(N__19544));
    InMux I__3665 (
            .O(N__19559),
            .I(N__19544));
    InMux I__3664 (
            .O(N__19556),
            .I(N__19541));
    LocalMux I__3663 (
            .O(N__19551),
            .I(N__19538));
    InMux I__3662 (
            .O(N__19550),
            .I(N__19533));
    InMux I__3661 (
            .O(N__19549),
            .I(N__19533));
    LocalMux I__3660 (
            .O(N__19544),
            .I(N__19530));
    LocalMux I__3659 (
            .O(N__19541),
            .I(N__19527));
    Span4Mux_v I__3658 (
            .O(N__19538),
            .I(N__19522));
    LocalMux I__3657 (
            .O(N__19533),
            .I(N__19522));
    Span4Mux_v I__3656 (
            .O(N__19530),
            .I(N__19519));
    Span4Mux_v I__3655 (
            .O(N__19527),
            .I(N__19516));
    Span4Mux_h I__3654 (
            .O(N__19522),
            .I(N__19513));
    Span4Mux_v I__3653 (
            .O(N__19519),
            .I(N__19508));
    Span4Mux_v I__3652 (
            .O(N__19516),
            .I(N__19508));
    Sp12to4 I__3651 (
            .O(N__19513),
            .I(N__19505));
    Span4Mux_v I__3650 (
            .O(N__19508),
            .I(N__19502));
    Span12Mux_v I__3649 (
            .O(N__19505),
            .I(N__19499));
    IoSpan4Mux I__3648 (
            .O(N__19502),
            .I(N__19496));
    Odrv12 I__3647 (
            .O(N__19499),
            .I(port_address_in_2));
    Odrv4 I__3646 (
            .O(N__19496),
            .I(port_address_in_2));
    InMux I__3645 (
            .O(N__19491),
            .I(N__19483));
    InMux I__3644 (
            .O(N__19490),
            .I(N__19483));
    InMux I__3643 (
            .O(N__19489),
            .I(N__19480));
    InMux I__3642 (
            .O(N__19488),
            .I(N__19477));
    LocalMux I__3641 (
            .O(N__19483),
            .I(\this_start_data_delay.N_48_0 ));
    LocalMux I__3640 (
            .O(N__19480),
            .I(\this_start_data_delay.N_48_0 ));
    LocalMux I__3639 (
            .O(N__19477),
            .I(\this_start_data_delay.N_48_0 ));
    CascadeMux I__3638 (
            .O(N__19470),
            .I(N__19467));
    InMux I__3637 (
            .O(N__19467),
            .I(N__19464));
    LocalMux I__3636 (
            .O(N__19464),
            .I(\this_start_data_delay.N_71 ));
    CascadeMux I__3635 (
            .O(N__19461),
            .I(\this_start_data_delay.N_127_cascade_ ));
    InMux I__3634 (
            .O(N__19458),
            .I(N__19452));
    InMux I__3633 (
            .O(N__19457),
            .I(N__19449));
    InMux I__3632 (
            .O(N__19456),
            .I(N__19444));
    InMux I__3631 (
            .O(N__19455),
            .I(N__19444));
    LocalMux I__3630 (
            .O(N__19452),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__3629 (
            .O(N__19449),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__3628 (
            .O(N__19444),
            .I(M_this_state_qZ0Z_11));
    CascadeMux I__3627 (
            .O(N__19437),
            .I(\this_start_data_delay.N_844_0_cascade_ ));
    CascadeMux I__3626 (
            .O(N__19434),
            .I(\this_start_data_delay.N_151_cascade_ ));
    InMux I__3625 (
            .O(N__19431),
            .I(N__19428));
    LocalMux I__3624 (
            .O(N__19428),
            .I(N__19424));
    InMux I__3623 (
            .O(N__19427),
            .I(N__19419));
    Span4Mux_v I__3622 (
            .O(N__19424),
            .I(N__19416));
    InMux I__3621 (
            .O(N__19423),
            .I(N__19411));
    InMux I__3620 (
            .O(N__19422),
            .I(N__19411));
    LocalMux I__3619 (
            .O(N__19419),
            .I(\this_start_data_delay.N_89_0 ));
    Odrv4 I__3618 (
            .O(N__19416),
            .I(\this_start_data_delay.N_89_0 ));
    LocalMux I__3617 (
            .O(N__19411),
            .I(\this_start_data_delay.N_89_0 ));
    InMux I__3616 (
            .O(N__19404),
            .I(N__19400));
    InMux I__3615 (
            .O(N__19403),
            .I(N__19396));
    LocalMux I__3614 (
            .O(N__19400),
            .I(N__19391));
    InMux I__3613 (
            .O(N__19399),
            .I(N__19387));
    LocalMux I__3612 (
            .O(N__19396),
            .I(N__19384));
    InMux I__3611 (
            .O(N__19395),
            .I(N__19381));
    InMux I__3610 (
            .O(N__19394),
            .I(N__19378));
    Span4Mux_v I__3609 (
            .O(N__19391),
            .I(N__19375));
    InMux I__3608 (
            .O(N__19390),
            .I(N__19372));
    LocalMux I__3607 (
            .O(N__19387),
            .I(N__19369));
    Span4Mux_h I__3606 (
            .O(N__19384),
            .I(N__19364));
    LocalMux I__3605 (
            .O(N__19381),
            .I(N__19364));
    LocalMux I__3604 (
            .O(N__19378),
            .I(M_this_state_qZ0Z_16));
    Odrv4 I__3603 (
            .O(N__19375),
            .I(M_this_state_qZ0Z_16));
    LocalMux I__3602 (
            .O(N__19372),
            .I(M_this_state_qZ0Z_16));
    Odrv4 I__3601 (
            .O(N__19369),
            .I(M_this_state_qZ0Z_16));
    Odrv4 I__3600 (
            .O(N__19364),
            .I(M_this_state_qZ0Z_16));
    InMux I__3599 (
            .O(N__19353),
            .I(N__19350));
    LocalMux I__3598 (
            .O(N__19350),
            .I(N__19347));
    Span4Mux_v I__3597 (
            .O(N__19347),
            .I(N__19344));
    Sp12to4 I__3596 (
            .O(N__19344),
            .I(N__19341));
    Span12Mux_h I__3595 (
            .O(N__19341),
            .I(N__19338));
    Odrv12 I__3594 (
            .O(N__19338),
            .I(\this_ppu.un3_sprites_addr_axb_0 ));
    CascadeMux I__3593 (
            .O(N__19335),
            .I(N__19331));
    InMux I__3592 (
            .O(N__19334),
            .I(N__19328));
    InMux I__3591 (
            .O(N__19331),
            .I(N__19325));
    LocalMux I__3590 (
            .O(N__19328),
            .I(N__19322));
    LocalMux I__3589 (
            .O(N__19325),
            .I(N__19319));
    Span4Mux_h I__3588 (
            .O(N__19322),
            .I(N__19315));
    Span4Mux_v I__3587 (
            .O(N__19319),
            .I(N__19312));
    CascadeMux I__3586 (
            .O(N__19318),
            .I(N__19308));
    Span4Mux_v I__3585 (
            .O(N__19315),
            .I(N__19303));
    Span4Mux_v I__3584 (
            .O(N__19312),
            .I(N__19300));
    InMux I__3583 (
            .O(N__19311),
            .I(N__19297));
    InMux I__3582 (
            .O(N__19308),
            .I(N__19294));
    CascadeMux I__3581 (
            .O(N__19307),
            .I(N__19291));
    CascadeMux I__3580 (
            .O(N__19306),
            .I(N__19287));
    Span4Mux_v I__3579 (
            .O(N__19303),
            .I(N__19282));
    Span4Mux_v I__3578 (
            .O(N__19300),
            .I(N__19275));
    LocalMux I__3577 (
            .O(N__19297),
            .I(N__19275));
    LocalMux I__3576 (
            .O(N__19294),
            .I(N__19275));
    InMux I__3575 (
            .O(N__19291),
            .I(N__19266));
    InMux I__3574 (
            .O(N__19290),
            .I(N__19266));
    InMux I__3573 (
            .O(N__19287),
            .I(N__19266));
    InMux I__3572 (
            .O(N__19286),
            .I(N__19266));
    InMux I__3571 (
            .O(N__19285),
            .I(N__19263));
    Span4Mux_v I__3570 (
            .O(N__19282),
            .I(N__19258));
    Span4Mux_h I__3569 (
            .O(N__19275),
            .I(N__19258));
    LocalMux I__3568 (
            .O(N__19266),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__3567 (
            .O(N__19263),
            .I(M_this_ppu_vram_addr_0));
    Odrv4 I__3566 (
            .O(N__19258),
            .I(M_this_ppu_vram_addr_0));
    CascadeMux I__3565 (
            .O(N__19251),
            .I(N__19248));
    CascadeBuf I__3564 (
            .O(N__19248),
            .I(N__19245));
    CascadeMux I__3563 (
            .O(N__19245),
            .I(N__19242));
    CascadeBuf I__3562 (
            .O(N__19242),
            .I(N__19239));
    CascadeMux I__3561 (
            .O(N__19239),
            .I(N__19236));
    CascadeBuf I__3560 (
            .O(N__19236),
            .I(N__19233));
    CascadeMux I__3559 (
            .O(N__19233),
            .I(N__19230));
    CascadeBuf I__3558 (
            .O(N__19230),
            .I(N__19227));
    CascadeMux I__3557 (
            .O(N__19227),
            .I(N__19224));
    CascadeBuf I__3556 (
            .O(N__19224),
            .I(N__19221));
    CascadeMux I__3555 (
            .O(N__19221),
            .I(N__19218));
    CascadeBuf I__3554 (
            .O(N__19218),
            .I(N__19215));
    CascadeMux I__3553 (
            .O(N__19215),
            .I(N__19212));
    CascadeBuf I__3552 (
            .O(N__19212),
            .I(N__19209));
    CascadeMux I__3551 (
            .O(N__19209),
            .I(N__19206));
    CascadeBuf I__3550 (
            .O(N__19206),
            .I(N__19203));
    CascadeMux I__3549 (
            .O(N__19203),
            .I(N__19200));
    CascadeBuf I__3548 (
            .O(N__19200),
            .I(N__19197));
    CascadeMux I__3547 (
            .O(N__19197),
            .I(N__19194));
    CascadeBuf I__3546 (
            .O(N__19194),
            .I(N__19191));
    CascadeMux I__3545 (
            .O(N__19191),
            .I(N__19188));
    CascadeBuf I__3544 (
            .O(N__19188),
            .I(N__19185));
    CascadeMux I__3543 (
            .O(N__19185),
            .I(N__19182));
    CascadeBuf I__3542 (
            .O(N__19182),
            .I(N__19179));
    CascadeMux I__3541 (
            .O(N__19179),
            .I(N__19176));
    CascadeBuf I__3540 (
            .O(N__19176),
            .I(N__19173));
    CascadeMux I__3539 (
            .O(N__19173),
            .I(N__19170));
    CascadeBuf I__3538 (
            .O(N__19170),
            .I(N__19167));
    CascadeMux I__3537 (
            .O(N__19167),
            .I(N__19164));
    CascadeBuf I__3536 (
            .O(N__19164),
            .I(N__19161));
    CascadeMux I__3535 (
            .O(N__19161),
            .I(N__19158));
    InMux I__3534 (
            .O(N__19158),
            .I(N__19155));
    LocalMux I__3533 (
            .O(N__19155),
            .I(N__19152));
    Span4Mux_h I__3532 (
            .O(N__19152),
            .I(N__19149));
    Odrv4 I__3531 (
            .O(N__19149),
            .I(M_this_ppu_sprites_addr_0));
    InMux I__3530 (
            .O(N__19146),
            .I(N__19141));
    CascadeMux I__3529 (
            .O(N__19145),
            .I(N__19138));
    InMux I__3528 (
            .O(N__19144),
            .I(N__19134));
    LocalMux I__3527 (
            .O(N__19141),
            .I(N__19131));
    InMux I__3526 (
            .O(N__19138),
            .I(N__19126));
    InMux I__3525 (
            .O(N__19137),
            .I(N__19126));
    LocalMux I__3524 (
            .O(N__19134),
            .I(M_this_state_qZ0Z_15));
    Odrv4 I__3523 (
            .O(N__19131),
            .I(M_this_state_qZ0Z_15));
    LocalMux I__3522 (
            .O(N__19126),
            .I(M_this_state_qZ0Z_15));
    InMux I__3521 (
            .O(N__19119),
            .I(N__19116));
    LocalMux I__3520 (
            .O(N__19116),
            .I(N__19112));
    InMux I__3519 (
            .O(N__19115),
            .I(N__19107));
    Span4Mux_h I__3518 (
            .O(N__19112),
            .I(N__19104));
    InMux I__3517 (
            .O(N__19111),
            .I(N__19099));
    InMux I__3516 (
            .O(N__19110),
            .I(N__19099));
    LocalMux I__3515 (
            .O(N__19107),
            .I(M_this_state_qZ0Z_14));
    Odrv4 I__3514 (
            .O(N__19104),
            .I(M_this_state_qZ0Z_14));
    LocalMux I__3513 (
            .O(N__19099),
            .I(M_this_state_qZ0Z_14));
    InMux I__3512 (
            .O(N__19092),
            .I(N__19088));
    InMux I__3511 (
            .O(N__19091),
            .I(N__19083));
    LocalMux I__3510 (
            .O(N__19088),
            .I(N__19080));
    InMux I__3509 (
            .O(N__19087),
            .I(N__19075));
    InMux I__3508 (
            .O(N__19086),
            .I(N__19075));
    LocalMux I__3507 (
            .O(N__19083),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__3506 (
            .O(N__19080),
            .I(M_this_state_qZ0Z_13));
    LocalMux I__3505 (
            .O(N__19075),
            .I(M_this_state_qZ0Z_13));
    InMux I__3504 (
            .O(N__19068),
            .I(N__19065));
    LocalMux I__3503 (
            .O(N__19065),
            .I(N__19062));
    Odrv4 I__3502 (
            .O(N__19062),
            .I(\this_start_data_delay.N_112_0 ));
    InMux I__3501 (
            .O(N__19059),
            .I(N__19053));
    InMux I__3500 (
            .O(N__19058),
            .I(N__19053));
    LocalMux I__3499 (
            .O(N__19053),
            .I(\this_start_data_delay.N_80_0 ));
    CascadeMux I__3498 (
            .O(N__19050),
            .I(\this_start_data_delay.un1_M_this_state_q_1_i_a2_0_aZ0Z2_cascade_ ));
    InMux I__3497 (
            .O(N__19047),
            .I(N__19043));
    InMux I__3496 (
            .O(N__19046),
            .I(N__19040));
    LocalMux I__3495 (
            .O(N__19043),
            .I(N__19037));
    LocalMux I__3494 (
            .O(N__19040),
            .I(N__19034));
    Span4Mux_h I__3493 (
            .O(N__19037),
            .I(N__19031));
    Span4Mux_h I__3492 (
            .O(N__19034),
            .I(N__19028));
    Odrv4 I__3491 (
            .O(N__19031),
            .I(\this_start_data_delay.N_76_1 ));
    Odrv4 I__3490 (
            .O(N__19028),
            .I(\this_start_data_delay.N_76_1 ));
    InMux I__3489 (
            .O(N__19023),
            .I(N__19020));
    LocalMux I__3488 (
            .O(N__19020),
            .I(\this_vga_signals.mult1_un54_sum_ac0_4_x1 ));
    CascadeMux I__3487 (
            .O(N__19017),
            .I(\this_vga_signals.mult1_un47_sum_c3_cascade_ ));
    InMux I__3486 (
            .O(N__19014),
            .I(N__19011));
    LocalMux I__3485 (
            .O(N__19011),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1 ));
    InMux I__3484 (
            .O(N__19008),
            .I(N__19005));
    LocalMux I__3483 (
            .O(N__19005),
            .I(N__19001));
    InMux I__3482 (
            .O(N__19004),
            .I(N__18997));
    Span4Mux_h I__3481 (
            .O(N__19001),
            .I(N__18994));
    InMux I__3480 (
            .O(N__19000),
            .I(N__18991));
    LocalMux I__3479 (
            .O(N__18997),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    Odrv4 I__3478 (
            .O(N__18994),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    LocalMux I__3477 (
            .O(N__18991),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    InMux I__3476 (
            .O(N__18984),
            .I(N__18981));
    LocalMux I__3475 (
            .O(N__18981),
            .I(\this_vga_signals.i1_mux ));
    InMux I__3474 (
            .O(N__18978),
            .I(N__18974));
    InMux I__3473 (
            .O(N__18977),
            .I(N__18971));
    LocalMux I__3472 (
            .O(N__18974),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1_0 ));
    LocalMux I__3471 (
            .O(N__18971),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1_0 ));
    CascadeMux I__3470 (
            .O(N__18966),
            .I(N__18963));
    InMux I__3469 (
            .O(N__18963),
            .I(N__18954));
    InMux I__3468 (
            .O(N__18962),
            .I(N__18954));
    InMux I__3467 (
            .O(N__18961),
            .I(N__18954));
    LocalMux I__3466 (
            .O(N__18954),
            .I(N__18948));
    InMux I__3465 (
            .O(N__18953),
            .I(N__18941));
    InMux I__3464 (
            .O(N__18952),
            .I(N__18941));
    InMux I__3463 (
            .O(N__18951),
            .I(N__18941));
    Span4Mux_h I__3462 (
            .O(N__18948),
            .I(N__18936));
    LocalMux I__3461 (
            .O(N__18941),
            .I(N__18936));
    Odrv4 I__3460 (
            .O(N__18936),
            .I(\this_vga_signals.vaddress_6 ));
    CascadeMux I__3459 (
            .O(N__18933),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_ ));
    InMux I__3458 (
            .O(N__18930),
            .I(N__18927));
    LocalMux I__3457 (
            .O(N__18927),
            .I(\this_vga_signals.mult1_un54_sum_ac0_4_x0 ));
    InMux I__3456 (
            .O(N__18924),
            .I(N__18921));
    LocalMux I__3455 (
            .O(N__18921),
            .I(N__18917));
    InMux I__3454 (
            .O(N__18920),
            .I(N__18914));
    Odrv4 I__3453 (
            .O(N__18917),
            .I(\this_vga_signals.g1_7 ));
    LocalMux I__3452 (
            .O(N__18914),
            .I(\this_vga_signals.g1_7 ));
    CascadeMux I__3451 (
            .O(N__18909),
            .I(N__18906));
    InMux I__3450 (
            .O(N__18906),
            .I(N__18903));
    LocalMux I__3449 (
            .O(N__18903),
            .I(N__18900));
    Odrv4 I__3448 (
            .O(N__18900),
            .I(\this_vga_signals.vaddress_3_6 ));
    InMux I__3447 (
            .O(N__18897),
            .I(N__18894));
    LocalMux I__3446 (
            .O(N__18894),
            .I(N__18891));
    Span4Mux_h I__3445 (
            .O(N__18891),
            .I(N__18888));
    Odrv4 I__3444 (
            .O(N__18888),
            .I(\this_vga_signals.g2_1_0 ));
    InMux I__3443 (
            .O(N__18885),
            .I(N__18879));
    InMux I__3442 (
            .O(N__18884),
            .I(N__18874));
    InMux I__3441 (
            .O(N__18883),
            .I(N__18874));
    CascadeMux I__3440 (
            .O(N__18882),
            .I(N__18871));
    LocalMux I__3439 (
            .O(N__18879),
            .I(N__18868));
    LocalMux I__3438 (
            .O(N__18874),
            .I(N__18865));
    InMux I__3437 (
            .O(N__18871),
            .I(N__18862));
    Odrv12 I__3436 (
            .O(N__18868),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0 ));
    Odrv4 I__3435 (
            .O(N__18865),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0 ));
    LocalMux I__3434 (
            .O(N__18862),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0 ));
    CascadeMux I__3433 (
            .O(N__18855),
            .I(N__18851));
    InMux I__3432 (
            .O(N__18854),
            .I(N__18846));
    InMux I__3431 (
            .O(N__18851),
            .I(N__18846));
    LocalMux I__3430 (
            .O(N__18846),
            .I(N__18843));
    Odrv4 I__3429 (
            .O(N__18843),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_2_1 ));
    InMux I__3428 (
            .O(N__18840),
            .I(N__18834));
    InMux I__3427 (
            .O(N__18839),
            .I(N__18834));
    LocalMux I__3426 (
            .O(N__18834),
            .I(N__18831));
    Odrv4 I__3425 (
            .O(N__18831),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_a4 ));
    InMux I__3424 (
            .O(N__18828),
            .I(N__18825));
    LocalMux I__3423 (
            .O(N__18825),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_1 ));
    CascadeMux I__3422 (
            .O(N__18822),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_3_cascade_ ));
    InMux I__3421 (
            .O(N__18819),
            .I(N__18810));
    InMux I__3420 (
            .O(N__18818),
            .I(N__18810));
    InMux I__3419 (
            .O(N__18817),
            .I(N__18810));
    LocalMux I__3418 (
            .O(N__18810),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_602_ns ));
    CascadeMux I__3417 (
            .O(N__18807),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ));
    InMux I__3416 (
            .O(N__18804),
            .I(N__18801));
    LocalMux I__3415 (
            .O(N__18801),
            .I(\this_vga_signals.g0_1_0 ));
    InMux I__3414 (
            .O(N__18798),
            .I(N__18794));
    InMux I__3413 (
            .O(N__18797),
            .I(N__18791));
    LocalMux I__3412 (
            .O(N__18794),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    LocalMux I__3411 (
            .O(N__18791),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    InMux I__3410 (
            .O(N__18786),
            .I(N__18778));
    InMux I__3409 (
            .O(N__18785),
            .I(N__18773));
    InMux I__3408 (
            .O(N__18784),
            .I(N__18769));
    InMux I__3407 (
            .O(N__18783),
            .I(N__18755));
    InMux I__3406 (
            .O(N__18782),
            .I(N__18755));
    InMux I__3405 (
            .O(N__18781),
            .I(N__18755));
    LocalMux I__3404 (
            .O(N__18778),
            .I(N__18752));
    InMux I__3403 (
            .O(N__18777),
            .I(N__18747));
    InMux I__3402 (
            .O(N__18776),
            .I(N__18747));
    LocalMux I__3401 (
            .O(N__18773),
            .I(N__18744));
    InMux I__3400 (
            .O(N__18772),
            .I(N__18741));
    LocalMux I__3399 (
            .O(N__18769),
            .I(N__18738));
    InMux I__3398 (
            .O(N__18768),
            .I(N__18731));
    InMux I__3397 (
            .O(N__18767),
            .I(N__18731));
    InMux I__3396 (
            .O(N__18766),
            .I(N__18731));
    InMux I__3395 (
            .O(N__18765),
            .I(N__18726));
    InMux I__3394 (
            .O(N__18764),
            .I(N__18726));
    InMux I__3393 (
            .O(N__18763),
            .I(N__18721));
    InMux I__3392 (
            .O(N__18762),
            .I(N__18721));
    LocalMux I__3391 (
            .O(N__18755),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__3390 (
            .O(N__18752),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__3389 (
            .O(N__18747),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__3388 (
            .O(N__18744),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__3387 (
            .O(N__18741),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__3386 (
            .O(N__18738),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__3385 (
            .O(N__18731),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__3384 (
            .O(N__18726),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__3383 (
            .O(N__18721),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    InMux I__3382 (
            .O(N__18702),
            .I(N__18699));
    LocalMux I__3381 (
            .O(N__18699),
            .I(N__18696));
    Span4Mux_h I__3380 (
            .O(N__18696),
            .I(N__18693));
    Odrv4 I__3379 (
            .O(N__18693),
            .I(\this_vga_signals.g0_5_2_0 ));
    InMux I__3378 (
            .O(N__18690),
            .I(N__18687));
    LocalMux I__3377 (
            .O(N__18687),
            .I(N_28_0));
    InMux I__3376 (
            .O(N__18684),
            .I(N__18681));
    LocalMux I__3375 (
            .O(N__18681),
            .I(\this_start_data_delay.N_82 ));
    CascadeMux I__3374 (
            .O(N__18678),
            .I(\this_start_data_delay.N_82_cascade_ ));
    InMux I__3373 (
            .O(N__18675),
            .I(N__18670));
    InMux I__3372 (
            .O(N__18674),
            .I(N__18665));
    InMux I__3371 (
            .O(N__18673),
            .I(N__18665));
    LocalMux I__3370 (
            .O(N__18670),
            .I(M_this_substate_qZ0));
    LocalMux I__3369 (
            .O(N__18665),
            .I(M_this_substate_qZ0));
    InMux I__3368 (
            .O(N__18660),
            .I(N__18657));
    LocalMux I__3367 (
            .O(N__18657),
            .I(N__18654));
    Span4Mux_v I__3366 (
            .O(N__18654),
            .I(N__18651));
    Odrv4 I__3365 (
            .O(N__18651),
            .I(\this_vga_signals.g0_0_x4_0_0 ));
    CascadeMux I__3364 (
            .O(N__18648),
            .I(\this_vga_signals.vaddress_c2_cascade_ ));
    CascadeMux I__3363 (
            .O(N__18645),
            .I(\this_vga_signals.N_5_2_1_cascade_ ));
    CascadeMux I__3362 (
            .O(N__18642),
            .I(\this_vga_signals.g0_5_0_cascade_ ));
    CascadeMux I__3361 (
            .O(N__18639),
            .I(\this_vga_signals.g0_1_1_cascade_ ));
    InMux I__3360 (
            .O(N__18636),
            .I(N__18633));
    LocalMux I__3359 (
            .O(N__18633),
            .I(N__18630));
    Span4Mux_v I__3358 (
            .O(N__18630),
            .I(N__18627));
    Odrv4 I__3357 (
            .O(N__18627),
            .I(\this_vga_signals.N_3_2 ));
    CascadeMux I__3356 (
            .O(N__18624),
            .I(N__18614));
    InMux I__3355 (
            .O(N__18623),
            .I(N__18611));
    CEMux I__3354 (
            .O(N__18622),
            .I(N__18605));
    CEMux I__3353 (
            .O(N__18621),
            .I(N__18602));
    InMux I__3352 (
            .O(N__18620),
            .I(N__18593));
    InMux I__3351 (
            .O(N__18619),
            .I(N__18572));
    InMux I__3350 (
            .O(N__18618),
            .I(N__18567));
    InMux I__3349 (
            .O(N__18617),
            .I(N__18567));
    InMux I__3348 (
            .O(N__18614),
            .I(N__18564));
    LocalMux I__3347 (
            .O(N__18611),
            .I(N__18561));
    InMux I__3346 (
            .O(N__18610),
            .I(N__18554));
    InMux I__3345 (
            .O(N__18609),
            .I(N__18554));
    InMux I__3344 (
            .O(N__18608),
            .I(N__18554));
    LocalMux I__3343 (
            .O(N__18605),
            .I(N__18549));
    LocalMux I__3342 (
            .O(N__18602),
            .I(N__18549));
    InMux I__3341 (
            .O(N__18601),
            .I(N__18536));
    InMux I__3340 (
            .O(N__18600),
            .I(N__18536));
    InMux I__3339 (
            .O(N__18599),
            .I(N__18536));
    InMux I__3338 (
            .O(N__18598),
            .I(N__18536));
    InMux I__3337 (
            .O(N__18597),
            .I(N__18536));
    InMux I__3336 (
            .O(N__18596),
            .I(N__18536));
    LocalMux I__3335 (
            .O(N__18593),
            .I(N__18533));
    InMux I__3334 (
            .O(N__18592),
            .I(N__18528));
    InMux I__3333 (
            .O(N__18591),
            .I(N__18528));
    InMux I__3332 (
            .O(N__18590),
            .I(N__18518));
    InMux I__3331 (
            .O(N__18589),
            .I(N__18518));
    InMux I__3330 (
            .O(N__18588),
            .I(N__18518));
    InMux I__3329 (
            .O(N__18587),
            .I(N__18518));
    InMux I__3328 (
            .O(N__18586),
            .I(N__18509));
    InMux I__3327 (
            .O(N__18585),
            .I(N__18509));
    InMux I__3326 (
            .O(N__18584),
            .I(N__18509));
    InMux I__3325 (
            .O(N__18583),
            .I(N__18509));
    InMux I__3324 (
            .O(N__18582),
            .I(N__18496));
    InMux I__3323 (
            .O(N__18581),
            .I(N__18496));
    InMux I__3322 (
            .O(N__18580),
            .I(N__18496));
    InMux I__3321 (
            .O(N__18579),
            .I(N__18496));
    InMux I__3320 (
            .O(N__18578),
            .I(N__18496));
    InMux I__3319 (
            .O(N__18577),
            .I(N__18496));
    InMux I__3318 (
            .O(N__18576),
            .I(N__18491));
    InMux I__3317 (
            .O(N__18575),
            .I(N__18491));
    LocalMux I__3316 (
            .O(N__18572),
            .I(N__18484));
    LocalMux I__3315 (
            .O(N__18567),
            .I(N__18484));
    LocalMux I__3314 (
            .O(N__18564),
            .I(N__18484));
    Span4Mux_v I__3313 (
            .O(N__18561),
            .I(N__18477));
    LocalMux I__3312 (
            .O(N__18554),
            .I(N__18477));
    Span4Mux_v I__3311 (
            .O(N__18549),
            .I(N__18472));
    LocalMux I__3310 (
            .O(N__18536),
            .I(N__18472));
    Span4Mux_v I__3309 (
            .O(N__18533),
            .I(N__18467));
    LocalMux I__3308 (
            .O(N__18528),
            .I(N__18467));
    InMux I__3307 (
            .O(N__18527),
            .I(N__18464));
    LocalMux I__3306 (
            .O(N__18518),
            .I(N__18457));
    LocalMux I__3305 (
            .O(N__18509),
            .I(N__18457));
    LocalMux I__3304 (
            .O(N__18496),
            .I(N__18457));
    LocalMux I__3303 (
            .O(N__18491),
            .I(N__18452));
    Span4Mux_v I__3302 (
            .O(N__18484),
            .I(N__18452));
    InMux I__3301 (
            .O(N__18483),
            .I(N__18449));
    InMux I__3300 (
            .O(N__18482),
            .I(N__18446));
    Span4Mux_v I__3299 (
            .O(N__18477),
            .I(N__18443));
    Span4Mux_h I__3298 (
            .O(N__18472),
            .I(N__18440));
    Span4Mux_h I__3297 (
            .O(N__18467),
            .I(N__18437));
    LocalMux I__3296 (
            .O(N__18464),
            .I(N__18434));
    Span4Mux_v I__3295 (
            .O(N__18457),
            .I(N__18429));
    Span4Mux_h I__3294 (
            .O(N__18452),
            .I(N__18429));
    LocalMux I__3293 (
            .O(N__18449),
            .I(N__18424));
    LocalMux I__3292 (
            .O(N__18446),
            .I(N__18424));
    Span4Mux_h I__3291 (
            .O(N__18443),
            .I(N__18421));
    Span4Mux_h I__3290 (
            .O(N__18440),
            .I(N__18418));
    Span4Mux_h I__3289 (
            .O(N__18437),
            .I(N__18415));
    Span4Mux_v I__3288 (
            .O(N__18434),
            .I(N__18408));
    Span4Mux_h I__3287 (
            .O(N__18429),
            .I(N__18408));
    Span4Mux_v I__3286 (
            .O(N__18424),
            .I(N__18408));
    Odrv4 I__3285 (
            .O(N__18421),
            .I(led23));
    Odrv4 I__3284 (
            .O(N__18418),
            .I(led23));
    Odrv4 I__3283 (
            .O(N__18415),
            .I(led23));
    Odrv4 I__3282 (
            .O(N__18408),
            .I(led23));
    CascadeMux I__3281 (
            .O(N__18399),
            .I(N__18396));
    InMux I__3280 (
            .O(N__18396),
            .I(N__18393));
    LocalMux I__3279 (
            .O(N__18393),
            .I(N__18390));
    Odrv4 I__3278 (
            .O(N__18390),
            .I(\this_start_data_delay.dmalto4_0_a2Z0Z_1 ));
    InMux I__3277 (
            .O(N__18387),
            .I(N__18384));
    LocalMux I__3276 (
            .O(N__18384),
            .I(\this_start_data_delay.N_115 ));
    CascadeMux I__3275 (
            .O(N__18381),
            .I(N__18378));
    InMux I__3274 (
            .O(N__18378),
            .I(N__18375));
    LocalMux I__3273 (
            .O(N__18375),
            .I(\this_start_data_delay.N_69 ));
    InMux I__3272 (
            .O(N__18372),
            .I(N__18369));
    LocalMux I__3271 (
            .O(N__18369),
            .I(N__18366));
    Span4Mux_v I__3270 (
            .O(N__18366),
            .I(N__18363));
    Sp12to4 I__3269 (
            .O(N__18363),
            .I(N__18360));
    Span12Mux_h I__3268 (
            .O(N__18360),
            .I(N__18357));
    Odrv12 I__3267 (
            .O(N__18357),
            .I(port_address_in_5));
    CascadeMux I__3266 (
            .O(N__18354),
            .I(N__18351));
    InMux I__3265 (
            .O(N__18351),
            .I(N__18348));
    LocalMux I__3264 (
            .O(N__18348),
            .I(N__18345));
    Sp12to4 I__3263 (
            .O(N__18345),
            .I(N__18342));
    Span12Mux_v I__3262 (
            .O(N__18342),
            .I(N__18339));
    Span12Mux_h I__3261 (
            .O(N__18339),
            .I(N__18336));
    Odrv12 I__3260 (
            .O(N__18336),
            .I(port_address_in_6));
    CascadeMux I__3259 (
            .O(N__18333),
            .I(\this_start_data_delay.N_47_0_cascade_ ));
    CascadeMux I__3258 (
            .O(N__18330),
            .I(\this_start_data_delay.N_48_0_cascade_ ));
    CascadeMux I__3257 (
            .O(N__18327),
            .I(\this_vga_signals.mult1_un54_sum_axb1_cascade_ ));
    InMux I__3256 (
            .O(N__18324),
            .I(N__18320));
    InMux I__3255 (
            .O(N__18323),
            .I(N__18317));
    LocalMux I__3254 (
            .O(N__18320),
            .I(N__18313));
    LocalMux I__3253 (
            .O(N__18317),
            .I(N__18310));
    InMux I__3252 (
            .O(N__18316),
            .I(N__18307));
    Span4Mux_v I__3251 (
            .O(N__18313),
            .I(N__18304));
    Odrv4 I__3250 (
            .O(N__18310),
            .I(\this_vga_signals.if_N_9_i ));
    LocalMux I__3249 (
            .O(N__18307),
            .I(\this_vga_signals.if_N_9_i ));
    Odrv4 I__3248 (
            .O(N__18304),
            .I(\this_vga_signals.if_N_9_i ));
    InMux I__3247 (
            .O(N__18297),
            .I(N__18294));
    LocalMux I__3246 (
            .O(N__18294),
            .I(N__18289));
    InMux I__3245 (
            .O(N__18293),
            .I(N__18286));
    InMux I__3244 (
            .O(N__18292),
            .I(N__18283));
    Odrv4 I__3243 (
            .O(N__18289),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__3242 (
            .O(N__18286),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__3241 (
            .O(N__18283),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    InMux I__3240 (
            .O(N__18276),
            .I(N__18273));
    LocalMux I__3239 (
            .O(N__18273),
            .I(\this_vga_signals.SUM_2_0_1 ));
    InMux I__3238 (
            .O(N__18270),
            .I(N__18267));
    LocalMux I__3237 (
            .O(N__18267),
            .I(\this_vga_signals.mult1_un47_sum_c3_1_0 ));
    CascadeMux I__3236 (
            .O(N__18264),
            .I(\this_vga_signals.mult1_un47_sum_c3_1_0_cascade_ ));
    InMux I__3235 (
            .O(N__18261),
            .I(N__18252));
    InMux I__3234 (
            .O(N__18260),
            .I(N__18252));
    InMux I__3233 (
            .O(N__18259),
            .I(N__18244));
    InMux I__3232 (
            .O(N__18258),
            .I(N__18237));
    InMux I__3231 (
            .O(N__18257),
            .I(N__18237));
    LocalMux I__3230 (
            .O(N__18252),
            .I(N__18226));
    InMux I__3229 (
            .O(N__18251),
            .I(N__18215));
    InMux I__3228 (
            .O(N__18250),
            .I(N__18215));
    InMux I__3227 (
            .O(N__18249),
            .I(N__18215));
    InMux I__3226 (
            .O(N__18248),
            .I(N__18215));
    InMux I__3225 (
            .O(N__18247),
            .I(N__18215));
    LocalMux I__3224 (
            .O(N__18244),
            .I(N__18212));
    InMux I__3223 (
            .O(N__18243),
            .I(N__18207));
    InMux I__3222 (
            .O(N__18242),
            .I(N__18207));
    LocalMux I__3221 (
            .O(N__18237),
            .I(N__18204));
    InMux I__3220 (
            .O(N__18236),
            .I(N__18201));
    InMux I__3219 (
            .O(N__18235),
            .I(N__18194));
    InMux I__3218 (
            .O(N__18234),
            .I(N__18194));
    InMux I__3217 (
            .O(N__18233),
            .I(N__18194));
    InMux I__3216 (
            .O(N__18232),
            .I(N__18185));
    InMux I__3215 (
            .O(N__18231),
            .I(N__18185));
    InMux I__3214 (
            .O(N__18230),
            .I(N__18185));
    InMux I__3213 (
            .O(N__18229),
            .I(N__18185));
    Odrv4 I__3212 (
            .O(N__18226),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__3211 (
            .O(N__18215),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    Odrv4 I__3210 (
            .O(N__18212),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__3209 (
            .O(N__18207),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    Odrv4 I__3208 (
            .O(N__18204),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__3207 (
            .O(N__18201),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__3206 (
            .O(N__18194),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__3205 (
            .O(N__18185),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    InMux I__3204 (
            .O(N__18168),
            .I(N__18165));
    LocalMux I__3203 (
            .O(N__18165),
            .I(\this_vga_signals.g2_4 ));
    InMux I__3202 (
            .O(N__18162),
            .I(N__18159));
    LocalMux I__3201 (
            .O(N__18159),
            .I(N__18156));
    Odrv4 I__3200 (
            .O(N__18156),
            .I(\this_vga_signals.m12_0_1 ));
    CascadeMux I__3199 (
            .O(N__18153),
            .I(N__18150));
    InMux I__3198 (
            .O(N__18150),
            .I(N__18147));
    LocalMux I__3197 (
            .O(N__18147),
            .I(N__18144));
    Odrv4 I__3196 (
            .O(N__18144),
            .I(\this_start_data_delay.N_400 ));
    CascadeMux I__3195 (
            .O(N__18141),
            .I(\this_vga_signals.N_4_3_0_cascade_ ));
    InMux I__3194 (
            .O(N__18138),
            .I(N__18135));
    LocalMux I__3193 (
            .O(N__18135),
            .I(\this_vga_signals.N_14_0 ));
    InMux I__3192 (
            .O(N__18132),
            .I(N__18129));
    LocalMux I__3191 (
            .O(N__18129),
            .I(\this_vga_signals.g1 ));
    InMux I__3190 (
            .O(N__18126),
            .I(N__18123));
    LocalMux I__3189 (
            .O(N__18123),
            .I(\this_vga_signals.g0_10_1 ));
    InMux I__3188 (
            .O(N__18120),
            .I(N__18117));
    LocalMux I__3187 (
            .O(N__18117),
            .I(\this_vga_signals.N_24_mux ));
    InMux I__3186 (
            .O(N__18114),
            .I(N__18111));
    LocalMux I__3185 (
            .O(N__18111),
            .I(\this_vga_signals.g1_2 ));
    CascadeMux I__3184 (
            .O(N__18108),
            .I(N__18105));
    InMux I__3183 (
            .O(N__18105),
            .I(N__18102));
    LocalMux I__3182 (
            .O(N__18102),
            .I(\this_vga_signals.g0_3_0_a3_3 ));
    InMux I__3181 (
            .O(N__18099),
            .I(N__18095));
    InMux I__3180 (
            .O(N__18098),
            .I(N__18092));
    LocalMux I__3179 (
            .O(N__18095),
            .I(N__18089));
    LocalMux I__3178 (
            .O(N__18092),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    Odrv4 I__3177 (
            .O(N__18089),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    CascadeMux I__3176 (
            .O(N__18084),
            .I(\this_vga_signals.mult1_un61_sum_axb2_0_cascade_ ));
    InMux I__3175 (
            .O(N__18081),
            .I(N__18075));
    InMux I__3174 (
            .O(N__18080),
            .I(N__18068));
    InMux I__3173 (
            .O(N__18079),
            .I(N__18068));
    InMux I__3172 (
            .O(N__18078),
            .I(N__18068));
    LocalMux I__3171 (
            .O(N__18075),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d));
    LocalMux I__3170 (
            .O(N__18068),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d));
    InMux I__3169 (
            .O(N__18063),
            .I(N__18060));
    LocalMux I__3168 (
            .O(N__18060),
            .I(\this_vga_signals.g2_0 ));
    CascadeMux I__3167 (
            .O(N__18057),
            .I(N__18054));
    InMux I__3166 (
            .O(N__18054),
            .I(N__18051));
    LocalMux I__3165 (
            .O(N__18051),
            .I(N__18048));
    Span4Mux_h I__3164 (
            .O(N__18048),
            .I(N__18044));
    InMux I__3163 (
            .O(N__18047),
            .I(N__18041));
    Odrv4 I__3162 (
            .O(N__18044),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2 ));
    LocalMux I__3161 (
            .O(N__18041),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2 ));
    CascadeMux I__3160 (
            .O(N__18036),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_cascade_));
    InMux I__3159 (
            .O(N__18033),
            .I(N__18030));
    LocalMux I__3158 (
            .O(N__18030),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_0 ));
    InMux I__3157 (
            .O(N__18027),
            .I(N__18023));
    InMux I__3156 (
            .O(N__18026),
            .I(N__18020));
    LocalMux I__3155 (
            .O(N__18023),
            .I(N__18017));
    LocalMux I__3154 (
            .O(N__18020),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_0 ));
    Odrv4 I__3153 (
            .O(N__18017),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_0 ));
    CascadeMux I__3152 (
            .O(N__18012),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_0_cascade_ ));
    CascadeMux I__3151 (
            .O(N__18009),
            .I(N__18004));
    InMux I__3150 (
            .O(N__18008),
            .I(N__18000));
    InMux I__3149 (
            .O(N__18007),
            .I(N__17995));
    InMux I__3148 (
            .O(N__18004),
            .I(N__17995));
    InMux I__3147 (
            .O(N__18003),
            .I(N__17992));
    LocalMux I__3146 (
            .O(N__18000),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__3145 (
            .O(N__17995),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__3144 (
            .O(N__17992),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    InMux I__3143 (
            .O(N__17985),
            .I(N__17982));
    LocalMux I__3142 (
            .O(N__17982),
            .I(\this_vga_signals.mult1_un75_sum_axb1_i_0 ));
    CascadeMux I__3141 (
            .O(N__17979),
            .I(\this_vga_signals.N_4_2_cascade_ ));
    InMux I__3140 (
            .O(N__17976),
            .I(N__17970));
    InMux I__3139 (
            .O(N__17975),
            .I(N__17970));
    LocalMux I__3138 (
            .O(N__17970),
            .I(\this_vga_signals.if_m1_0_0 ));
    InMux I__3137 (
            .O(N__17967),
            .I(N__17964));
    LocalMux I__3136 (
            .O(N__17964),
            .I(N__17961));
    Odrv12 I__3135 (
            .O(N__17961),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d_0_0 ));
    CascadeMux I__3134 (
            .O(N__17958),
            .I(N__17954));
    InMux I__3133 (
            .O(N__17957),
            .I(N__17950));
    InMux I__3132 (
            .O(N__17954),
            .I(N__17947));
    InMux I__3131 (
            .O(N__17953),
            .I(N__17944));
    LocalMux I__3130 (
            .O(N__17950),
            .I(N__17939));
    LocalMux I__3129 (
            .O(N__17947),
            .I(N__17939));
    LocalMux I__3128 (
            .O(N__17944),
            .I(\this_vga_signals.mult1_un61_sum_axb2_0 ));
    Odrv4 I__3127 (
            .O(N__17939),
            .I(\this_vga_signals.mult1_un61_sum_axb2_0 ));
    CascadeMux I__3126 (
            .O(N__17934),
            .I(N__17930));
    InMux I__3125 (
            .O(N__17933),
            .I(N__17925));
    InMux I__3124 (
            .O(N__17930),
            .I(N__17920));
    InMux I__3123 (
            .O(N__17929),
            .I(N__17920));
    InMux I__3122 (
            .O(N__17928),
            .I(N__17917));
    LocalMux I__3121 (
            .O(N__17925),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1));
    LocalMux I__3120 (
            .O(N__17920),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1));
    LocalMux I__3119 (
            .O(N__17917),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1));
    CascadeMux I__3118 (
            .O(N__17910),
            .I(N__17907));
    InMux I__3117 (
            .O(N__17907),
            .I(N__17903));
    InMux I__3116 (
            .O(N__17906),
            .I(N__17900));
    LocalMux I__3115 (
            .O(N__17903),
            .I(\this_vga_signals.mult1_un75_sum_axb1_1 ));
    LocalMux I__3114 (
            .O(N__17900),
            .I(\this_vga_signals.mult1_un75_sum_axb1_1 ));
    CascadeMux I__3113 (
            .O(N__17895),
            .I(\this_vga_signals.mult1_un54_sum_ac0_4_cascade_ ));
    CascadeMux I__3112 (
            .O(N__17892),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ));
    CascadeMux I__3111 (
            .O(N__17889),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_0_2_cascade_ ));
    InMux I__3110 (
            .O(N__17886),
            .I(N__17877));
    InMux I__3109 (
            .O(N__17885),
            .I(N__17877));
    InMux I__3108 (
            .O(N__17884),
            .I(N__17877));
    LocalMux I__3107 (
            .O(N__17877),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3));
    CascadeMux I__3106 (
            .O(N__17874),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_cascade_));
    InMux I__3105 (
            .O(N__17871),
            .I(N__17868));
    LocalMux I__3104 (
            .O(N__17868),
            .I(\this_vga_signals.mult1_un61_sum_c3_0 ));
    InMux I__3103 (
            .O(N__17865),
            .I(N__17862));
    LocalMux I__3102 (
            .O(N__17862),
            .I(N__17859));
    Span4Mux_h I__3101 (
            .O(N__17859),
            .I(N__17856));
    Span4Mux_h I__3100 (
            .O(N__17856),
            .I(N__17853));
    Span4Mux_h I__3099 (
            .O(N__17853),
            .I(N__17850));
    Odrv4 I__3098 (
            .O(N__17850),
            .I(\this_vga_signals.if_m2 ));
    InMux I__3097 (
            .O(N__17847),
            .I(N__17844));
    LocalMux I__3096 (
            .O(N__17844),
            .I(\this_vga_signals.if_m1_9_0 ));
    CascadeMux I__3095 (
            .O(N__17841),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_cascade_ ));
    InMux I__3094 (
            .O(N__17838),
            .I(N__17834));
    InMux I__3093 (
            .O(N__17837),
            .I(N__17831));
    LocalMux I__3092 (
            .O(N__17834),
            .I(\this_vga_signals.if_m2_3_1 ));
    LocalMux I__3091 (
            .O(N__17831),
            .I(\this_vga_signals.if_m2_3_1 ));
    InMux I__3090 (
            .O(N__17826),
            .I(N__17823));
    LocalMux I__3089 (
            .O(N__17823),
            .I(\this_vga_signals.if_i4_mux ));
    InMux I__3088 (
            .O(N__17820),
            .I(N__17817));
    LocalMux I__3087 (
            .O(N__17817),
            .I(\this_vga_signals.g0_1 ));
    CascadeMux I__3086 (
            .O(N__17814),
            .I(N__17811));
    InMux I__3085 (
            .O(N__17811),
            .I(N__17808));
    LocalMux I__3084 (
            .O(N__17808),
            .I(N__17805));
    Span4Mux_h I__3083 (
            .O(N__17805),
            .I(N__17802));
    Odrv4 I__3082 (
            .O(N__17802),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0 ));
    InMux I__3081 (
            .O(N__17799),
            .I(N__17796));
    LocalMux I__3080 (
            .O(N__17796),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_0_2_1 ));
    CascadeMux I__3079 (
            .O(N__17793),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_0_2_1_cascade_ ));
    CascadeMux I__3078 (
            .O(N__17790),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_cascade_ ));
    CascadeMux I__3077 (
            .O(N__17787),
            .I(N__17784));
    InMux I__3076 (
            .O(N__17784),
            .I(N__17781));
    LocalMux I__3075 (
            .O(N__17781),
            .I(M_this_state_d_0_sqmuxa_2));
    CascadeMux I__3074 (
            .O(N__17778),
            .I(\this_start_data_delay.N_65_cascade_ ));
    InMux I__3073 (
            .O(N__17775),
            .I(N__17772));
    LocalMux I__3072 (
            .O(N__17772),
            .I(N__17769));
    Odrv4 I__3071 (
            .O(N__17769),
            .I(\this_start_data_delay.N_42_0 ));
    InMux I__3070 (
            .O(N__17766),
            .I(N__17763));
    LocalMux I__3069 (
            .O(N__17763),
            .I(N__17759));
    InMux I__3068 (
            .O(N__17762),
            .I(N__17756));
    Span4Mux_v I__3067 (
            .O(N__17759),
            .I(N__17753));
    LocalMux I__3066 (
            .O(N__17756),
            .I(N__17750));
    Odrv4 I__3065 (
            .O(N__17753),
            .I(\this_start_data_delay.N_43_0 ));
    Odrv4 I__3064 (
            .O(N__17750),
            .I(\this_start_data_delay.N_43_0 ));
    IoInMux I__3063 (
            .O(N__17745),
            .I(N__17742));
    LocalMux I__3062 (
            .O(N__17742),
            .I(N__17739));
    Span4Mux_s1_h I__3061 (
            .O(N__17739),
            .I(N__17736));
    Span4Mux_h I__3060 (
            .O(N__17736),
            .I(N__17731));
    InMux I__3059 (
            .O(N__17735),
            .I(N__17728));
    InMux I__3058 (
            .O(N__17734),
            .I(N__17725));
    Sp12to4 I__3057 (
            .O(N__17731),
            .I(N__17721));
    LocalMux I__3056 (
            .O(N__17728),
            .I(N__17718));
    LocalMux I__3055 (
            .O(N__17725),
            .I(N__17715));
    CascadeMux I__3054 (
            .O(N__17724),
            .I(N__17712));
    Span12Mux_v I__3053 (
            .O(N__17721),
            .I(N__17707));
    Span12Mux_s5_h I__3052 (
            .O(N__17718),
            .I(N__17707));
    Span4Mux_h I__3051 (
            .O(N__17715),
            .I(N__17704));
    InMux I__3050 (
            .O(N__17712),
            .I(N__17701));
    Span12Mux_h I__3049 (
            .O(N__17707),
            .I(N__17698));
    Span4Mux_v I__3048 (
            .O(N__17704),
            .I(N__17693));
    LocalMux I__3047 (
            .O(N__17701),
            .I(N__17693));
    Odrv12 I__3046 (
            .O(N__17698),
            .I(dma_0));
    Odrv4 I__3045 (
            .O(N__17693),
            .I(dma_0));
    CascadeMux I__3044 (
            .O(N__17688),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2_cascade_ ));
    CascadeMux I__3043 (
            .O(N__17685),
            .I(\this_vga_signals.g0_i_x4_1_cascade_ ));
    CascadeMux I__3042 (
            .O(N__17682),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_1_0_0_cascade_ ));
    InMux I__3041 (
            .O(N__17679),
            .I(N__17676));
    LocalMux I__3040 (
            .O(N__17676),
            .I(\this_vga_signals.g0_9_N_3L3 ));
    InMux I__3039 (
            .O(N__17673),
            .I(N__17670));
    LocalMux I__3038 (
            .O(N__17670),
            .I(N__17667));
    Odrv4 I__3037 (
            .O(N__17667),
            .I(\this_vga_signals.g0_i_a4_4_0_0 ));
    CEMux I__3036 (
            .O(N__17664),
            .I(N__17660));
    CEMux I__3035 (
            .O(N__17663),
            .I(N__17656));
    LocalMux I__3034 (
            .O(N__17660),
            .I(N__17653));
    CEMux I__3033 (
            .O(N__17659),
            .I(N__17650));
    LocalMux I__3032 (
            .O(N__17656),
            .I(N__17646));
    Span4Mux_v I__3031 (
            .O(N__17653),
            .I(N__17642));
    LocalMux I__3030 (
            .O(N__17650),
            .I(N__17639));
    CEMux I__3029 (
            .O(N__17649),
            .I(N__17636));
    Span4Mux_v I__3028 (
            .O(N__17646),
            .I(N__17633));
    CEMux I__3027 (
            .O(N__17645),
            .I(N__17630));
    Span4Mux_h I__3026 (
            .O(N__17642),
            .I(N__17625));
    Span4Mux_v I__3025 (
            .O(N__17639),
            .I(N__17625));
    LocalMux I__3024 (
            .O(N__17636),
            .I(N__17622));
    Span4Mux_h I__3023 (
            .O(N__17633),
            .I(N__17617));
    LocalMux I__3022 (
            .O(N__17630),
            .I(N__17617));
    Span4Mux_h I__3021 (
            .O(N__17625),
            .I(N__17612));
    Span4Mux_h I__3020 (
            .O(N__17622),
            .I(N__17612));
    Sp12to4 I__3019 (
            .O(N__17617),
            .I(N__17609));
    Span4Mux_h I__3018 (
            .O(N__17612),
            .I(N__17606));
    Odrv12 I__3017 (
            .O(N__17609),
            .I(N_1422_0));
    Odrv4 I__3016 (
            .O(N__17606),
            .I(N_1422_0));
    CascadeMux I__3015 (
            .O(N__17601),
            .I(M_this_state_d_0_sqmuxa_2_cascade_));
    InMux I__3014 (
            .O(N__17598),
            .I(N__17594));
    InMux I__3013 (
            .O(N__17597),
            .I(N__17591));
    LocalMux I__3012 (
            .O(N__17594),
            .I(\this_vga_signals.if_m1_0 ));
    LocalMux I__3011 (
            .O(N__17591),
            .I(\this_vga_signals.if_m1_0 ));
    InMux I__3010 (
            .O(N__17586),
            .I(N__17583));
    LocalMux I__3009 (
            .O(N__17583),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0 ));
    CascadeMux I__3008 (
            .O(N__17580),
            .I(N__17577));
    InMux I__3007 (
            .O(N__17577),
            .I(N__17574));
    LocalMux I__3006 (
            .O(N__17574),
            .I(\this_vga_signals.g0_3_0_a3 ));
    InMux I__3005 (
            .O(N__17571),
            .I(N__17568));
    LocalMux I__3004 (
            .O(N__17568),
            .I(\this_vga_signals.g1_0 ));
    CascadeMux I__3003 (
            .O(N__17565),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_1_0_cascade_ ));
    InMux I__3002 (
            .O(N__17562),
            .I(N__17559));
    LocalMux I__3001 (
            .O(N__17559),
            .I(\this_vga_signals.g0_i_x4_7_0_0 ));
    CascadeMux I__3000 (
            .O(N__17556),
            .I(\this_vga_signals.g0_9_N_2L1_cascade_ ));
    CascadeMux I__2999 (
            .O(N__17553),
            .I(\this_vga_signals.mult1_un68_sum_c3_cascade_ ));
    CascadeMux I__2998 (
            .O(N__17550),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_ ));
    InMux I__2997 (
            .O(N__17547),
            .I(N__17543));
    InMux I__2996 (
            .O(N__17546),
            .I(N__17540));
    LocalMux I__2995 (
            .O(N__17543),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    LocalMux I__2994 (
            .O(N__17540),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    CascadeMux I__2993 (
            .O(N__17535),
            .I(\this_vga_signals.if_m2_3_1_cascade_ ));
    CascadeMux I__2992 (
            .O(N__17532),
            .I(\this_vga_signals.g2_cascade_ ));
    InMux I__2991 (
            .O(N__17529),
            .I(N__17526));
    LocalMux I__2990 (
            .O(N__17526),
            .I(\this_vga_signals.g0_4 ));
    InMux I__2989 (
            .O(N__17523),
            .I(N__17520));
    LocalMux I__2988 (
            .O(N__17520),
            .I(\this_vga_signals.g1_0_0 ));
    CascadeMux I__2987 (
            .O(N__17517),
            .I(\this_vga_signals.if_m1_0_cascade_ ));
    InMux I__2986 (
            .O(N__17514),
            .I(N__17511));
    LocalMux I__2985 (
            .O(N__17511),
            .I(N__17508));
    Odrv4 I__2984 (
            .O(N__17508),
            .I(\this_vga_signals.N_129_i ));
    InMux I__2983 (
            .O(N__17505),
            .I(N__17502));
    LocalMux I__2982 (
            .O(N__17502),
            .I(N__17499));
    Sp12to4 I__2981 (
            .O(N__17499),
            .I(N__17496));
    Span12Mux_v I__2980 (
            .O(N__17496),
            .I(N__17493));
    Odrv12 I__2979 (
            .O(N__17493),
            .I(\this_sprites_ram.mem_out_bus7_2 ));
    InMux I__2978 (
            .O(N__17490),
            .I(N__17487));
    LocalMux I__2977 (
            .O(N__17487),
            .I(N__17484));
    Span4Mux_h I__2976 (
            .O(N__17484),
            .I(N__17481));
    Span4Mux_h I__2975 (
            .O(N__17481),
            .I(N__17478));
    Odrv4 I__2974 (
            .O(N__17478),
            .I(\this_sprites_ram.mem_out_bus3_2 ));
    InMux I__2973 (
            .O(N__17475),
            .I(N__17472));
    LocalMux I__2972 (
            .O(N__17472),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ));
    InMux I__2971 (
            .O(N__17469),
            .I(N__17463));
    CascadeMux I__2970 (
            .O(N__17468),
            .I(N__17460));
    InMux I__2969 (
            .O(N__17467),
            .I(N__17456));
    InMux I__2968 (
            .O(N__17466),
            .I(N__17453));
    LocalMux I__2967 (
            .O(N__17463),
            .I(N__17450));
    InMux I__2966 (
            .O(N__17460),
            .I(N__17447));
    InMux I__2965 (
            .O(N__17459),
            .I(N__17444));
    LocalMux I__2964 (
            .O(N__17456),
            .I(N__17439));
    LocalMux I__2963 (
            .O(N__17453),
            .I(N__17439));
    Span4Mux_h I__2962 (
            .O(N__17450),
            .I(N__17430));
    LocalMux I__2961 (
            .O(N__17447),
            .I(N__17430));
    LocalMux I__2960 (
            .O(N__17444),
            .I(N__17430));
    Span4Mux_v I__2959 (
            .O(N__17439),
            .I(N__17430));
    Odrv4 I__2958 (
            .O(N__17430),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    InMux I__2957 (
            .O(N__17427),
            .I(N__17424));
    LocalMux I__2956 (
            .O(N__17424),
            .I(N__17421));
    Span4Mux_h I__2955 (
            .O(N__17421),
            .I(N__17417));
    InMux I__2954 (
            .O(N__17420),
            .I(N__17414));
    Odrv4 I__2953 (
            .O(N__17417),
            .I(\this_ppu.M_state_q_srsts_i_a3_5_2 ));
    LocalMux I__2952 (
            .O(N__17414),
            .I(\this_ppu.M_state_q_srsts_i_a3_5_2 ));
    InMux I__2951 (
            .O(N__17409),
            .I(N__17406));
    LocalMux I__2950 (
            .O(N__17406),
            .I(N__17403));
    Span4Mux_h I__2949 (
            .O(N__17403),
            .I(N__17399));
    InMux I__2948 (
            .O(N__17402),
            .I(N__17396));
    Odrv4 I__2947 (
            .O(N__17399),
            .I(\this_ppu.M_state_q_srsts_i_a3_4_2 ));
    LocalMux I__2946 (
            .O(N__17396),
            .I(\this_ppu.M_state_q_srsts_i_a3_4_2 ));
    CascadeMux I__2945 (
            .O(N__17391),
            .I(N_2_cascade_));
    CascadeMux I__2944 (
            .O(N__17388),
            .I(\this_vga_signals.N_6_1_cascade_ ));
    InMux I__2943 (
            .O(N__17385),
            .I(N__17382));
    LocalMux I__2942 (
            .O(N__17382),
            .I(\this_vga_signals.vaddress_N_4_0 ));
    InMux I__2941 (
            .O(N__17379),
            .I(N__17376));
    LocalMux I__2940 (
            .O(N__17376),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    InMux I__2939 (
            .O(N__17373),
            .I(N__17370));
    LocalMux I__2938 (
            .O(N__17370),
            .I(\this_vga_signals.mult1_un75_sum_axb1_i_1 ));
    InMux I__2937 (
            .O(N__17367),
            .I(N__17364));
    LocalMux I__2936 (
            .O(N__17364),
            .I(\this_vga_signals.N_7_0 ));
    CEMux I__2935 (
            .O(N__17361),
            .I(N__17358));
    LocalMux I__2934 (
            .O(N__17358),
            .I(N__17354));
    CEMux I__2933 (
            .O(N__17357),
            .I(N__17349));
    Span4Mux_v I__2932 (
            .O(N__17354),
            .I(N__17346));
    CEMux I__2931 (
            .O(N__17353),
            .I(N__17343));
    CEMux I__2930 (
            .O(N__17352),
            .I(N__17340));
    LocalMux I__2929 (
            .O(N__17349),
            .I(N__17336));
    Span4Mux_h I__2928 (
            .O(N__17346),
            .I(N__17331));
    LocalMux I__2927 (
            .O(N__17343),
            .I(N__17331));
    LocalMux I__2926 (
            .O(N__17340),
            .I(N__17328));
    CEMux I__2925 (
            .O(N__17339),
            .I(N__17325));
    Span4Mux_h I__2924 (
            .O(N__17336),
            .I(N__17322));
    Span4Mux_h I__2923 (
            .O(N__17331),
            .I(N__17315));
    Span4Mux_v I__2922 (
            .O(N__17328),
            .I(N__17315));
    LocalMux I__2921 (
            .O(N__17325),
            .I(N__17315));
    Span4Mux_h I__2920 (
            .O(N__17322),
            .I(N__17312));
    Sp12to4 I__2919 (
            .O(N__17315),
            .I(N__17309));
    Odrv4 I__2918 (
            .O(N__17312),
            .I(N_1438_0));
    Odrv12 I__2917 (
            .O(N__17309),
            .I(N_1438_0));
    InMux I__2916 (
            .O(N__17304),
            .I(N__17301));
    LocalMux I__2915 (
            .O(N__17301),
            .I(\this_start_data_delay.port_data_rw_0_a2Z0Z_1 ));
    IoInMux I__2914 (
            .O(N__17298),
            .I(N__17295));
    LocalMux I__2913 (
            .O(N__17295),
            .I(N__17292));
    Span4Mux_s1_h I__2912 (
            .O(N__17292),
            .I(N__17289));
    Span4Mux_h I__2911 (
            .O(N__17289),
            .I(N__17286));
    Span4Mux_h I__2910 (
            .O(N__17286),
            .I(N__17283));
    Sp12to4 I__2909 (
            .O(N__17283),
            .I(N__17280));
    Span12Mux_v I__2908 (
            .O(N__17280),
            .I(N__17277));
    Odrv12 I__2907 (
            .O(N__17277),
            .I(port_data_rw_0_i));
    InMux I__2906 (
            .O(N__17274),
            .I(N__17271));
    LocalMux I__2905 (
            .O(N__17271),
            .I(N__17268));
    Span12Mux_v I__2904 (
            .O(N__17268),
            .I(N__17265));
    Odrv12 I__2903 (
            .O(N__17265),
            .I(\this_sprites_ram.mem_out_bus5_2 ));
    InMux I__2902 (
            .O(N__17262),
            .I(N__17259));
    LocalMux I__2901 (
            .O(N__17259),
            .I(N__17256));
    Span12Mux_v I__2900 (
            .O(N__17256),
            .I(N__17253));
    Odrv12 I__2899 (
            .O(N__17253),
            .I(\this_sprites_ram.mem_out_bus1_2 ));
    InMux I__2898 (
            .O(N__17250),
            .I(N__17247));
    LocalMux I__2897 (
            .O(N__17247),
            .I(N__17244));
    Span4Mux_h I__2896 (
            .O(N__17244),
            .I(N__17241));
    Span4Mux_h I__2895 (
            .O(N__17241),
            .I(N__17238));
    Span4Mux_h I__2894 (
            .O(N__17238),
            .I(N__17235));
    Odrv4 I__2893 (
            .O(N__17235),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    InMux I__2892 (
            .O(N__17232),
            .I(N__17229));
    LocalMux I__2891 (
            .O(N__17229),
            .I(N__17226));
    Span4Mux_h I__2890 (
            .O(N__17226),
            .I(N__17223));
    Span4Mux_h I__2889 (
            .O(N__17223),
            .I(N__17220));
    Odrv4 I__2888 (
            .O(N__17220),
            .I(\this_sprites_ram.mem_out_bus4_2 ));
    InMux I__2887 (
            .O(N__17217),
            .I(N__17214));
    LocalMux I__2886 (
            .O(N__17214),
            .I(N__17211));
    Span12Mux_v I__2885 (
            .O(N__17211),
            .I(N__17208));
    Span12Mux_v I__2884 (
            .O(N__17208),
            .I(N__17205));
    Odrv12 I__2883 (
            .O(N__17205),
            .I(\this_sprites_ram.mem_out_bus0_2 ));
    CascadeMux I__2882 (
            .O(N__17202),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ));
    InMux I__2881 (
            .O(N__17199),
            .I(N__17196));
    LocalMux I__2880 (
            .O(N__17196),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ));
    CascadeMux I__2879 (
            .O(N__17193),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ));
    InMux I__2878 (
            .O(N__17190),
            .I(N__17186));
    InMux I__2877 (
            .O(N__17189),
            .I(N__17183));
    LocalMux I__2876 (
            .O(N__17186),
            .I(N__17179));
    LocalMux I__2875 (
            .O(N__17183),
            .I(N__17176));
    InMux I__2874 (
            .O(N__17182),
            .I(N__17173));
    Span12Mux_h I__2873 (
            .O(N__17179),
            .I(N__17170));
    Span4Mux_h I__2872 (
            .O(N__17176),
            .I(N__17167));
    LocalMux I__2871 (
            .O(N__17173),
            .I(N__17164));
    Odrv12 I__2870 (
            .O(N__17170),
            .I(M_this_ppu_vram_data_2));
    Odrv4 I__2869 (
            .O(N__17167),
            .I(M_this_ppu_vram_data_2));
    Odrv12 I__2868 (
            .O(N__17164),
            .I(M_this_ppu_vram_data_2));
    InMux I__2867 (
            .O(N__17157),
            .I(N__17154));
    LocalMux I__2866 (
            .O(N__17154),
            .I(\this_ppu.un10_sprites_addr_cry_2_c_RNIQP7BZ0 ));
    InMux I__2865 (
            .O(N__17151),
            .I(N__17148));
    LocalMux I__2864 (
            .O(N__17148),
            .I(N__17145));
    Span4Mux_v I__2863 (
            .O(N__17145),
            .I(N__17142));
    Span4Mux_v I__2862 (
            .O(N__17142),
            .I(N__17139));
    Span4Mux_h I__2861 (
            .O(N__17139),
            .I(N__17136));
    Span4Mux_h I__2860 (
            .O(N__17136),
            .I(N__17133));
    Odrv4 I__2859 (
            .O(N__17133),
            .I(M_this_map_ram_read_data_5));
    InMux I__2858 (
            .O(N__17130),
            .I(N__17125));
    InMux I__2857 (
            .O(N__17129),
            .I(N__17122));
    InMux I__2856 (
            .O(N__17128),
            .I(N__17115));
    LocalMux I__2855 (
            .O(N__17125),
            .I(N__17112));
    LocalMux I__2854 (
            .O(N__17122),
            .I(N__17109));
    InMux I__2853 (
            .O(N__17121),
            .I(N__17106));
    InMux I__2852 (
            .O(N__17120),
            .I(N__17103));
    InMux I__2851 (
            .O(N__17119),
            .I(N__17098));
    InMux I__2850 (
            .O(N__17118),
            .I(N__17098));
    LocalMux I__2849 (
            .O(N__17115),
            .I(N__17095));
    Span4Mux_h I__2848 (
            .O(N__17112),
            .I(N__17092));
    Span4Mux_h I__2847 (
            .O(N__17109),
            .I(N__17089));
    LocalMux I__2846 (
            .O(N__17106),
            .I(N__17086));
    LocalMux I__2845 (
            .O(N__17103),
            .I(N__17083));
    LocalMux I__2844 (
            .O(N__17098),
            .I(N__17080));
    Span4Mux_h I__2843 (
            .O(N__17095),
            .I(N__17071));
    Span4Mux_v I__2842 (
            .O(N__17092),
            .I(N__17071));
    Span4Mux_v I__2841 (
            .O(N__17089),
            .I(N__17071));
    Span4Mux_h I__2840 (
            .O(N__17086),
            .I(N__17068));
    Span4Mux_v I__2839 (
            .O(N__17083),
            .I(N__17063));
    Span4Mux_h I__2838 (
            .O(N__17080),
            .I(N__17063));
    InMux I__2837 (
            .O(N__17079),
            .I(N__17058));
    InMux I__2836 (
            .O(N__17078),
            .I(N__17058));
    Odrv4 I__2835 (
            .O(N__17071),
            .I(M_this_vga_ramdac_en_0));
    Odrv4 I__2834 (
            .O(N__17068),
            .I(M_this_vga_ramdac_en_0));
    Odrv4 I__2833 (
            .O(N__17063),
            .I(M_this_vga_ramdac_en_0));
    LocalMux I__2832 (
            .O(N__17058),
            .I(M_this_vga_ramdac_en_0));
    CascadeMux I__2831 (
            .O(N__17049),
            .I(\this_vga_signals.mult1_un75_sum_c3_0_0_0_0_cascade_ ));
    CascadeMux I__2830 (
            .O(N__17046),
            .I(N__17043));
    InMux I__2829 (
            .O(N__17043),
            .I(N__17040));
    LocalMux I__2828 (
            .O(N__17040),
            .I(N__17037));
    Span4Mux_v I__2827 (
            .O(N__17037),
            .I(N__17034));
    Span4Mux_h I__2826 (
            .O(N__17034),
            .I(N__17031));
    Span4Mux_h I__2825 (
            .O(N__17031),
            .I(N__17028));
    Odrv4 I__2824 (
            .O(N__17028),
            .I(M_this_vga_signals_address_7));
    InMux I__2823 (
            .O(N__17025),
            .I(N__17022));
    LocalMux I__2822 (
            .O(N__17022),
            .I(\this_vga_signals.un6_vvisibilitylt9_0 ));
    InMux I__2821 (
            .O(N__17019),
            .I(N__17016));
    LocalMux I__2820 (
            .O(N__17016),
            .I(\this_vga_signals.g2_2 ));
    CascadeMux I__2819 (
            .O(N__17013),
            .I(\this_vga_signals.SUM_2_1_cascade_ ));
    CascadeMux I__2818 (
            .O(N__17010),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_1_1_cascade_ ));
    InMux I__2817 (
            .O(N__17007),
            .I(N__17004));
    LocalMux I__2816 (
            .O(N__17004),
            .I(\this_vga_signals.N_4_0_0_0 ));
    InMux I__2815 (
            .O(N__17001),
            .I(N__16998));
    LocalMux I__2814 (
            .O(N__16998),
            .I(\this_vga_signals.g3_2_0 ));
    CascadeMux I__2813 (
            .O(N__16995),
            .I(\this_vga_signals.N_6_cascade_ ));
    InMux I__2812 (
            .O(N__16992),
            .I(N__16989));
    LocalMux I__2811 (
            .O(N__16989),
            .I(\this_vga_signals.g4 ));
    InMux I__2810 (
            .O(N__16986),
            .I(N__16983));
    LocalMux I__2809 (
            .O(N__16983),
            .I(N__16979));
    InMux I__2808 (
            .O(N__16982),
            .I(N__16975));
    Span4Mux_v I__2807 (
            .O(N__16979),
            .I(N__16969));
    InMux I__2806 (
            .O(N__16978),
            .I(N__16966));
    LocalMux I__2805 (
            .O(N__16975),
            .I(N__16963));
    InMux I__2804 (
            .O(N__16974),
            .I(N__16956));
    InMux I__2803 (
            .O(N__16973),
            .I(N__16956));
    InMux I__2802 (
            .O(N__16972),
            .I(N__16956));
    Odrv4 I__2801 (
            .O(N__16969),
            .I(\this_ppu.M_last_q ));
    LocalMux I__2800 (
            .O(N__16966),
            .I(\this_ppu.M_last_q ));
    Odrv4 I__2799 (
            .O(N__16963),
            .I(\this_ppu.M_last_q ));
    LocalMux I__2798 (
            .O(N__16956),
            .I(\this_ppu.M_last_q ));
    InMux I__2797 (
            .O(N__16947),
            .I(N__16940));
    InMux I__2796 (
            .O(N__16946),
            .I(N__16937));
    InMux I__2795 (
            .O(N__16945),
            .I(N__16930));
    InMux I__2794 (
            .O(N__16944),
            .I(N__16930));
    InMux I__2793 (
            .O(N__16943),
            .I(N__16930));
    LocalMux I__2792 (
            .O(N__16940),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__2791 (
            .O(N__16937),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__2790 (
            .O(N__16930),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    InMux I__2789 (
            .O(N__16923),
            .I(N__16918));
    CascadeMux I__2788 (
            .O(N__16922),
            .I(N__16913));
    InMux I__2787 (
            .O(N__16921),
            .I(N__16910));
    LocalMux I__2786 (
            .O(N__16918),
            .I(N__16907));
    InMux I__2785 (
            .O(N__16917),
            .I(N__16904));
    InMux I__2784 (
            .O(N__16916),
            .I(N__16901));
    InMux I__2783 (
            .O(N__16913),
            .I(N__16898));
    LocalMux I__2782 (
            .O(N__16910),
            .I(M_this_vga_signals_line_clk_0));
    Odrv4 I__2781 (
            .O(N__16907),
            .I(M_this_vga_signals_line_clk_0));
    LocalMux I__2780 (
            .O(N__16904),
            .I(M_this_vga_signals_line_clk_0));
    LocalMux I__2779 (
            .O(N__16901),
            .I(M_this_vga_signals_line_clk_0));
    LocalMux I__2778 (
            .O(N__16898),
            .I(M_this_vga_signals_line_clk_0));
    CascadeMux I__2777 (
            .O(N__16887),
            .I(N__16882));
    InMux I__2776 (
            .O(N__16886),
            .I(N__16877));
    InMux I__2775 (
            .O(N__16885),
            .I(N__16877));
    InMux I__2774 (
            .O(N__16882),
            .I(N__16873));
    LocalMux I__2773 (
            .O(N__16877),
            .I(N__16868));
    InMux I__2772 (
            .O(N__16876),
            .I(N__16865));
    LocalMux I__2771 (
            .O(N__16873),
            .I(N__16862));
    InMux I__2770 (
            .O(N__16872),
            .I(N__16857));
    InMux I__2769 (
            .O(N__16871),
            .I(N__16857));
    Odrv4 I__2768 (
            .O(N__16868),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    LocalMux I__2767 (
            .O(N__16865),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    Odrv4 I__2766 (
            .O(N__16862),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    LocalMux I__2765 (
            .O(N__16857),
            .I(\this_ppu.M_state_d_0_sqmuxa ));
    CascadeMux I__2764 (
            .O(N__16848),
            .I(N__16845));
    InMux I__2763 (
            .O(N__16845),
            .I(N__16842));
    LocalMux I__2762 (
            .O(N__16842),
            .I(N__16839));
    Span4Mux_h I__2761 (
            .O(N__16839),
            .I(N__16836));
    Sp12to4 I__2760 (
            .O(N__16836),
            .I(N__16829));
    CascadeMux I__2759 (
            .O(N__16835),
            .I(N__16826));
    CascadeMux I__2758 (
            .O(N__16834),
            .I(N__16822));
    InMux I__2757 (
            .O(N__16833),
            .I(N__16817));
    CascadeMux I__2756 (
            .O(N__16832),
            .I(N__16814));
    Span12Mux_v I__2755 (
            .O(N__16829),
            .I(N__16811));
    InMux I__2754 (
            .O(N__16826),
            .I(N__16804));
    InMux I__2753 (
            .O(N__16825),
            .I(N__16804));
    InMux I__2752 (
            .O(N__16822),
            .I(N__16804));
    InMux I__2751 (
            .O(N__16821),
            .I(N__16799));
    InMux I__2750 (
            .O(N__16820),
            .I(N__16799));
    LocalMux I__2749 (
            .O(N__16817),
            .I(N__16796));
    InMux I__2748 (
            .O(N__16814),
            .I(N__16793));
    Odrv12 I__2747 (
            .O(N__16811),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__2746 (
            .O(N__16804),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__2745 (
            .O(N__16799),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__2744 (
            .O(N__16796),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__2743 (
            .O(N__16793),
            .I(M_this_ppu_vram_addr_7));
    CascadeMux I__2742 (
            .O(N__16782),
            .I(N__16779));
    CascadeBuf I__2741 (
            .O(N__16779),
            .I(N__16776));
    CascadeMux I__2740 (
            .O(N__16776),
            .I(N__16772));
    InMux I__2739 (
            .O(N__16775),
            .I(N__16768));
    InMux I__2738 (
            .O(N__16772),
            .I(N__16765));
    InMux I__2737 (
            .O(N__16771),
            .I(N__16762));
    LocalMux I__2736 (
            .O(N__16768),
            .I(N__16759));
    LocalMux I__2735 (
            .O(N__16765),
            .I(N__16756));
    LocalMux I__2734 (
            .O(N__16762),
            .I(N__16752));
    Span4Mux_v I__2733 (
            .O(N__16759),
            .I(N__16748));
    Sp12to4 I__2732 (
            .O(N__16756),
            .I(N__16745));
    InMux I__2731 (
            .O(N__16755),
            .I(N__16742));
    Span4Mux_v I__2730 (
            .O(N__16752),
            .I(N__16739));
    InMux I__2729 (
            .O(N__16751),
            .I(N__16736));
    Sp12to4 I__2728 (
            .O(N__16748),
            .I(N__16731));
    Span12Mux_v I__2727 (
            .O(N__16745),
            .I(N__16731));
    LocalMux I__2726 (
            .O(N__16742),
            .I(M_this_ppu_map_addr_7));
    Odrv4 I__2725 (
            .O(N__16739),
            .I(M_this_ppu_map_addr_7));
    LocalMux I__2724 (
            .O(N__16736),
            .I(M_this_ppu_map_addr_7));
    Odrv12 I__2723 (
            .O(N__16731),
            .I(M_this_ppu_map_addr_7));
    InMux I__2722 (
            .O(N__16722),
            .I(N__16713));
    InMux I__2721 (
            .O(N__16721),
            .I(N__16713));
    InMux I__2720 (
            .O(N__16720),
            .I(N__16713));
    LocalMux I__2719 (
            .O(N__16713),
            .I(N__16709));
    InMux I__2718 (
            .O(N__16712),
            .I(N__16706));
    Odrv4 I__2717 (
            .O(N__16709),
            .I(\this_ppu.un1_M_vaddress_q_c3 ));
    LocalMux I__2716 (
            .O(N__16706),
            .I(\this_ppu.un1_M_vaddress_q_c3 ));
    CascadeMux I__2715 (
            .O(N__16701),
            .I(N__16698));
    CascadeBuf I__2714 (
            .O(N__16698),
            .I(N__16695));
    CascadeMux I__2713 (
            .O(N__16695),
            .I(N__16692));
    InMux I__2712 (
            .O(N__16692),
            .I(N__16688));
    InMux I__2711 (
            .O(N__16691),
            .I(N__16683));
    LocalMux I__2710 (
            .O(N__16688),
            .I(N__16679));
    CascadeMux I__2709 (
            .O(N__16687),
            .I(N__16676));
    CascadeMux I__2708 (
            .O(N__16686),
            .I(N__16673));
    LocalMux I__2707 (
            .O(N__16683),
            .I(N__16669));
    CascadeMux I__2706 (
            .O(N__16682),
            .I(N__16666));
    Sp12to4 I__2705 (
            .O(N__16679),
            .I(N__16663));
    InMux I__2704 (
            .O(N__16676),
            .I(N__16656));
    InMux I__2703 (
            .O(N__16673),
            .I(N__16656));
    InMux I__2702 (
            .O(N__16672),
            .I(N__16656));
    Span4Mux_v I__2701 (
            .O(N__16669),
            .I(N__16653));
    InMux I__2700 (
            .O(N__16666),
            .I(N__16650));
    Span12Mux_v I__2699 (
            .O(N__16663),
            .I(N__16647));
    LocalMux I__2698 (
            .O(N__16656),
            .I(M_this_ppu_map_addr_5));
    Odrv4 I__2697 (
            .O(N__16653),
            .I(M_this_ppu_map_addr_5));
    LocalMux I__2696 (
            .O(N__16650),
            .I(M_this_ppu_map_addr_5));
    Odrv12 I__2695 (
            .O(N__16647),
            .I(M_this_ppu_map_addr_5));
    CascadeMux I__2694 (
            .O(N__16638),
            .I(N__16635));
    CascadeBuf I__2693 (
            .O(N__16635),
            .I(N__16632));
    CascadeMux I__2692 (
            .O(N__16632),
            .I(N__16629));
    InMux I__2691 (
            .O(N__16629),
            .I(N__16626));
    LocalMux I__2690 (
            .O(N__16626),
            .I(N__16622));
    InMux I__2689 (
            .O(N__16625),
            .I(N__16619));
    Span4Mux_h I__2688 (
            .O(N__16622),
            .I(N__16616));
    LocalMux I__2687 (
            .O(N__16619),
            .I(N__16611));
    Span4Mux_h I__2686 (
            .O(N__16616),
            .I(N__16607));
    InMux I__2685 (
            .O(N__16615),
            .I(N__16602));
    InMux I__2684 (
            .O(N__16614),
            .I(N__16602));
    Span4Mux_v I__2683 (
            .O(N__16611),
            .I(N__16599));
    InMux I__2682 (
            .O(N__16610),
            .I(N__16596));
    Span4Mux_v I__2681 (
            .O(N__16607),
            .I(N__16593));
    LocalMux I__2680 (
            .O(N__16602),
            .I(M_this_ppu_map_addr_6));
    Odrv4 I__2679 (
            .O(N__16599),
            .I(M_this_ppu_map_addr_6));
    LocalMux I__2678 (
            .O(N__16596),
            .I(M_this_ppu_map_addr_6));
    Odrv4 I__2677 (
            .O(N__16593),
            .I(M_this_ppu_map_addr_6));
    SRMux I__2676 (
            .O(N__16584),
            .I(N__16579));
    SRMux I__2675 (
            .O(N__16583),
            .I(N__16576));
    SRMux I__2674 (
            .O(N__16582),
            .I(N__16573));
    LocalMux I__2673 (
            .O(N__16579),
            .I(N__16570));
    LocalMux I__2672 (
            .O(N__16576),
            .I(N__16567));
    LocalMux I__2671 (
            .O(N__16573),
            .I(N__16564));
    Span4Mux_v I__2670 (
            .O(N__16570),
            .I(N__16561));
    Span4Mux_v I__2669 (
            .O(N__16567),
            .I(N__16558));
    Span4Mux_h I__2668 (
            .O(N__16564),
            .I(N__16555));
    Odrv4 I__2667 (
            .O(N__16561),
            .I(\this_ppu.M_state_q_RNIELANCZ0Z_0 ));
    Odrv4 I__2666 (
            .O(N__16558),
            .I(\this_ppu.M_state_q_RNIELANCZ0Z_0 ));
    Odrv4 I__2665 (
            .O(N__16555),
            .I(\this_ppu.M_state_q_RNIELANCZ0Z_0 ));
    IoInMux I__2664 (
            .O(N__16548),
            .I(N__16545));
    LocalMux I__2663 (
            .O(N__16545),
            .I(N__16542));
    Span12Mux_s5_h I__2662 (
            .O(N__16542),
            .I(N__16538));
    InMux I__2661 (
            .O(N__16541),
            .I(N__16535));
    Span12Mux_h I__2660 (
            .O(N__16538),
            .I(N__16532));
    LocalMux I__2659 (
            .O(N__16535),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI4KCU6Z0Z_9 ));
    Odrv12 I__2658 (
            .O(N__16532),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI4KCU6Z0Z_9 ));
    CascadeMux I__2657 (
            .O(N__16527),
            .I(\this_vga_signals.g1_2_0_0_cascade_ ));
    CascadeMux I__2656 (
            .O(N__16524),
            .I(M_this_state_q_ns_17_cascade_));
    CEMux I__2655 (
            .O(N__16521),
            .I(N__16517));
    CEMux I__2654 (
            .O(N__16520),
            .I(N__16513));
    LocalMux I__2653 (
            .O(N__16517),
            .I(N__16509));
    CEMux I__2652 (
            .O(N__16516),
            .I(N__16506));
    LocalMux I__2651 (
            .O(N__16513),
            .I(N__16503));
    CEMux I__2650 (
            .O(N__16512),
            .I(N__16500));
    Span4Mux_v I__2649 (
            .O(N__16509),
            .I(N__16494));
    LocalMux I__2648 (
            .O(N__16506),
            .I(N__16494));
    Span4Mux_v I__2647 (
            .O(N__16503),
            .I(N__16489));
    LocalMux I__2646 (
            .O(N__16500),
            .I(N__16489));
    CEMux I__2645 (
            .O(N__16499),
            .I(N__16486));
    Span4Mux_h I__2644 (
            .O(N__16494),
            .I(N__16483));
    Span4Mux_h I__2643 (
            .O(N__16489),
            .I(N__16480));
    LocalMux I__2642 (
            .O(N__16486),
            .I(N__16477));
    Odrv4 I__2641 (
            .O(N__16483),
            .I(M_this_state_q_ns_0_17));
    Odrv4 I__2640 (
            .O(N__16480),
            .I(M_this_state_q_ns_0_17));
    Odrv12 I__2639 (
            .O(N__16477),
            .I(M_this_state_q_ns_0_17));
    CascadeMux I__2638 (
            .O(N__16470),
            .I(N__16467));
    InMux I__2637 (
            .O(N__16467),
            .I(N__16464));
    LocalMux I__2636 (
            .O(N__16464),
            .I(N__16461));
    Span4Mux_v I__2635 (
            .O(N__16461),
            .I(N__16458));
    Sp12to4 I__2634 (
            .O(N__16458),
            .I(N__16455));
    Span12Mux_h I__2633 (
            .O(N__16455),
            .I(N__16452));
    Odrv12 I__2632 (
            .O(N__16452),
            .I(M_this_map_ram_read_data_6));
    InMux I__2631 (
            .O(N__16449),
            .I(N__16445));
    InMux I__2630 (
            .O(N__16448),
            .I(N__16442));
    LocalMux I__2629 (
            .O(N__16445),
            .I(N__16437));
    LocalMux I__2628 (
            .O(N__16442),
            .I(N__16437));
    Span4Mux_h I__2627 (
            .O(N__16437),
            .I(N__16434));
    Span4Mux_h I__2626 (
            .O(N__16434),
            .I(N__16431));
    Odrv4 I__2625 (
            .O(N__16431),
            .I(M_this_oam_ram_read_data_8));
    InMux I__2624 (
            .O(N__16428),
            .I(N__16425));
    LocalMux I__2623 (
            .O(N__16425),
            .I(\this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ));
    InMux I__2622 (
            .O(N__16422),
            .I(N__16419));
    LocalMux I__2621 (
            .O(N__16419),
            .I(M_this_oam_ram_read_data_i_9));
    InMux I__2620 (
            .O(N__16416),
            .I(N__16413));
    LocalMux I__2619 (
            .O(N__16413),
            .I(\this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5BZ0 ));
    InMux I__2618 (
            .O(N__16410),
            .I(\this_ppu.un10_sprites_addr_cry_0 ));
    InMux I__2617 (
            .O(N__16407),
            .I(N__16404));
    LocalMux I__2616 (
            .O(N__16404),
            .I(N__16401));
    Span4Mux_h I__2615 (
            .O(N__16401),
            .I(N__16398));
    Span4Mux_h I__2614 (
            .O(N__16398),
            .I(N__16395));
    Odrv4 I__2613 (
            .O(N__16395),
            .I(M_this_oam_ram_read_data_i_10));
    InMux I__2612 (
            .O(N__16392),
            .I(\this_ppu.un10_sprites_addr_cry_1 ));
    InMux I__2611 (
            .O(N__16389),
            .I(N__16386));
    LocalMux I__2610 (
            .O(N__16386),
            .I(N__16383));
    Span4Mux_h I__2609 (
            .O(N__16383),
            .I(N__16380));
    Span4Mux_h I__2608 (
            .O(N__16380),
            .I(N__16377));
    Odrv4 I__2607 (
            .O(N__16377),
            .I(M_this_oam_ram_read_data_i_11));
    InMux I__2606 (
            .O(N__16374),
            .I(\this_ppu.un10_sprites_addr_cry_2 ));
    CascadeMux I__2605 (
            .O(N__16371),
            .I(N__16368));
    InMux I__2604 (
            .O(N__16368),
            .I(N__16365));
    LocalMux I__2603 (
            .O(N__16365),
            .I(N__16362));
    Span4Mux_h I__2602 (
            .O(N__16362),
            .I(N__16359));
    Span4Mux_h I__2601 (
            .O(N__16359),
            .I(N__16356));
    Odrv4 I__2600 (
            .O(N__16356),
            .I(M_this_oam_ram_read_data_i_12));
    InMux I__2599 (
            .O(N__16353),
            .I(N__16350));
    LocalMux I__2598 (
            .O(N__16350),
            .I(\this_ppu.un10_sprites_addr_cry_3_c_RNISS8BZ0 ));
    InMux I__2597 (
            .O(N__16347),
            .I(\this_ppu.un10_sprites_addr_cry_3 ));
    InMux I__2596 (
            .O(N__16344),
            .I(N__16341));
    LocalMux I__2595 (
            .O(N__16341),
            .I(N__16338));
    Span4Mux_v I__2594 (
            .O(N__16338),
            .I(N__16335));
    Span4Mux_h I__2593 (
            .O(N__16335),
            .I(N__16332));
    Odrv4 I__2592 (
            .O(N__16332),
            .I(M_this_oam_ram_read_data_13));
    InMux I__2591 (
            .O(N__16329),
            .I(\this_ppu.un10_sprites_addr_cry_4 ));
    InMux I__2590 (
            .O(N__16326),
            .I(N__16323));
    LocalMux I__2589 (
            .O(N__16323),
            .I(\this_reset_cond.M_stage_qZ0Z_6 ));
    InMux I__2588 (
            .O(N__16320),
            .I(N__16305));
    InMux I__2587 (
            .O(N__16319),
            .I(N__16305));
    InMux I__2586 (
            .O(N__16318),
            .I(N__16305));
    InMux I__2585 (
            .O(N__16317),
            .I(N__16305));
    InMux I__2584 (
            .O(N__16316),
            .I(N__16305));
    LocalMux I__2583 (
            .O(N__16305),
            .I(N__16299));
    InMux I__2582 (
            .O(N__16304),
            .I(N__16294));
    InMux I__2581 (
            .O(N__16303),
            .I(N__16294));
    InMux I__2580 (
            .O(N__16302),
            .I(N__16290));
    Span4Mux_v I__2579 (
            .O(N__16299),
            .I(N__16287));
    LocalMux I__2578 (
            .O(N__16294),
            .I(N__16284));
    InMux I__2577 (
            .O(N__16293),
            .I(N__16281));
    LocalMux I__2576 (
            .O(N__16290),
            .I(N__16277));
    Span4Mux_v I__2575 (
            .O(N__16287),
            .I(N__16270));
    Span4Mux_h I__2574 (
            .O(N__16284),
            .I(N__16270));
    LocalMux I__2573 (
            .O(N__16281),
            .I(N__16270));
    InMux I__2572 (
            .O(N__16280),
            .I(N__16267));
    Span4Mux_h I__2571 (
            .O(N__16277),
            .I(N__16264));
    Span4Mux_v I__2570 (
            .O(N__16270),
            .I(N__16261));
    LocalMux I__2569 (
            .O(N__16267),
            .I(N__16258));
    Span4Mux_v I__2568 (
            .O(N__16264),
            .I(N__16255));
    Span4Mux_v I__2567 (
            .O(N__16261),
            .I(N__16252));
    Span12Mux_h I__2566 (
            .O(N__16258),
            .I(N__16249));
    Span4Mux_v I__2565 (
            .O(N__16255),
            .I(N__16246));
    Span4Mux_v I__2564 (
            .O(N__16252),
            .I(N__16243));
    Span12Mux_v I__2563 (
            .O(N__16249),
            .I(N__16240));
    Span4Mux_v I__2562 (
            .O(N__16246),
            .I(N__16237));
    IoSpan4Mux I__2561 (
            .O(N__16243),
            .I(N__16234));
    Odrv12 I__2560 (
            .O(N__16240),
            .I(rst_n_c));
    Odrv4 I__2559 (
            .O(N__16237),
            .I(rst_n_c));
    Odrv4 I__2558 (
            .O(N__16234),
            .I(rst_n_c));
    InMux I__2557 (
            .O(N__16227),
            .I(N__16224));
    LocalMux I__2556 (
            .O(N__16224),
            .I(\this_reset_cond.M_stage_qZ0Z_7 ));
    InMux I__2555 (
            .O(N__16221),
            .I(N__16218));
    LocalMux I__2554 (
            .O(N__16218),
            .I(\this_reset_cond.M_stage_qZ0Z_8 ));
    CascadeMux I__2553 (
            .O(N__16215),
            .I(N__16212));
    InMux I__2552 (
            .O(N__16212),
            .I(N__16209));
    LocalMux I__2551 (
            .O(N__16209),
            .I(\this_vga_signals.vaddress_ac0_9_0_a0_2 ));
    InMux I__2550 (
            .O(N__16206),
            .I(N__16202));
    InMux I__2549 (
            .O(N__16205),
            .I(N__16199));
    LocalMux I__2548 (
            .O(N__16202),
            .I(N__16192));
    LocalMux I__2547 (
            .O(N__16199),
            .I(N__16192));
    InMux I__2546 (
            .O(N__16198),
            .I(N__16189));
    InMux I__2545 (
            .O(N__16197),
            .I(N__16186));
    Span4Mux_v I__2544 (
            .O(N__16192),
            .I(N__16183));
    LocalMux I__2543 (
            .O(N__16189),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    LocalMux I__2542 (
            .O(N__16186),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    Odrv4 I__2541 (
            .O(N__16183),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    InMux I__2540 (
            .O(N__16176),
            .I(N__16172));
    InMux I__2539 (
            .O(N__16175),
            .I(N__16169));
    LocalMux I__2538 (
            .O(N__16172),
            .I(N__16166));
    LocalMux I__2537 (
            .O(N__16169),
            .I(N__16163));
    Odrv4 I__2536 (
            .O(N__16166),
            .I(\this_ppu.un1_M_vaddress_q_c5 ));
    Odrv4 I__2535 (
            .O(N__16163),
            .I(\this_ppu.un1_M_vaddress_q_c5 ));
    InMux I__2534 (
            .O(N__16158),
            .I(N__16154));
    CascadeMux I__2533 (
            .O(N__16157),
            .I(N__16151));
    LocalMux I__2532 (
            .O(N__16154),
            .I(N__16148));
    InMux I__2531 (
            .O(N__16151),
            .I(N__16145));
    Span4Mux_v I__2530 (
            .O(N__16148),
            .I(N__16142));
    LocalMux I__2529 (
            .O(N__16145),
            .I(\this_ppu.M_vaddress_qZ0Z_7 ));
    Odrv4 I__2528 (
            .O(N__16142),
            .I(\this_ppu.M_vaddress_qZ0Z_7 ));
    IoInMux I__2527 (
            .O(N__16137),
            .I(N__16132));
    IoInMux I__2526 (
            .O(N__16136),
            .I(N__16127));
    IoInMux I__2525 (
            .O(N__16135),
            .I(N__16124));
    LocalMux I__2524 (
            .O(N__16132),
            .I(N__16117));
    IoInMux I__2523 (
            .O(N__16131),
            .I(N__16114));
    IoInMux I__2522 (
            .O(N__16130),
            .I(N__16109));
    LocalMux I__2521 (
            .O(N__16127),
            .I(N__16104));
    LocalMux I__2520 (
            .O(N__16124),
            .I(N__16104));
    IoInMux I__2519 (
            .O(N__16123),
            .I(N__16101));
    IoInMux I__2518 (
            .O(N__16122),
            .I(N__16098));
    IoInMux I__2517 (
            .O(N__16121),
            .I(N__16095));
    IoInMux I__2516 (
            .O(N__16120),
            .I(N__16092));
    IoSpan4Mux I__2515 (
            .O(N__16117),
            .I(N__16086));
    LocalMux I__2514 (
            .O(N__16114),
            .I(N__16086));
    IoInMux I__2513 (
            .O(N__16113),
            .I(N__16083));
    IoInMux I__2512 (
            .O(N__16112),
            .I(N__16080));
    LocalMux I__2511 (
            .O(N__16109),
            .I(N__16076));
    IoSpan4Mux I__2510 (
            .O(N__16104),
            .I(N__16073));
    LocalMux I__2509 (
            .O(N__16101),
            .I(N__16064));
    LocalMux I__2508 (
            .O(N__16098),
            .I(N__16064));
    LocalMux I__2507 (
            .O(N__16095),
            .I(N__16064));
    LocalMux I__2506 (
            .O(N__16092),
            .I(N__16064));
    IoInMux I__2505 (
            .O(N__16091),
            .I(N__16061));
    IoSpan4Mux I__2504 (
            .O(N__16086),
            .I(N__16056));
    LocalMux I__2503 (
            .O(N__16083),
            .I(N__16056));
    LocalMux I__2502 (
            .O(N__16080),
            .I(N__16053));
    IoInMux I__2501 (
            .O(N__16079),
            .I(N__16050));
    IoSpan4Mux I__2500 (
            .O(N__16076),
            .I(N__16045));
    IoSpan4Mux I__2499 (
            .O(N__16073),
            .I(N__16042));
    IoSpan4Mux I__2498 (
            .O(N__16064),
            .I(N__16037));
    LocalMux I__2497 (
            .O(N__16061),
            .I(N__16037));
    IoSpan4Mux I__2496 (
            .O(N__16056),
            .I(N__16030));
    IoSpan4Mux I__2495 (
            .O(N__16053),
            .I(N__16030));
    LocalMux I__2494 (
            .O(N__16050),
            .I(N__16030));
    IoInMux I__2493 (
            .O(N__16049),
            .I(N__16027));
    IoInMux I__2492 (
            .O(N__16048),
            .I(N__16024));
    IoSpan4Mux I__2491 (
            .O(N__16045),
            .I(N__16021));
    IoSpan4Mux I__2490 (
            .O(N__16042),
            .I(N__16016));
    IoSpan4Mux I__2489 (
            .O(N__16037),
            .I(N__16016));
    IoSpan4Mux I__2488 (
            .O(N__16030),
            .I(N__16012));
    LocalMux I__2487 (
            .O(N__16027),
            .I(N__16008));
    LocalMux I__2486 (
            .O(N__16024),
            .I(N__16005));
    Span4Mux_s2_h I__2485 (
            .O(N__16021),
            .I(N__16002));
    Span4Mux_s1_h I__2484 (
            .O(N__16016),
            .I(N__15999));
    IoInMux I__2483 (
            .O(N__16015),
            .I(N__15996));
    Span4Mux_s2_v I__2482 (
            .O(N__16012),
            .I(N__15993));
    IoInMux I__2481 (
            .O(N__16011),
            .I(N__15990));
    Span12Mux_s6_h I__2480 (
            .O(N__16008),
            .I(N__15985));
    Span12Mux_s4_v I__2479 (
            .O(N__16005),
            .I(N__15985));
    Sp12to4 I__2478 (
            .O(N__16002),
            .I(N__15982));
    Sp12to4 I__2477 (
            .O(N__15999),
            .I(N__15977));
    LocalMux I__2476 (
            .O(N__15996),
            .I(N__15977));
    Sp12to4 I__2475 (
            .O(N__15993),
            .I(N__15972));
    LocalMux I__2474 (
            .O(N__15990),
            .I(N__15972));
    Span12Mux_v I__2473 (
            .O(N__15985),
            .I(N__15965));
    Span12Mux_h I__2472 (
            .O(N__15982),
            .I(N__15965));
    Span12Mux_s6_h I__2471 (
            .O(N__15977),
            .I(N__15965));
    Span12Mux_s10_v I__2470 (
            .O(N__15972),
            .I(N__15962));
    Odrv12 I__2469 (
            .O(N__15965),
            .I(dma_0_i));
    Odrv12 I__2468 (
            .O(N__15962),
            .I(dma_0_i));
    CEMux I__2467 (
            .O(N__15957),
            .I(N__15954));
    LocalMux I__2466 (
            .O(N__15954),
            .I(N__15951));
    Span4Mux_v I__2465 (
            .O(N__15951),
            .I(N__15948));
    Span4Mux_h I__2464 (
            .O(N__15948),
            .I(N__15944));
    CEMux I__2463 (
            .O(N__15947),
            .I(N__15941));
    Odrv4 I__2462 (
            .O(N__15944),
            .I(N_1430_0));
    LocalMux I__2461 (
            .O(N__15941),
            .I(N_1430_0));
    CascadeMux I__2460 (
            .O(N__15936),
            .I(\this_vga_signals.N_1028_cascade_ ));
    InMux I__2459 (
            .O(N__15933),
            .I(N__15929));
    InMux I__2458 (
            .O(N__15932),
            .I(N__15926));
    LocalMux I__2457 (
            .O(N__15929),
            .I(\this_vga_signals.N_999 ));
    LocalMux I__2456 (
            .O(N__15926),
            .I(\this_vga_signals.N_999 ));
    CascadeMux I__2455 (
            .O(N__15921),
            .I(\this_vga_signals.N_1004_cascade_ ));
    CascadeMux I__2454 (
            .O(N__15918),
            .I(N__15915));
    InMux I__2453 (
            .O(N__15915),
            .I(N__15912));
    LocalMux I__2452 (
            .O(N__15912),
            .I(\this_vga_signals.N_1013 ));
    CascadeMux I__2451 (
            .O(N__15909),
            .I(\this_vga_signals.N_1013_cascade_ ));
    CascadeMux I__2450 (
            .O(N__15906),
            .I(\this_vga_signals.N_105_mux_cascade_ ));
    InMux I__2449 (
            .O(N__15903),
            .I(N__15899));
    InMux I__2448 (
            .O(N__15902),
            .I(N__15896));
    LocalMux I__2447 (
            .O(N__15899),
            .I(\this_vga_signals.N_113_mux ));
    LocalMux I__2446 (
            .O(N__15896),
            .I(\this_vga_signals.N_113_mux ));
    InMux I__2445 (
            .O(N__15891),
            .I(N__15888));
    LocalMux I__2444 (
            .O(N__15888),
            .I(\this_reset_cond.M_stage_qZ0Z_4 ));
    InMux I__2443 (
            .O(N__15885),
            .I(N__15882));
    LocalMux I__2442 (
            .O(N__15882),
            .I(\this_reset_cond.M_stage_qZ0Z_5 ));
    InMux I__2441 (
            .O(N__15879),
            .I(N__15876));
    LocalMux I__2440 (
            .O(N__15876),
            .I(N__15873));
    Span4Mux_v I__2439 (
            .O(N__15873),
            .I(N__15869));
    InMux I__2438 (
            .O(N__15872),
            .I(N__15866));
    Span4Mux_v I__2437 (
            .O(N__15869),
            .I(N__15862));
    LocalMux I__2436 (
            .O(N__15866),
            .I(N__15859));
    CascadeMux I__2435 (
            .O(N__15865),
            .I(N__15856));
    Span4Mux_v I__2434 (
            .O(N__15862),
            .I(N__15851));
    Span4Mux_v I__2433 (
            .O(N__15859),
            .I(N__15851));
    InMux I__2432 (
            .O(N__15856),
            .I(N__15847));
    Sp12to4 I__2431 (
            .O(N__15851),
            .I(N__15844));
    InMux I__2430 (
            .O(N__15850),
            .I(N__15841));
    LocalMux I__2429 (
            .O(N__15847),
            .I(N__15838));
    Span12Mux_h I__2428 (
            .O(N__15844),
            .I(N__15835));
    LocalMux I__2427 (
            .O(N__15841),
            .I(N__15832));
    Span4Mux_v I__2426 (
            .O(N__15838),
            .I(N__15829));
    Odrv12 I__2425 (
            .O(N__15835),
            .I(this_vga_signals_vvisibility));
    Odrv4 I__2424 (
            .O(N__15832),
            .I(this_vga_signals_vvisibility));
    Odrv4 I__2423 (
            .O(N__15829),
            .I(this_vga_signals_vvisibility));
    InMux I__2422 (
            .O(N__15822),
            .I(N__15818));
    CascadeMux I__2421 (
            .O(N__15821),
            .I(N__15811));
    LocalMux I__2420 (
            .O(N__15818),
            .I(N__15806));
    InMux I__2419 (
            .O(N__15817),
            .I(N__15803));
    InMux I__2418 (
            .O(N__15816),
            .I(N__15800));
    InMux I__2417 (
            .O(N__15815),
            .I(N__15797));
    InMux I__2416 (
            .O(N__15814),
            .I(N__15790));
    InMux I__2415 (
            .O(N__15811),
            .I(N__15790));
    InMux I__2414 (
            .O(N__15810),
            .I(N__15790));
    IoInMux I__2413 (
            .O(N__15809),
            .I(N__15787));
    Span4Mux_v I__2412 (
            .O(N__15806),
            .I(N__15782));
    LocalMux I__2411 (
            .O(N__15803),
            .I(N__15782));
    LocalMux I__2410 (
            .O(N__15800),
            .I(N__15779));
    LocalMux I__2409 (
            .O(N__15797),
            .I(N__15774));
    LocalMux I__2408 (
            .O(N__15790),
            .I(N__15774));
    LocalMux I__2407 (
            .O(N__15787),
            .I(N__15768));
    Span4Mux_h I__2406 (
            .O(N__15782),
            .I(N__15765));
    Span4Mux_v I__2405 (
            .O(N__15779),
            .I(N__15760));
    Span4Mux_v I__2404 (
            .O(N__15774),
            .I(N__15760));
    InMux I__2403 (
            .O(N__15773),
            .I(N__15757));
    InMux I__2402 (
            .O(N__15772),
            .I(N__15754));
    InMux I__2401 (
            .O(N__15771),
            .I(N__15751));
    Span4Mux_s3_v I__2400 (
            .O(N__15768),
            .I(N__15748));
    Span4Mux_v I__2399 (
            .O(N__15765),
            .I(N__15745));
    Span4Mux_h I__2398 (
            .O(N__15760),
            .I(N__15736));
    LocalMux I__2397 (
            .O(N__15757),
            .I(N__15736));
    LocalMux I__2396 (
            .O(N__15754),
            .I(N__15736));
    LocalMux I__2395 (
            .O(N__15751),
            .I(N__15736));
    Span4Mux_v I__2394 (
            .O(N__15748),
            .I(N__15733));
    Odrv4 I__2393 (
            .O(N__15745),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__2392 (
            .O(N__15736),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__2391 (
            .O(N__15733),
            .I(M_this_reset_cond_out_0));
    InMux I__2390 (
            .O(N__15726),
            .I(N__15723));
    LocalMux I__2389 (
            .O(N__15723),
            .I(N__15720));
    Span4Mux_h I__2388 (
            .O(N__15720),
            .I(N__15717));
    Odrv4 I__2387 (
            .O(N__15717),
            .I(\this_ppu.un3_sprites_addr_cry_2_c_RNIVRCZ0Z8 ));
    CascadeMux I__2386 (
            .O(N__15714),
            .I(N__15711));
    CascadeBuf I__2385 (
            .O(N__15711),
            .I(N__15708));
    CascadeMux I__2384 (
            .O(N__15708),
            .I(N__15705));
    CascadeBuf I__2383 (
            .O(N__15705),
            .I(N__15702));
    CascadeMux I__2382 (
            .O(N__15702),
            .I(N__15699));
    CascadeBuf I__2381 (
            .O(N__15699),
            .I(N__15696));
    CascadeMux I__2380 (
            .O(N__15696),
            .I(N__15693));
    CascadeBuf I__2379 (
            .O(N__15693),
            .I(N__15690));
    CascadeMux I__2378 (
            .O(N__15690),
            .I(N__15687));
    CascadeBuf I__2377 (
            .O(N__15687),
            .I(N__15684));
    CascadeMux I__2376 (
            .O(N__15684),
            .I(N__15681));
    CascadeBuf I__2375 (
            .O(N__15681),
            .I(N__15678));
    CascadeMux I__2374 (
            .O(N__15678),
            .I(N__15675));
    CascadeBuf I__2373 (
            .O(N__15675),
            .I(N__15672));
    CascadeMux I__2372 (
            .O(N__15672),
            .I(N__15669));
    CascadeBuf I__2371 (
            .O(N__15669),
            .I(N__15666));
    CascadeMux I__2370 (
            .O(N__15666),
            .I(N__15663));
    CascadeBuf I__2369 (
            .O(N__15663),
            .I(N__15660));
    CascadeMux I__2368 (
            .O(N__15660),
            .I(N__15657));
    CascadeBuf I__2367 (
            .O(N__15657),
            .I(N__15654));
    CascadeMux I__2366 (
            .O(N__15654),
            .I(N__15651));
    CascadeBuf I__2365 (
            .O(N__15651),
            .I(N__15648));
    CascadeMux I__2364 (
            .O(N__15648),
            .I(N__15645));
    CascadeBuf I__2363 (
            .O(N__15645),
            .I(N__15642));
    CascadeMux I__2362 (
            .O(N__15642),
            .I(N__15639));
    CascadeBuf I__2361 (
            .O(N__15639),
            .I(N__15636));
    CascadeMux I__2360 (
            .O(N__15636),
            .I(N__15633));
    CascadeBuf I__2359 (
            .O(N__15633),
            .I(N__15630));
    CascadeMux I__2358 (
            .O(N__15630),
            .I(N__15627));
    CascadeBuf I__2357 (
            .O(N__15627),
            .I(N__15624));
    CascadeMux I__2356 (
            .O(N__15624),
            .I(N__15621));
    InMux I__2355 (
            .O(N__15621),
            .I(N__15618));
    LocalMux I__2354 (
            .O(N__15618),
            .I(N__15615));
    Span12Mux_h I__2353 (
            .O(N__15615),
            .I(N__15612));
    Span12Mux_v I__2352 (
            .O(N__15612),
            .I(N__15609));
    Odrv12 I__2351 (
            .O(N__15609),
            .I(M_this_ppu_sprites_addr_3));
    InMux I__2350 (
            .O(N__15606),
            .I(N__15603));
    LocalMux I__2349 (
            .O(N__15603),
            .I(N__15600));
    Span4Mux_h I__2348 (
            .O(N__15600),
            .I(N__15597));
    Span4Mux_h I__2347 (
            .O(N__15597),
            .I(N__15594));
    Odrv4 I__2346 (
            .O(N__15594),
            .I(\this_oam_ram.M_this_oam_ram_read_data_9 ));
    CascadeMux I__2345 (
            .O(N__15591),
            .I(N__15588));
    InMux I__2344 (
            .O(N__15588),
            .I(N__15585));
    LocalMux I__2343 (
            .O(N__15585),
            .I(N__15582));
    Span4Mux_v I__2342 (
            .O(N__15582),
            .I(N__15579));
    Span4Mux_h I__2341 (
            .O(N__15579),
            .I(N__15576));
    Span4Mux_h I__2340 (
            .O(N__15576),
            .I(N__15573));
    Odrv4 I__2339 (
            .O(N__15573),
            .I(M_this_map_ram_read_data_3));
    CascadeMux I__2338 (
            .O(N__15570),
            .I(N__15567));
    CascadeBuf I__2337 (
            .O(N__15567),
            .I(N__15564));
    CascadeMux I__2336 (
            .O(N__15564),
            .I(N__15561));
    CascadeBuf I__2335 (
            .O(N__15561),
            .I(N__15558));
    CascadeMux I__2334 (
            .O(N__15558),
            .I(N__15555));
    CascadeBuf I__2333 (
            .O(N__15555),
            .I(N__15552));
    CascadeMux I__2332 (
            .O(N__15552),
            .I(N__15549));
    CascadeBuf I__2331 (
            .O(N__15549),
            .I(N__15546));
    CascadeMux I__2330 (
            .O(N__15546),
            .I(N__15543));
    CascadeBuf I__2329 (
            .O(N__15543),
            .I(N__15540));
    CascadeMux I__2328 (
            .O(N__15540),
            .I(N__15537));
    CascadeBuf I__2327 (
            .O(N__15537),
            .I(N__15534));
    CascadeMux I__2326 (
            .O(N__15534),
            .I(N__15531));
    CascadeBuf I__2325 (
            .O(N__15531),
            .I(N__15528));
    CascadeMux I__2324 (
            .O(N__15528),
            .I(N__15525));
    CascadeBuf I__2323 (
            .O(N__15525),
            .I(N__15522));
    CascadeMux I__2322 (
            .O(N__15522),
            .I(N__15519));
    CascadeBuf I__2321 (
            .O(N__15519),
            .I(N__15516));
    CascadeMux I__2320 (
            .O(N__15516),
            .I(N__15513));
    CascadeBuf I__2319 (
            .O(N__15513),
            .I(N__15510));
    CascadeMux I__2318 (
            .O(N__15510),
            .I(N__15507));
    CascadeBuf I__2317 (
            .O(N__15507),
            .I(N__15504));
    CascadeMux I__2316 (
            .O(N__15504),
            .I(N__15501));
    CascadeBuf I__2315 (
            .O(N__15501),
            .I(N__15498));
    CascadeMux I__2314 (
            .O(N__15498),
            .I(N__15495));
    CascadeBuf I__2313 (
            .O(N__15495),
            .I(N__15492));
    CascadeMux I__2312 (
            .O(N__15492),
            .I(N__15489));
    CascadeBuf I__2311 (
            .O(N__15489),
            .I(N__15486));
    CascadeMux I__2310 (
            .O(N__15486),
            .I(N__15483));
    CascadeBuf I__2309 (
            .O(N__15483),
            .I(N__15480));
    CascadeMux I__2308 (
            .O(N__15480),
            .I(N__15477));
    InMux I__2307 (
            .O(N__15477),
            .I(N__15474));
    LocalMux I__2306 (
            .O(N__15474),
            .I(N__15471));
    Span4Mux_h I__2305 (
            .O(N__15471),
            .I(N__15468));
    Sp12to4 I__2304 (
            .O(N__15468),
            .I(N__15465));
    Span12Mux_s6_v I__2303 (
            .O(N__15465),
            .I(N__15462));
    Span12Mux_h I__2302 (
            .O(N__15462),
            .I(N__15459));
    Odrv12 I__2301 (
            .O(N__15459),
            .I(M_this_ppu_sprites_addr_9));
    CascadeMux I__2300 (
            .O(N__15456),
            .I(N__15453));
    InMux I__2299 (
            .O(N__15453),
            .I(N__15447));
    InMux I__2298 (
            .O(N__15452),
            .I(N__15447));
    LocalMux I__2297 (
            .O(N__15447),
            .I(\this_ppu.M_state_d_0_sqmuxa_1 ));
    InMux I__2296 (
            .O(N__15444),
            .I(N__15441));
    LocalMux I__2295 (
            .O(N__15441),
            .I(N__15438));
    Odrv4 I__2294 (
            .O(N__15438),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_7 ));
    CascadeMux I__2293 (
            .O(N__15435),
            .I(N__15431));
    InMux I__2292 (
            .O(N__15434),
            .I(N__15428));
    InMux I__2291 (
            .O(N__15431),
            .I(N__15425));
    LocalMux I__2290 (
            .O(N__15428),
            .I(N__15420));
    LocalMux I__2289 (
            .O(N__15425),
            .I(N__15420));
    Odrv4 I__2288 (
            .O(N__15420),
            .I(\this_ppu.M_count_qZ0Z_7 ));
    CascadeMux I__2287 (
            .O(N__15417),
            .I(N__15414));
    InMux I__2286 (
            .O(N__15414),
            .I(N__15411));
    LocalMux I__2285 (
            .O(N__15411),
            .I(\this_vga_signals.N_129_mux ));
    InMux I__2284 (
            .O(N__15408),
            .I(N__15405));
    LocalMux I__2283 (
            .O(N__15405),
            .I(\this_vga_signals.N_1028 ));
    InMux I__2282 (
            .O(N__15402),
            .I(N__15399));
    LocalMux I__2281 (
            .O(N__15399),
            .I(M_this_data_tmp_qZ0Z_10));
    InMux I__2280 (
            .O(N__15396),
            .I(N__15393));
    LocalMux I__2279 (
            .O(N__15393),
            .I(N__15390));
    Span4Mux_h I__2278 (
            .O(N__15390),
            .I(N__15387));
    Odrv4 I__2277 (
            .O(N__15387),
            .I(M_this_data_tmp_qZ0Z_17));
    CascadeMux I__2276 (
            .O(N__15384),
            .I(N__15381));
    InMux I__2275 (
            .O(N__15381),
            .I(N__15378));
    LocalMux I__2274 (
            .O(N__15378),
            .I(\this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ));
    InMux I__2273 (
            .O(N__15375),
            .I(N__15370));
    InMux I__2272 (
            .O(N__15374),
            .I(N__15367));
    InMux I__2271 (
            .O(N__15373),
            .I(N__15364));
    LocalMux I__2270 (
            .O(N__15370),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    LocalMux I__2269 (
            .O(N__15367),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    LocalMux I__2268 (
            .O(N__15364),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    InMux I__2267 (
            .O(N__15357),
            .I(N__15352));
    InMux I__2266 (
            .O(N__15356),
            .I(N__15349));
    InMux I__2265 (
            .O(N__15355),
            .I(N__15346));
    LocalMux I__2264 (
            .O(N__15352),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    LocalMux I__2263 (
            .O(N__15349),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    LocalMux I__2262 (
            .O(N__15346),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    CascadeMux I__2261 (
            .O(N__15339),
            .I(N__15336));
    InMux I__2260 (
            .O(N__15336),
            .I(N__15333));
    LocalMux I__2259 (
            .O(N__15333),
            .I(\this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ));
    CascadeMux I__2258 (
            .O(N__15330),
            .I(N__15327));
    InMux I__2257 (
            .O(N__15327),
            .I(N__15322));
    InMux I__2256 (
            .O(N__15326),
            .I(N__15317));
    InMux I__2255 (
            .O(N__15325),
            .I(N__15317));
    LocalMux I__2254 (
            .O(N__15322),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    LocalMux I__2253 (
            .O(N__15317),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    InMux I__2252 (
            .O(N__15312),
            .I(N__15309));
    LocalMux I__2251 (
            .O(N__15309),
            .I(N__15306));
    Span4Mux_h I__2250 (
            .O(N__15306),
            .I(N__15303));
    Span4Mux_v I__2249 (
            .O(N__15303),
            .I(N__15300));
    Span4Mux_h I__2248 (
            .O(N__15300),
            .I(N__15297));
    Odrv4 I__2247 (
            .O(N__15297),
            .I(M_this_map_ram_read_data_2));
    CascadeMux I__2246 (
            .O(N__15294),
            .I(\this_ppu.un10_sprites_addr_axb_0_cascade_ ));
    CascadeMux I__2245 (
            .O(N__15291),
            .I(N__15288));
    CascadeBuf I__2244 (
            .O(N__15288),
            .I(N__15285));
    CascadeMux I__2243 (
            .O(N__15285),
            .I(N__15282));
    CascadeBuf I__2242 (
            .O(N__15282),
            .I(N__15279));
    CascadeMux I__2241 (
            .O(N__15279),
            .I(N__15276));
    CascadeBuf I__2240 (
            .O(N__15276),
            .I(N__15273));
    CascadeMux I__2239 (
            .O(N__15273),
            .I(N__15270));
    CascadeBuf I__2238 (
            .O(N__15270),
            .I(N__15267));
    CascadeMux I__2237 (
            .O(N__15267),
            .I(N__15264));
    CascadeBuf I__2236 (
            .O(N__15264),
            .I(N__15261));
    CascadeMux I__2235 (
            .O(N__15261),
            .I(N__15258));
    CascadeBuf I__2234 (
            .O(N__15258),
            .I(N__15255));
    CascadeMux I__2233 (
            .O(N__15255),
            .I(N__15252));
    CascadeBuf I__2232 (
            .O(N__15252),
            .I(N__15249));
    CascadeMux I__2231 (
            .O(N__15249),
            .I(N__15246));
    CascadeBuf I__2230 (
            .O(N__15246),
            .I(N__15243));
    CascadeMux I__2229 (
            .O(N__15243),
            .I(N__15240));
    CascadeBuf I__2228 (
            .O(N__15240),
            .I(N__15237));
    CascadeMux I__2227 (
            .O(N__15237),
            .I(N__15234));
    CascadeBuf I__2226 (
            .O(N__15234),
            .I(N__15231));
    CascadeMux I__2225 (
            .O(N__15231),
            .I(N__15228));
    CascadeBuf I__2224 (
            .O(N__15228),
            .I(N__15225));
    CascadeMux I__2223 (
            .O(N__15225),
            .I(N__15222));
    CascadeBuf I__2222 (
            .O(N__15222),
            .I(N__15219));
    CascadeMux I__2221 (
            .O(N__15219),
            .I(N__15216));
    CascadeBuf I__2220 (
            .O(N__15216),
            .I(N__15213));
    CascadeMux I__2219 (
            .O(N__15213),
            .I(N__15210));
    CascadeBuf I__2218 (
            .O(N__15210),
            .I(N__15207));
    CascadeMux I__2217 (
            .O(N__15207),
            .I(N__15204));
    CascadeBuf I__2216 (
            .O(N__15204),
            .I(N__15201));
    CascadeMux I__2215 (
            .O(N__15201),
            .I(N__15198));
    InMux I__2214 (
            .O(N__15198),
            .I(N__15195));
    LocalMux I__2213 (
            .O(N__15195),
            .I(N__15192));
    Span4Mux_h I__2212 (
            .O(N__15192),
            .I(N__15189));
    Span4Mux_h I__2211 (
            .O(N__15189),
            .I(N__15186));
    Span4Mux_v I__2210 (
            .O(N__15186),
            .I(N__15183));
    Span4Mux_v I__2209 (
            .O(N__15183),
            .I(N__15180));
    Span4Mux_v I__2208 (
            .O(N__15180),
            .I(N__15177));
    Odrv4 I__2207 (
            .O(N__15177),
            .I(M_this_ppu_sprites_addr_8));
    InMux I__2206 (
            .O(N__15174),
            .I(N__15166));
    InMux I__2205 (
            .O(N__15173),
            .I(N__15166));
    CascadeMux I__2204 (
            .O(N__15172),
            .I(N__15162));
    InMux I__2203 (
            .O(N__15171),
            .I(N__15157));
    LocalMux I__2202 (
            .O(N__15166),
            .I(N__15154));
    InMux I__2201 (
            .O(N__15165),
            .I(N__15151));
    InMux I__2200 (
            .O(N__15162),
            .I(N__15144));
    InMux I__2199 (
            .O(N__15161),
            .I(N__15144));
    InMux I__2198 (
            .O(N__15160),
            .I(N__15144));
    LocalMux I__2197 (
            .O(N__15157),
            .I(N__15141));
    Odrv4 I__2196 (
            .O(N__15154),
            .I(\this_ppu.un10_0 ));
    LocalMux I__2195 (
            .O(N__15151),
            .I(\this_ppu.un10_0 ));
    LocalMux I__2194 (
            .O(N__15144),
            .I(\this_ppu.un10_0 ));
    Odrv12 I__2193 (
            .O(N__15141),
            .I(\this_ppu.un10_0 ));
    CascadeMux I__2192 (
            .O(N__15132),
            .I(N__15129));
    InMux I__2191 (
            .O(N__15129),
            .I(N__15126));
    LocalMux I__2190 (
            .O(N__15126),
            .I(N__15123));
    Odrv4 I__2189 (
            .O(N__15123),
            .I(\this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ));
    InMux I__2188 (
            .O(N__15120),
            .I(N__15112));
    InMux I__2187 (
            .O(N__15119),
            .I(N__15107));
    InMux I__2186 (
            .O(N__15118),
            .I(N__15107));
    InMux I__2185 (
            .O(N__15117),
            .I(N__15104));
    InMux I__2184 (
            .O(N__15116),
            .I(N__15099));
    InMux I__2183 (
            .O(N__15115),
            .I(N__15099));
    LocalMux I__2182 (
            .O(N__15112),
            .I(N__15096));
    LocalMux I__2181 (
            .O(N__15107),
            .I(\this_ppu.N_1456_0 ));
    LocalMux I__2180 (
            .O(N__15104),
            .I(\this_ppu.N_1456_0 ));
    LocalMux I__2179 (
            .O(N__15099),
            .I(\this_ppu.N_1456_0 ));
    Odrv4 I__2178 (
            .O(N__15096),
            .I(\this_ppu.N_1456_0 ));
    CascadeMux I__2177 (
            .O(N__15087),
            .I(N__15082));
    CascadeMux I__2176 (
            .O(N__15086),
            .I(N__15079));
    InMux I__2175 (
            .O(N__15085),
            .I(N__15076));
    InMux I__2174 (
            .O(N__15082),
            .I(N__15073));
    InMux I__2173 (
            .O(N__15079),
            .I(N__15070));
    LocalMux I__2172 (
            .O(N__15076),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    LocalMux I__2171 (
            .O(N__15073),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    LocalMux I__2170 (
            .O(N__15070),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    InMux I__2169 (
            .O(N__15063),
            .I(N__15060));
    LocalMux I__2168 (
            .O(N__15060),
            .I(N__15057));
    Odrv12 I__2167 (
            .O(N__15057),
            .I(\this_reset_cond.M_stage_qZ0Z_3 ));
    InMux I__2166 (
            .O(N__15054),
            .I(N__15046));
    InMux I__2165 (
            .O(N__15053),
            .I(N__15046));
    InMux I__2164 (
            .O(N__15052),
            .I(N__15041));
    InMux I__2163 (
            .O(N__15051),
            .I(N__15041));
    LocalMux I__2162 (
            .O(N__15046),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    LocalMux I__2161 (
            .O(N__15041),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    CascadeMux I__2160 (
            .O(N__15036),
            .I(\this_vga_signals.i21_mux_cascade_ ));
    InMux I__2159 (
            .O(N__15033),
            .I(N__15027));
    InMux I__2158 (
            .O(N__15032),
            .I(N__15024));
    InMux I__2157 (
            .O(N__15031),
            .I(N__15019));
    InMux I__2156 (
            .O(N__15030),
            .I(N__15019));
    LocalMux I__2155 (
            .O(N__15027),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    LocalMux I__2154 (
            .O(N__15024),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    LocalMux I__2153 (
            .O(N__15019),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    InMux I__2152 (
            .O(N__15012),
            .I(N__15009));
    LocalMux I__2151 (
            .O(N__15009),
            .I(N__15006));
    Span4Mux_h I__2150 (
            .O(N__15006),
            .I(N__15003));
    Span4Mux_h I__2149 (
            .O(N__15003),
            .I(N__15000));
    Odrv4 I__2148 (
            .O(N__15000),
            .I(N_817_0));
    InMux I__2147 (
            .O(N__14997),
            .I(N__14994));
    LocalMux I__2146 (
            .O(N__14994),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__2145 (
            .O(N__14991),
            .I(N__14988));
    LocalMux I__2144 (
            .O(N__14988),
            .I(\this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ));
    CascadeMux I__2143 (
            .O(N__14985),
            .I(N__14982));
    InMux I__2142 (
            .O(N__14982),
            .I(N__14979));
    LocalMux I__2141 (
            .O(N__14979),
            .I(N__14976));
    Odrv4 I__2140 (
            .O(N__14976),
            .I(\this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ));
    InMux I__2139 (
            .O(N__14973),
            .I(N__14968));
    InMux I__2138 (
            .O(N__14972),
            .I(N__14965));
    InMux I__2137 (
            .O(N__14971),
            .I(N__14962));
    LocalMux I__2136 (
            .O(N__14968),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    LocalMux I__2135 (
            .O(N__14965),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    LocalMux I__2134 (
            .O(N__14962),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    CascadeMux I__2133 (
            .O(N__14955),
            .I(N__14952));
    InMux I__2132 (
            .O(N__14952),
            .I(N__14947));
    InMux I__2131 (
            .O(N__14951),
            .I(N__14942));
    InMux I__2130 (
            .O(N__14950),
            .I(N__14942));
    LocalMux I__2129 (
            .O(N__14947),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    LocalMux I__2128 (
            .O(N__14942),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    InMux I__2127 (
            .O(N__14937),
            .I(N__14932));
    InMux I__2126 (
            .O(N__14936),
            .I(N__14927));
    InMux I__2125 (
            .O(N__14935),
            .I(N__14927));
    LocalMux I__2124 (
            .O(N__14932),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    LocalMux I__2123 (
            .O(N__14927),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    SRMux I__2122 (
            .O(N__14922),
            .I(N__14919));
    LocalMux I__2121 (
            .O(N__14919),
            .I(N__14915));
    SRMux I__2120 (
            .O(N__14918),
            .I(N__14912));
    Span4Mux_v I__2119 (
            .O(N__14915),
            .I(N__14909));
    LocalMux I__2118 (
            .O(N__14912),
            .I(N__14906));
    Odrv4 I__2117 (
            .O(N__14909),
            .I(\this_ppu.M_state_q_RNIE20V4Z0Z_0 ));
    Odrv4 I__2116 (
            .O(N__14906),
            .I(\this_ppu.M_state_q_RNIE20V4Z0Z_0 ));
    CascadeMux I__2115 (
            .O(N__14901),
            .I(M_this_vga_signals_line_clk_0_cascade_));
    CascadeMux I__2114 (
            .O(N__14898),
            .I(\this_ppu.M_state_d_0_sqmuxa_cascade_ ));
    CascadeMux I__2113 (
            .O(N__14895),
            .I(\this_vga_signals.N_1000_cascade_ ));
    InMux I__2112 (
            .O(N__14892),
            .I(\this_ppu.un1_M_count_q_1_cry_1_s1 ));
    InMux I__2111 (
            .O(N__14889),
            .I(\this_ppu.un1_M_count_q_1_cry_2_s1 ));
    InMux I__2110 (
            .O(N__14886),
            .I(\this_ppu.un1_M_count_q_1_cry_3_s1 ));
    InMux I__2109 (
            .O(N__14883),
            .I(\this_ppu.un1_M_count_q_1_cry_4_s1 ));
    InMux I__2108 (
            .O(N__14880),
            .I(\this_ppu.un1_M_count_q_1_cry_5_s1 ));
    InMux I__2107 (
            .O(N__14877),
            .I(\this_ppu.un1_M_count_q_1_cry_6_s1 ));
    CascadeMux I__2106 (
            .O(N__14874),
            .I(\this_ppu.M_state_d_0_sqmuxa_1_cascade_ ));
    InMux I__2105 (
            .O(N__14871),
            .I(N__14868));
    LocalMux I__2104 (
            .O(N__14868),
            .I(\this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ));
    CascadeMux I__2103 (
            .O(N__14865),
            .I(\this_ppu.N_1456_0_cascade_ ));
    CEMux I__2102 (
            .O(N__14862),
            .I(N__14859));
    LocalMux I__2101 (
            .O(N__14859),
            .I(N__14856));
    Odrv4 I__2100 (
            .O(N__14856),
            .I(\this_vga_signals.N_1090_1 ));
    CascadeMux I__2099 (
            .O(N__14853),
            .I(N__14850));
    InMux I__2098 (
            .O(N__14850),
            .I(N__14845));
    InMux I__2097 (
            .O(N__14849),
            .I(N__14842));
    InMux I__2096 (
            .O(N__14848),
            .I(N__14839));
    LocalMux I__2095 (
            .O(N__14845),
            .I(N__14834));
    LocalMux I__2094 (
            .O(N__14842),
            .I(N__14829));
    LocalMux I__2093 (
            .O(N__14839),
            .I(N__14829));
    InMux I__2092 (
            .O(N__14838),
            .I(N__14823));
    InMux I__2091 (
            .O(N__14837),
            .I(N__14823));
    Span4Mux_v I__2090 (
            .O(N__14834),
            .I(N__14818));
    Span4Mux_v I__2089 (
            .O(N__14829),
            .I(N__14818));
    InMux I__2088 (
            .O(N__14828),
            .I(N__14815));
    LocalMux I__2087 (
            .O(N__14823),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    Odrv4 I__2086 (
            .O(N__14818),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__2085 (
            .O(N__14815),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    CascadeMux I__2084 (
            .O(N__14808),
            .I(N__14803));
    CascadeMux I__2083 (
            .O(N__14807),
            .I(N__14800));
    InMux I__2082 (
            .O(N__14806),
            .I(N__14795));
    InMux I__2081 (
            .O(N__14803),
            .I(N__14792));
    InMux I__2080 (
            .O(N__14800),
            .I(N__14789));
    InMux I__2079 (
            .O(N__14799),
            .I(N__14784));
    InMux I__2078 (
            .O(N__14798),
            .I(N__14784));
    LocalMux I__2077 (
            .O(N__14795),
            .I(N__14776));
    LocalMux I__2076 (
            .O(N__14792),
            .I(N__14776));
    LocalMux I__2075 (
            .O(N__14789),
            .I(N__14776));
    LocalMux I__2074 (
            .O(N__14784),
            .I(N__14773));
    InMux I__2073 (
            .O(N__14783),
            .I(N__14769));
    Span4Mux_v I__2072 (
            .O(N__14776),
            .I(N__14766));
    Span4Mux_h I__2071 (
            .O(N__14773),
            .I(N__14763));
    InMux I__2070 (
            .O(N__14772),
            .I(N__14760));
    LocalMux I__2069 (
            .O(N__14769),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__2068 (
            .O(N__14766),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__2067 (
            .O(N__14763),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2066 (
            .O(N__14760),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    SRMux I__2065 (
            .O(N__14751),
            .I(N__14746));
    SRMux I__2064 (
            .O(N__14750),
            .I(N__14743));
    SRMux I__2063 (
            .O(N__14749),
            .I(N__14739));
    LocalMux I__2062 (
            .O(N__14746),
            .I(N__14736));
    LocalMux I__2061 (
            .O(N__14743),
            .I(N__14733));
    InMux I__2060 (
            .O(N__14742),
            .I(N__14730));
    LocalMux I__2059 (
            .O(N__14739),
            .I(G_464));
    Odrv12 I__2058 (
            .O(N__14736),
            .I(G_464));
    Odrv4 I__2057 (
            .O(N__14733),
            .I(G_464));
    LocalMux I__2056 (
            .O(N__14730),
            .I(G_464));
    InMux I__2055 (
            .O(N__14721),
            .I(N__14718));
    LocalMux I__2054 (
            .O(N__14718),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__2053 (
            .O(N__14715),
            .I(N__14712));
    LocalMux I__2052 (
            .O(N__14712),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    InMux I__2051 (
            .O(N__14709),
            .I(N__14706));
    LocalMux I__2050 (
            .O(N__14706),
            .I(N__14703));
    Span4Mux_h I__2049 (
            .O(N__14703),
            .I(N__14700));
    Odrv4 I__2048 (
            .O(N__14700),
            .I(M_this_oam_ram_write_data_10));
    InMux I__2047 (
            .O(N__14697),
            .I(\this_ppu.un1_M_count_q_1_cry_0_s1 ));
    CascadeMux I__2046 (
            .O(N__14694),
            .I(N__14691));
    InMux I__2045 (
            .O(N__14691),
            .I(N__14688));
    LocalMux I__2044 (
            .O(N__14688),
            .I(\this_ppu.M_state_qc_1_3 ));
    InMux I__2043 (
            .O(N__14685),
            .I(N__14682));
    LocalMux I__2042 (
            .O(N__14682),
            .I(N__14679));
    Span4Mux_h I__2041 (
            .O(N__14679),
            .I(N__14676));
    Sp12to4 I__2040 (
            .O(N__14676),
            .I(N__14673));
    Span12Mux_v I__2039 (
            .O(N__14673),
            .I(N__14669));
    InMux I__2038 (
            .O(N__14672),
            .I(N__14666));
    Odrv12 I__2037 (
            .O(N__14669),
            .I(M_this_ppu_vram_data_0));
    LocalMux I__2036 (
            .O(N__14666),
            .I(M_this_ppu_vram_data_0));
    CascadeMux I__2035 (
            .O(N__14661),
            .I(\this_ppu.M_state_qc_1_1_cascade_ ));
    InMux I__2034 (
            .O(N__14658),
            .I(N__14652));
    InMux I__2033 (
            .O(N__14657),
            .I(N__14652));
    LocalMux I__2032 (
            .O(N__14652),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    CascadeMux I__2031 (
            .O(N__14649),
            .I(N__14644));
    CascadeMux I__2030 (
            .O(N__14648),
            .I(N__14641));
    InMux I__2029 (
            .O(N__14647),
            .I(N__14635));
    InMux I__2028 (
            .O(N__14644),
            .I(N__14635));
    InMux I__2027 (
            .O(N__14641),
            .I(N__14632));
    InMux I__2026 (
            .O(N__14640),
            .I(N__14629));
    LocalMux I__2025 (
            .O(N__14635),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    LocalMux I__2024 (
            .O(N__14632),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    LocalMux I__2023 (
            .O(N__14629),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    CascadeMux I__2022 (
            .O(N__14622),
            .I(N__14619));
    InMux I__2021 (
            .O(N__14619),
            .I(N__14614));
    InMux I__2020 (
            .O(N__14618),
            .I(N__14608));
    InMux I__2019 (
            .O(N__14617),
            .I(N__14604));
    LocalMux I__2018 (
            .O(N__14614),
            .I(N__14601));
    CascadeMux I__2017 (
            .O(N__14613),
            .I(N__14596));
    InMux I__2016 (
            .O(N__14612),
            .I(N__14593));
    CascadeMux I__2015 (
            .O(N__14611),
            .I(N__14590));
    LocalMux I__2014 (
            .O(N__14608),
            .I(N__14587));
    InMux I__2013 (
            .O(N__14607),
            .I(N__14584));
    LocalMux I__2012 (
            .O(N__14604),
            .I(N__14579));
    Span4Mux_v I__2011 (
            .O(N__14601),
            .I(N__14579));
    InMux I__2010 (
            .O(N__14600),
            .I(N__14572));
    InMux I__2009 (
            .O(N__14599),
            .I(N__14572));
    InMux I__2008 (
            .O(N__14596),
            .I(N__14572));
    LocalMux I__2007 (
            .O(N__14593),
            .I(N__14569));
    InMux I__2006 (
            .O(N__14590),
            .I(N__14566));
    Odrv4 I__2005 (
            .O(N__14587),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2004 (
            .O(N__14584),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__2003 (
            .O(N__14579),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2002 (
            .O(N__14572),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__2001 (
            .O(N__14569),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2000 (
            .O(N__14566),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__1999 (
            .O(N__14553),
            .I(N__14542));
    InMux I__1998 (
            .O(N__14552),
            .I(N__14542));
    CascadeMux I__1997 (
            .O(N__14551),
            .I(N__14539));
    CascadeMux I__1996 (
            .O(N__14550),
            .I(N__14536));
    CascadeMux I__1995 (
            .O(N__14549),
            .I(N__14532));
    InMux I__1994 (
            .O(N__14548),
            .I(N__14529));
    InMux I__1993 (
            .O(N__14547),
            .I(N__14525));
    LocalMux I__1992 (
            .O(N__14542),
            .I(N__14522));
    InMux I__1991 (
            .O(N__14539),
            .I(N__14512));
    InMux I__1990 (
            .O(N__14536),
            .I(N__14512));
    InMux I__1989 (
            .O(N__14535),
            .I(N__14512));
    InMux I__1988 (
            .O(N__14532),
            .I(N__14512));
    LocalMux I__1987 (
            .O(N__14529),
            .I(N__14509));
    InMux I__1986 (
            .O(N__14528),
            .I(N__14506));
    LocalMux I__1985 (
            .O(N__14525),
            .I(N__14503));
    Span4Mux_h I__1984 (
            .O(N__14522),
            .I(N__14500));
    InMux I__1983 (
            .O(N__14521),
            .I(N__14497));
    LocalMux I__1982 (
            .O(N__14512),
            .I(N__14494));
    Odrv4 I__1981 (
            .O(N__14509),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1980 (
            .O(N__14506),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1979 (
            .O(N__14503),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1978 (
            .O(N__14500),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1977 (
            .O(N__14497),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1976 (
            .O(N__14494),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__1975 (
            .O(N__14481),
            .I(N__14463));
    InMux I__1974 (
            .O(N__14480),
            .I(N__14463));
    InMux I__1973 (
            .O(N__14479),
            .I(N__14463));
    InMux I__1972 (
            .O(N__14478),
            .I(N__14463));
    InMux I__1971 (
            .O(N__14477),
            .I(N__14458));
    InMux I__1970 (
            .O(N__14476),
            .I(N__14458));
    InMux I__1969 (
            .O(N__14475),
            .I(N__14455));
    InMux I__1968 (
            .O(N__14474),
            .I(N__14451));
    InMux I__1967 (
            .O(N__14473),
            .I(N__14448));
    InMux I__1966 (
            .O(N__14472),
            .I(N__14445));
    LocalMux I__1965 (
            .O(N__14463),
            .I(N__14442));
    LocalMux I__1964 (
            .O(N__14458),
            .I(N__14437));
    LocalMux I__1963 (
            .O(N__14455),
            .I(N__14437));
    InMux I__1962 (
            .O(N__14454),
            .I(N__14434));
    LocalMux I__1961 (
            .O(N__14451),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1960 (
            .O(N__14448),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1959 (
            .O(N__14445),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1958 (
            .O(N__14442),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1957 (
            .O(N__14437),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1956 (
            .O(N__14434),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__1955 (
            .O(N__14421),
            .I(N__14413));
    InMux I__1954 (
            .O(N__14420),
            .I(N__14413));
    CascadeMux I__1953 (
            .O(N__14419),
            .I(N__14407));
    CascadeMux I__1952 (
            .O(N__14418),
            .I(N__14403));
    LocalMux I__1951 (
            .O(N__14413),
            .I(N__14398));
    InMux I__1950 (
            .O(N__14412),
            .I(N__14395));
    InMux I__1949 (
            .O(N__14411),
            .I(N__14392));
    InMux I__1948 (
            .O(N__14410),
            .I(N__14387));
    InMux I__1947 (
            .O(N__14407),
            .I(N__14387));
    InMux I__1946 (
            .O(N__14406),
            .I(N__14378));
    InMux I__1945 (
            .O(N__14403),
            .I(N__14378));
    InMux I__1944 (
            .O(N__14402),
            .I(N__14378));
    InMux I__1943 (
            .O(N__14401),
            .I(N__14378));
    Odrv4 I__1942 (
            .O(N__14398),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1941 (
            .O(N__14395),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1940 (
            .O(N__14392),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1939 (
            .O(N__14387),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1938 (
            .O(N__14378),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    CascadeMux I__1937 (
            .O(N__14367),
            .I(\this_vga_signals.N_18_0_cascade_ ));
    InMux I__1936 (
            .O(N__14364),
            .I(N__14360));
    InMux I__1935 (
            .O(N__14363),
            .I(N__14356));
    LocalMux I__1934 (
            .O(N__14360),
            .I(N__14353));
    InMux I__1933 (
            .O(N__14359),
            .I(N__14343));
    LocalMux I__1932 (
            .O(N__14356),
            .I(N__14338));
    Span4Mux_v I__1931 (
            .O(N__14353),
            .I(N__14338));
    InMux I__1930 (
            .O(N__14352),
            .I(N__14335));
    InMux I__1929 (
            .O(N__14351),
            .I(N__14332));
    InMux I__1928 (
            .O(N__14350),
            .I(N__14321));
    InMux I__1927 (
            .O(N__14349),
            .I(N__14321));
    InMux I__1926 (
            .O(N__14348),
            .I(N__14321));
    InMux I__1925 (
            .O(N__14347),
            .I(N__14321));
    InMux I__1924 (
            .O(N__14346),
            .I(N__14321));
    LocalMux I__1923 (
            .O(N__14343),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1922 (
            .O(N__14338),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1921 (
            .O(N__14335),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1920 (
            .O(N__14332),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1919 (
            .O(N__14321),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    CascadeMux I__1918 (
            .O(N__14310),
            .I(N__14306));
    CascadeMux I__1917 (
            .O(N__14309),
            .I(N__14302));
    InMux I__1916 (
            .O(N__14306),
            .I(N__14299));
    InMux I__1915 (
            .O(N__14305),
            .I(N__14296));
    InMux I__1914 (
            .O(N__14302),
            .I(N__14293));
    LocalMux I__1913 (
            .O(N__14299),
            .I(N__14287));
    LocalMux I__1912 (
            .O(N__14296),
            .I(N__14282));
    LocalMux I__1911 (
            .O(N__14293),
            .I(N__14282));
    InMux I__1910 (
            .O(N__14292),
            .I(N__14279));
    CascadeMux I__1909 (
            .O(N__14291),
            .I(N__14275));
    InMux I__1908 (
            .O(N__14290),
            .I(N__14271));
    Sp12to4 I__1907 (
            .O(N__14287),
            .I(N__14264));
    Sp12to4 I__1906 (
            .O(N__14282),
            .I(N__14264));
    LocalMux I__1905 (
            .O(N__14279),
            .I(N__14264));
    InMux I__1904 (
            .O(N__14278),
            .I(N__14261));
    InMux I__1903 (
            .O(N__14275),
            .I(N__14256));
    InMux I__1902 (
            .O(N__14274),
            .I(N__14256));
    LocalMux I__1901 (
            .O(N__14271),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv12 I__1900 (
            .O(N__14264),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1899 (
            .O(N__14261),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1898 (
            .O(N__14256),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    InMux I__1897 (
            .O(N__14247),
            .I(N__14242));
    InMux I__1896 (
            .O(N__14246),
            .I(N__14237));
    InMux I__1895 (
            .O(N__14245),
            .I(N__14237));
    LocalMux I__1894 (
            .O(N__14242),
            .I(N__14230));
    LocalMux I__1893 (
            .O(N__14237),
            .I(N__14230));
    InMux I__1892 (
            .O(N__14236),
            .I(N__14227));
    InMux I__1891 (
            .O(N__14235),
            .I(N__14221));
    Sp12to4 I__1890 (
            .O(N__14230),
            .I(N__14216));
    LocalMux I__1889 (
            .O(N__14227),
            .I(N__14216));
    InMux I__1888 (
            .O(N__14226),
            .I(N__14213));
    InMux I__1887 (
            .O(N__14225),
            .I(N__14208));
    InMux I__1886 (
            .O(N__14224),
            .I(N__14208));
    LocalMux I__1885 (
            .O(N__14221),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv12 I__1884 (
            .O(N__14216),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1883 (
            .O(N__14213),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1882 (
            .O(N__14208),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    CascadeMux I__1881 (
            .O(N__14199),
            .I(\this_vga_signals.m23_1_cascade_ ));
    CascadeMux I__1880 (
            .O(N__14196),
            .I(N__14193));
    InMux I__1879 (
            .O(N__14193),
            .I(N__14188));
    InMux I__1878 (
            .O(N__14192),
            .I(N__14183));
    InMux I__1877 (
            .O(N__14191),
            .I(N__14183));
    LocalMux I__1876 (
            .O(N__14188),
            .I(N__14175));
    LocalMux I__1875 (
            .O(N__14183),
            .I(N__14175));
    InMux I__1874 (
            .O(N__14182),
            .I(N__14172));
    CascadeMux I__1873 (
            .O(N__14181),
            .I(N__14167));
    InMux I__1872 (
            .O(N__14180),
            .I(N__14164));
    Sp12to4 I__1871 (
            .O(N__14175),
            .I(N__14159));
    LocalMux I__1870 (
            .O(N__14172),
            .I(N__14159));
    InMux I__1869 (
            .O(N__14171),
            .I(N__14156));
    InMux I__1868 (
            .O(N__14170),
            .I(N__14151));
    InMux I__1867 (
            .O(N__14167),
            .I(N__14151));
    LocalMux I__1866 (
            .O(N__14164),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv12 I__1865 (
            .O(N__14159),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1864 (
            .O(N__14156),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1863 (
            .O(N__14151),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__1862 (
            .O(N__14142),
            .I(N__14139));
    LocalMux I__1861 (
            .O(N__14139),
            .I(N__14136));
    Span4Mux_v I__1860 (
            .O(N__14136),
            .I(N__14133));
    Odrv4 I__1859 (
            .O(N__14133),
            .I(M_this_data_tmp_qZ0Z_6));
    InMux I__1858 (
            .O(N__14130),
            .I(N__14127));
    LocalMux I__1857 (
            .O(N__14127),
            .I(N__14124));
    Odrv12 I__1856 (
            .O(N__14124),
            .I(\this_ppu.un3_sprites_addr_cry_1_c_RNITOBZ0Z8 ));
    CascadeMux I__1855 (
            .O(N__14121),
            .I(N__14118));
    CascadeBuf I__1854 (
            .O(N__14118),
            .I(N__14115));
    CascadeMux I__1853 (
            .O(N__14115),
            .I(N__14112));
    CascadeBuf I__1852 (
            .O(N__14112),
            .I(N__14109));
    CascadeMux I__1851 (
            .O(N__14109),
            .I(N__14106));
    CascadeBuf I__1850 (
            .O(N__14106),
            .I(N__14103));
    CascadeMux I__1849 (
            .O(N__14103),
            .I(N__14100));
    CascadeBuf I__1848 (
            .O(N__14100),
            .I(N__14097));
    CascadeMux I__1847 (
            .O(N__14097),
            .I(N__14094));
    CascadeBuf I__1846 (
            .O(N__14094),
            .I(N__14091));
    CascadeMux I__1845 (
            .O(N__14091),
            .I(N__14088));
    CascadeBuf I__1844 (
            .O(N__14088),
            .I(N__14085));
    CascadeMux I__1843 (
            .O(N__14085),
            .I(N__14082));
    CascadeBuf I__1842 (
            .O(N__14082),
            .I(N__14079));
    CascadeMux I__1841 (
            .O(N__14079),
            .I(N__14076));
    CascadeBuf I__1840 (
            .O(N__14076),
            .I(N__14073));
    CascadeMux I__1839 (
            .O(N__14073),
            .I(N__14070));
    CascadeBuf I__1838 (
            .O(N__14070),
            .I(N__14067));
    CascadeMux I__1837 (
            .O(N__14067),
            .I(N__14064));
    CascadeBuf I__1836 (
            .O(N__14064),
            .I(N__14061));
    CascadeMux I__1835 (
            .O(N__14061),
            .I(N__14058));
    CascadeBuf I__1834 (
            .O(N__14058),
            .I(N__14055));
    CascadeMux I__1833 (
            .O(N__14055),
            .I(N__14052));
    CascadeBuf I__1832 (
            .O(N__14052),
            .I(N__14049));
    CascadeMux I__1831 (
            .O(N__14049),
            .I(N__14046));
    CascadeBuf I__1830 (
            .O(N__14046),
            .I(N__14043));
    CascadeMux I__1829 (
            .O(N__14043),
            .I(N__14040));
    CascadeBuf I__1828 (
            .O(N__14040),
            .I(N__14037));
    CascadeMux I__1827 (
            .O(N__14037),
            .I(N__14034));
    CascadeBuf I__1826 (
            .O(N__14034),
            .I(N__14031));
    CascadeMux I__1825 (
            .O(N__14031),
            .I(N__14028));
    InMux I__1824 (
            .O(N__14028),
            .I(N__14025));
    LocalMux I__1823 (
            .O(N__14025),
            .I(N__14022));
    Span12Mux_s5_v I__1822 (
            .O(N__14022),
            .I(N__14019));
    Span12Mux_h I__1821 (
            .O(N__14019),
            .I(N__14016));
    Odrv12 I__1820 (
            .O(N__14016),
            .I(M_this_ppu_sprites_addr_2));
    CascadeMux I__1819 (
            .O(N__14013),
            .I(\this_ppu.un1_M_haddress_q_c1_cascade_ ));
    CEMux I__1818 (
            .O(N__14010),
            .I(N__14007));
    LocalMux I__1817 (
            .O(N__14007),
            .I(N__14004));
    Span4Mux_h I__1816 (
            .O(N__14004),
            .I(N__14001));
    Span4Mux_v I__1815 (
            .O(N__14001),
            .I(N__13998));
    Span4Mux_v I__1814 (
            .O(N__13998),
            .I(N__13992));
    InMux I__1813 (
            .O(N__13997),
            .I(N__13987));
    InMux I__1812 (
            .O(N__13996),
            .I(N__13987));
    InMux I__1811 (
            .O(N__13995),
            .I(N__13984));
    Odrv4 I__1810 (
            .O(N__13992),
            .I(M_this_ppu_vram_en_0));
    LocalMux I__1809 (
            .O(N__13987),
            .I(M_this_ppu_vram_en_0));
    LocalMux I__1808 (
            .O(N__13984),
            .I(M_this_ppu_vram_en_0));
    InMux I__1807 (
            .O(N__13977),
            .I(N__13972));
    InMux I__1806 (
            .O(N__13976),
            .I(N__13967));
    InMux I__1805 (
            .O(N__13975),
            .I(N__13967));
    LocalMux I__1804 (
            .O(N__13972),
            .I(\this_ppu.N_134 ));
    LocalMux I__1803 (
            .O(N__13967),
            .I(\this_ppu.N_134 ));
    CascadeMux I__1802 (
            .O(N__13962),
            .I(N__13959));
    CascadeBuf I__1801 (
            .O(N__13959),
            .I(N__13956));
    CascadeMux I__1800 (
            .O(N__13956),
            .I(N__13953));
    InMux I__1799 (
            .O(N__13953),
            .I(N__13949));
    CascadeMux I__1798 (
            .O(N__13952),
            .I(N__13946));
    LocalMux I__1797 (
            .O(N__13949),
            .I(N__13942));
    InMux I__1796 (
            .O(N__13946),
            .I(N__13939));
    CascadeMux I__1795 (
            .O(N__13945),
            .I(N__13936));
    Span4Mux_h I__1794 (
            .O(N__13942),
            .I(N__13933));
    LocalMux I__1793 (
            .O(N__13939),
            .I(N__13930));
    InMux I__1792 (
            .O(N__13936),
            .I(N__13924));
    Span4Mux_h I__1791 (
            .O(N__13933),
            .I(N__13921));
    Sp12to4 I__1790 (
            .O(N__13930),
            .I(N__13918));
    InMux I__1789 (
            .O(N__13929),
            .I(N__13915));
    InMux I__1788 (
            .O(N__13928),
            .I(N__13912));
    InMux I__1787 (
            .O(N__13927),
            .I(N__13909));
    LocalMux I__1786 (
            .O(N__13924),
            .I(N__13906));
    Sp12to4 I__1785 (
            .O(N__13921),
            .I(N__13901));
    Span12Mux_h I__1784 (
            .O(N__13918),
            .I(N__13901));
    LocalMux I__1783 (
            .O(N__13915),
            .I(M_this_ppu_map_addr_0));
    LocalMux I__1782 (
            .O(N__13912),
            .I(M_this_ppu_map_addr_0));
    LocalMux I__1781 (
            .O(N__13909),
            .I(M_this_ppu_map_addr_0));
    Odrv12 I__1780 (
            .O(N__13906),
            .I(M_this_ppu_map_addr_0));
    Odrv12 I__1779 (
            .O(N__13901),
            .I(M_this_ppu_map_addr_0));
    CascadeMux I__1778 (
            .O(N__13890),
            .I(N__13887));
    InMux I__1777 (
            .O(N__13887),
            .I(N__13884));
    LocalMux I__1776 (
            .O(N__13884),
            .I(N__13881));
    Span4Mux_v I__1775 (
            .O(N__13881),
            .I(N__13877));
    CascadeMux I__1774 (
            .O(N__13880),
            .I(N__13874));
    Span4Mux_v I__1773 (
            .O(N__13877),
            .I(N__13870));
    InMux I__1772 (
            .O(N__13874),
            .I(N__13867));
    InMux I__1771 (
            .O(N__13873),
            .I(N__13860));
    Span4Mux_v I__1770 (
            .O(N__13870),
            .I(N__13855));
    LocalMux I__1769 (
            .O(N__13867),
            .I(N__13855));
    InMux I__1768 (
            .O(N__13866),
            .I(N__13850));
    InMux I__1767 (
            .O(N__13865),
            .I(N__13850));
    InMux I__1766 (
            .O(N__13864),
            .I(N__13845));
    InMux I__1765 (
            .O(N__13863),
            .I(N__13845));
    LocalMux I__1764 (
            .O(N__13860),
            .I(N__13840));
    Span4Mux_h I__1763 (
            .O(N__13855),
            .I(N__13840));
    LocalMux I__1762 (
            .O(N__13850),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__1761 (
            .O(N__13845),
            .I(M_this_ppu_vram_addr_2));
    Odrv4 I__1760 (
            .O(N__13840),
            .I(M_this_ppu_vram_addr_2));
    InMux I__1759 (
            .O(N__13833),
            .I(N__13830));
    LocalMux I__1758 (
            .O(N__13830),
            .I(\this_ppu.un1_M_haddress_q_c2 ));
    CascadeMux I__1757 (
            .O(N__13827),
            .I(N__13824));
    CascadeBuf I__1756 (
            .O(N__13824),
            .I(N__13821));
    CascadeMux I__1755 (
            .O(N__13821),
            .I(N__13817));
    CascadeMux I__1754 (
            .O(N__13820),
            .I(N__13814));
    InMux I__1753 (
            .O(N__13817),
            .I(N__13810));
    InMux I__1752 (
            .O(N__13814),
            .I(N__13807));
    CascadeMux I__1751 (
            .O(N__13813),
            .I(N__13804));
    LocalMux I__1750 (
            .O(N__13810),
            .I(N__13801));
    LocalMux I__1749 (
            .O(N__13807),
            .I(N__13798));
    InMux I__1748 (
            .O(N__13804),
            .I(N__13793));
    Span4Mux_v I__1747 (
            .O(N__13801),
            .I(N__13788));
    Span4Mux_v I__1746 (
            .O(N__13798),
            .I(N__13788));
    CascadeMux I__1745 (
            .O(N__13797),
            .I(N__13785));
    InMux I__1744 (
            .O(N__13796),
            .I(N__13782));
    LocalMux I__1743 (
            .O(N__13793),
            .I(N__13779));
    Span4Mux_h I__1742 (
            .O(N__13788),
            .I(N__13776));
    InMux I__1741 (
            .O(N__13785),
            .I(N__13773));
    LocalMux I__1740 (
            .O(N__13782),
            .I(N__13768));
    Span4Mux_h I__1739 (
            .O(N__13779),
            .I(N__13768));
    Span4Mux_v I__1738 (
            .O(N__13776),
            .I(N__13765));
    LocalMux I__1737 (
            .O(N__13773),
            .I(M_this_ppu_map_addr_1));
    Odrv4 I__1736 (
            .O(N__13768),
            .I(M_this_ppu_map_addr_1));
    Odrv4 I__1735 (
            .O(N__13765),
            .I(M_this_ppu_map_addr_1));
    InMux I__1734 (
            .O(N__13758),
            .I(N__13755));
    LocalMux I__1733 (
            .O(N__13755),
            .I(\this_ppu.N_128 ));
    InMux I__1732 (
            .O(N__13752),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__1731 (
            .O(N__13749),
            .I(bfn_12_22_0_));
    InMux I__1730 (
            .O(N__13746),
            .I(N__13742));
    InMux I__1729 (
            .O(N__13745),
            .I(N__13739));
    LocalMux I__1728 (
            .O(N__13742),
            .I(\this_vga_signals.M_pcounter_q_i_3_0 ));
    LocalMux I__1727 (
            .O(N__13739),
            .I(\this_vga_signals.M_pcounter_q_i_3_0 ));
    CascadeMux I__1726 (
            .O(N__13734),
            .I(N__13729));
    InMux I__1725 (
            .O(N__13733),
            .I(N__13725));
    InMux I__1724 (
            .O(N__13732),
            .I(N__13722));
    InMux I__1723 (
            .O(N__13729),
            .I(N__13717));
    InMux I__1722 (
            .O(N__13728),
            .I(N__13717));
    LocalMux I__1721 (
            .O(N__13725),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    LocalMux I__1720 (
            .O(N__13722),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    LocalMux I__1719 (
            .O(N__13717),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    CascadeMux I__1718 (
            .O(N__13710),
            .I(N__13705));
    InMux I__1717 (
            .O(N__13709),
            .I(N__13702));
    InMux I__1716 (
            .O(N__13708),
            .I(N__13697));
    InMux I__1715 (
            .O(N__13705),
            .I(N__13697));
    LocalMux I__1714 (
            .O(N__13702),
            .I(N__13692));
    LocalMux I__1713 (
            .O(N__13697),
            .I(N__13692));
    Odrv4 I__1712 (
            .O(N__13692),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    InMux I__1711 (
            .O(N__13689),
            .I(N__13686));
    LocalMux I__1710 (
            .O(N__13686),
            .I(N__13683));
    Span4Mux_v I__1709 (
            .O(N__13683),
            .I(N__13680));
    Odrv4 I__1708 (
            .O(N__13680),
            .I(N_815_0));
    InMux I__1707 (
            .O(N__13677),
            .I(N__13674));
    LocalMux I__1706 (
            .O(N__13674),
            .I(N__13671));
    Span4Mux_h I__1705 (
            .O(N__13671),
            .I(N__13668));
    Span4Mux_h I__1704 (
            .O(N__13668),
            .I(N__13665));
    Odrv4 I__1703 (
            .O(N__13665),
            .I(N_814_0));
    CascadeMux I__1702 (
            .O(N__13662),
            .I(N__13659));
    CascadeBuf I__1701 (
            .O(N__13659),
            .I(N__13656));
    CascadeMux I__1700 (
            .O(N__13656),
            .I(N__13653));
    InMux I__1699 (
            .O(N__13653),
            .I(N__13650));
    LocalMux I__1698 (
            .O(N__13650),
            .I(N__13647));
    Odrv12 I__1697 (
            .O(N__13647),
            .I(this_ppu_M_vaddress_q_i_6));
    InMux I__1696 (
            .O(N__13644),
            .I(N__13641));
    LocalMux I__1695 (
            .O(N__13641),
            .I(N__13638));
    Odrv12 I__1694 (
            .O(N__13638),
            .I(M_this_data_tmp_qZ0Z_1));
    InMux I__1693 (
            .O(N__13635),
            .I(N__13632));
    LocalMux I__1692 (
            .O(N__13632),
            .I(N__13629));
    Span4Mux_h I__1691 (
            .O(N__13629),
            .I(N__13626));
    Odrv4 I__1690 (
            .O(N__13626),
            .I(M_this_data_tmp_qZ0Z_24));
    CascadeMux I__1689 (
            .O(N__13623),
            .I(N__13620));
    InMux I__1688 (
            .O(N__13620),
            .I(N__13617));
    LocalMux I__1687 (
            .O(N__13617),
            .I(N__13614));
    Span4Mux_h I__1686 (
            .O(N__13614),
            .I(N__13611));
    Span4Mux_v I__1685 (
            .O(N__13611),
            .I(N__13608));
    Span4Mux_v I__1684 (
            .O(N__13608),
            .I(N__13601));
    InMux I__1683 (
            .O(N__13607),
            .I(N__13596));
    InMux I__1682 (
            .O(N__13606),
            .I(N__13596));
    InMux I__1681 (
            .O(N__13605),
            .I(N__13591));
    InMux I__1680 (
            .O(N__13604),
            .I(N__13591));
    Odrv4 I__1679 (
            .O(N__13601),
            .I(M_this_ppu_vram_addr_6));
    LocalMux I__1678 (
            .O(N__13596),
            .I(M_this_ppu_vram_addr_6));
    LocalMux I__1677 (
            .O(N__13591),
            .I(M_this_ppu_vram_addr_6));
    CascadeMux I__1676 (
            .O(N__13584),
            .I(N__13581));
    CascadeBuf I__1675 (
            .O(N__13581),
            .I(N__13578));
    CascadeMux I__1674 (
            .O(N__13578),
            .I(N__13573));
    CascadeMux I__1673 (
            .O(N__13577),
            .I(N__13570));
    CascadeMux I__1672 (
            .O(N__13576),
            .I(N__13567));
    InMux I__1671 (
            .O(N__13573),
            .I(N__13564));
    InMux I__1670 (
            .O(N__13570),
            .I(N__13561));
    InMux I__1669 (
            .O(N__13567),
            .I(N__13555));
    LocalMux I__1668 (
            .O(N__13564),
            .I(N__13550));
    LocalMux I__1667 (
            .O(N__13561),
            .I(N__13550));
    InMux I__1666 (
            .O(N__13560),
            .I(N__13545));
    InMux I__1665 (
            .O(N__13559),
            .I(N__13545));
    InMux I__1664 (
            .O(N__13558),
            .I(N__13542));
    LocalMux I__1663 (
            .O(N__13555),
            .I(N__13537));
    Span12Mux_v I__1662 (
            .O(N__13550),
            .I(N__13537));
    LocalMux I__1661 (
            .O(N__13545),
            .I(M_this_ppu_map_addr_2));
    LocalMux I__1660 (
            .O(N__13542),
            .I(M_this_ppu_map_addr_2));
    Odrv12 I__1659 (
            .O(N__13537),
            .I(M_this_ppu_map_addr_2));
    CascadeMux I__1658 (
            .O(N__13530),
            .I(\this_ppu.un1_M_haddress_q_c5_cascade_ ));
    InMux I__1657 (
            .O(N__13527),
            .I(N__13523));
    InMux I__1656 (
            .O(N__13526),
            .I(N__13520));
    LocalMux I__1655 (
            .O(N__13523),
            .I(\this_ppu.M_haddress_qZ0Z_7 ));
    LocalMux I__1654 (
            .O(N__13520),
            .I(\this_ppu.M_haddress_qZ0Z_7 ));
    InMux I__1653 (
            .O(N__13515),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__1652 (
            .O(N__13512),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__1651 (
            .O(N__13509),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__1650 (
            .O(N__13506),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__1649 (
            .O(N__13503),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__1648 (
            .O(N__13500),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__1647 (
            .O(N__13497),
            .I(N__13494));
    LocalMux I__1646 (
            .O(N__13494),
            .I(N__13491));
    Odrv4 I__1645 (
            .O(N__13491),
            .I(M_this_data_tmp_qZ0Z_13));
    InMux I__1644 (
            .O(N__13488),
            .I(N__13485));
    LocalMux I__1643 (
            .O(N__13485),
            .I(N__13482));
    Odrv4 I__1642 (
            .O(N__13482),
            .I(M_this_data_tmp_qZ0Z_9));
    InMux I__1641 (
            .O(N__13479),
            .I(N__13476));
    LocalMux I__1640 (
            .O(N__13476),
            .I(N__13473));
    Span4Mux_h I__1639 (
            .O(N__13473),
            .I(N__13470));
    Odrv4 I__1638 (
            .O(N__13470),
            .I(M_this_data_tmp_qZ0Z_0));
    CascadeMux I__1637 (
            .O(N__13467),
            .I(M_this_ppu_vram_data_0_cascade_));
    CascadeMux I__1636 (
            .O(N__13464),
            .I(\this_ppu.N_134_cascade_ ));
    CascadeMux I__1635 (
            .O(N__13461),
            .I(\this_ppu.un1_M_haddress_q_c2_cascade_ ));
    InMux I__1634 (
            .O(N__13458),
            .I(N__13452));
    InMux I__1633 (
            .O(N__13457),
            .I(N__13452));
    LocalMux I__1632 (
            .O(N__13452),
            .I(\this_ppu.un1_M_haddress_q_c5 ));
    InMux I__1631 (
            .O(N__13449),
            .I(N__13446));
    LocalMux I__1630 (
            .O(N__13446),
            .I(\this_vga_signals.i5_mux ));
    IoInMux I__1629 (
            .O(N__13443),
            .I(N__13440));
    LocalMux I__1628 (
            .O(N__13440),
            .I(N__13437));
    Span12Mux_s7_v I__1627 (
            .O(N__13437),
            .I(N__13434));
    Odrv12 I__1626 (
            .O(N__13434),
            .I(this_vga_signals_hsync_1_i));
    CascadeMux I__1625 (
            .O(N__13431),
            .I(N__13428));
    CascadeBuf I__1624 (
            .O(N__13428),
            .I(N__13425));
    CascadeMux I__1623 (
            .O(N__13425),
            .I(N__13422));
    InMux I__1622 (
            .O(N__13422),
            .I(N__13419));
    LocalMux I__1621 (
            .O(N__13419),
            .I(N__13416));
    Span4Mux_h I__1620 (
            .O(N__13416),
            .I(N__13413));
    Odrv4 I__1619 (
            .O(N__13413),
            .I(M_this_ppu_map_addr_9));
    InMux I__1618 (
            .O(N__13410),
            .I(N__13407));
    LocalMux I__1617 (
            .O(N__13407),
            .I(N__13404));
    Span4Mux_v I__1616 (
            .O(N__13404),
            .I(N__13401));
    Odrv4 I__1615 (
            .O(N__13401),
            .I(N_63_0));
    InMux I__1614 (
            .O(N__13398),
            .I(N__13395));
    LocalMux I__1613 (
            .O(N__13395),
            .I(N__13391));
    CascadeMux I__1612 (
            .O(N__13394),
            .I(N__13387));
    Span4Mux_v I__1611 (
            .O(N__13391),
            .I(N__13383));
    InMux I__1610 (
            .O(N__13390),
            .I(N__13380));
    InMux I__1609 (
            .O(N__13387),
            .I(N__13375));
    InMux I__1608 (
            .O(N__13386),
            .I(N__13375));
    Odrv4 I__1607 (
            .O(N__13383),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    LocalMux I__1606 (
            .O(N__13380),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    LocalMux I__1605 (
            .O(N__13375),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    InMux I__1604 (
            .O(N__13368),
            .I(N__13365));
    LocalMux I__1603 (
            .O(N__13365),
            .I(N__13359));
    InMux I__1602 (
            .O(N__13364),
            .I(N__13356));
    InMux I__1601 (
            .O(N__13363),
            .I(N__13351));
    InMux I__1600 (
            .O(N__13362),
            .I(N__13351));
    Odrv12 I__1599 (
            .O(N__13359),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3 ));
    LocalMux I__1598 (
            .O(N__13356),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3 ));
    LocalMux I__1597 (
            .O(N__13351),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3 ));
    CascadeMux I__1596 (
            .O(N__13344),
            .I(N__13341));
    InMux I__1595 (
            .O(N__13341),
            .I(N__13338));
    LocalMux I__1594 (
            .O(N__13338),
            .I(N__13335));
    Span4Mux_h I__1593 (
            .O(N__13335),
            .I(N__13332));
    Odrv4 I__1592 (
            .O(N__13332),
            .I(M_this_vga_signals_address_3));
    InMux I__1591 (
            .O(N__13329),
            .I(N__13326));
    LocalMux I__1590 (
            .O(N__13326),
            .I(\this_vga_signals.SUM_3_1 ));
    CascadeMux I__1589 (
            .O(N__13323),
            .I(N__13320));
    InMux I__1588 (
            .O(N__13320),
            .I(N__13317));
    LocalMux I__1587 (
            .O(N__13317),
            .I(N__13314));
    Span4Mux_h I__1586 (
            .O(N__13314),
            .I(N__13311));
    Odrv4 I__1585 (
            .O(N__13311),
            .I(M_this_vga_signals_address_6));
    InMux I__1584 (
            .O(N__13308),
            .I(N__13305));
    LocalMux I__1583 (
            .O(N__13305),
            .I(N__13302));
    Span4Mux_h I__1582 (
            .O(N__13302),
            .I(N__13299));
    Odrv4 I__1581 (
            .O(N__13299),
            .I(M_this_data_tmp_qZ0Z_29));
    InMux I__1580 (
            .O(N__13296),
            .I(N__13293));
    LocalMux I__1579 (
            .O(N__13293),
            .I(N__13290));
    Odrv12 I__1578 (
            .O(N__13290),
            .I(M_this_data_tmp_qZ0Z_5));
    InMux I__1577 (
            .O(N__13287),
            .I(N__13284));
    LocalMux I__1576 (
            .O(N__13284),
            .I(N__13281));
    Odrv4 I__1575 (
            .O(N__13281),
            .I(M_this_data_tmp_qZ0Z_12));
    InMux I__1574 (
            .O(N__13278),
            .I(N__13272));
    InMux I__1573 (
            .O(N__13277),
            .I(N__13265));
    InMux I__1572 (
            .O(N__13276),
            .I(N__13265));
    InMux I__1571 (
            .O(N__13275),
            .I(N__13265));
    LocalMux I__1570 (
            .O(N__13272),
            .I(\this_vga_signals.SUM_3 ));
    LocalMux I__1569 (
            .O(N__13265),
            .I(\this_vga_signals.SUM_3 ));
    InMux I__1568 (
            .O(N__13260),
            .I(N__13256));
    InMux I__1567 (
            .O(N__13259),
            .I(N__13253));
    LocalMux I__1566 (
            .O(N__13256),
            .I(N_3_0));
    LocalMux I__1565 (
            .O(N__13253),
            .I(N_3_0));
    InMux I__1564 (
            .O(N__13248),
            .I(N__13245));
    LocalMux I__1563 (
            .O(N__13245),
            .I(\this_vga_signals.M_pcounter_q_3_0 ));
    InMux I__1562 (
            .O(N__13242),
            .I(N__13236));
    InMux I__1561 (
            .O(N__13241),
            .I(N__13236));
    LocalMux I__1560 (
            .O(N__13236),
            .I(\this_vga_signals.N_17_0 ));
    InMux I__1559 (
            .O(N__13233),
            .I(N__13230));
    LocalMux I__1558 (
            .O(N__13230),
            .I(\this_vga_signals.M_hcounter_q_RNI9JJM1Z0Z_0 ));
    CascadeMux I__1557 (
            .O(N__13227),
            .I(\this_vga_signals.M_hcounter_q_RNIADGD1Z0Z_5_cascade_ ));
    IoInMux I__1556 (
            .O(N__13224),
            .I(N__13221));
    LocalMux I__1555 (
            .O(N__13221),
            .I(N__13218));
    Span4Mux_s1_v I__1554 (
            .O(N__13218),
            .I(N__13215));
    Sp12to4 I__1553 (
            .O(N__13215),
            .I(N__13212));
    Span12Mux_s10_h I__1552 (
            .O(N__13212),
            .I(N__13209));
    Odrv12 I__1551 (
            .O(N__13209),
            .I(this_vga_signals_hvisibility_i));
    CascadeMux I__1550 (
            .O(N__13206),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_2_cascade_ ));
    InMux I__1549 (
            .O(N__13203),
            .I(N__13200));
    LocalMux I__1548 (
            .O(N__13200),
            .I(\this_vga_signals.mult1_un89_sum_c3_0 ));
    CascadeMux I__1547 (
            .O(N__13197),
            .I(N__13194));
    InMux I__1546 (
            .O(N__13194),
            .I(N__13191));
    LocalMux I__1545 (
            .O(N__13191),
            .I(N__13188));
    Span4Mux_v I__1544 (
            .O(N__13188),
            .I(N__13185));
    Span4Mux_v I__1543 (
            .O(N__13185),
            .I(N__13182));
    Odrv4 I__1542 (
            .O(N__13182),
            .I(M_this_vga_signals_address_0));
    InMux I__1541 (
            .O(N__13179),
            .I(N__13176));
    LocalMux I__1540 (
            .O(N__13176),
            .I(N__13173));
    Span4Mux_v I__1539 (
            .O(N__13173),
            .I(N__13169));
    CascadeMux I__1538 (
            .O(N__13172),
            .I(N__13166));
    Span4Mux_v I__1537 (
            .O(N__13169),
            .I(N__13162));
    InMux I__1536 (
            .O(N__13166),
            .I(N__13157));
    InMux I__1535 (
            .O(N__13165),
            .I(N__13157));
    Odrv4 I__1534 (
            .O(N__13162),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__1533 (
            .O(N__13157),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    InMux I__1532 (
            .O(N__13152),
            .I(N__13149));
    LocalMux I__1531 (
            .O(N__13149),
            .I(\this_vga_signals.mult1_un82_sum_axb1 ));
    InMux I__1530 (
            .O(N__13146),
            .I(N__13143));
    LocalMux I__1529 (
            .O(N__13143),
            .I(N__13139));
    InMux I__1528 (
            .O(N__13142),
            .I(N__13136));
    Odrv4 I__1527 (
            .O(N__13139),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_1 ));
    LocalMux I__1526 (
            .O(N__13136),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_1 ));
    InMux I__1525 (
            .O(N__13131),
            .I(N__13128));
    LocalMux I__1524 (
            .O(N__13128),
            .I(N__13125));
    Span4Mux_v I__1523 (
            .O(N__13125),
            .I(N__13121));
    InMux I__1522 (
            .O(N__13124),
            .I(N__13118));
    Odrv4 I__1521 (
            .O(N__13121),
            .I(\this_vga_signals.mult1_un82_sum_c3 ));
    LocalMux I__1520 (
            .O(N__13118),
            .I(\this_vga_signals.mult1_un82_sum_c3 ));
    InMux I__1519 (
            .O(N__13113),
            .I(N__13107));
    InMux I__1518 (
            .O(N__13112),
            .I(N__13107));
    LocalMux I__1517 (
            .O(N__13107),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3 ));
    InMux I__1516 (
            .O(N__13104),
            .I(N__13101));
    LocalMux I__1515 (
            .O(N__13101),
            .I(N__13098));
    Span4Mux_h I__1514 (
            .O(N__13098),
            .I(N__13095));
    Span4Mux_v I__1513 (
            .O(N__13095),
            .I(N__13091));
    InMux I__1512 (
            .O(N__13094),
            .I(N__13088));
    Odrv4 I__1511 (
            .O(N__13091),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__1510 (
            .O(N__13088),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    InMux I__1509 (
            .O(N__13083),
            .I(N__13077));
    InMux I__1508 (
            .O(N__13082),
            .I(N__13077));
    LocalMux I__1507 (
            .O(N__13077),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    CascadeMux I__1506 (
            .O(N__13074),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_ ));
    CascadeMux I__1505 (
            .O(N__13071),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_ ));
    CascadeMux I__1504 (
            .O(N__13068),
            .I(N__13065));
    InMux I__1503 (
            .O(N__13065),
            .I(N__13056));
    InMux I__1502 (
            .O(N__13064),
            .I(N__13056));
    InMux I__1501 (
            .O(N__13063),
            .I(N__13056));
    LocalMux I__1500 (
            .O(N__13056),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9 ));
    InMux I__1499 (
            .O(N__13053),
            .I(N__13050));
    LocalMux I__1498 (
            .O(N__13050),
            .I(N__13046));
    InMux I__1497 (
            .O(N__13049),
            .I(N__13043));
    Span12Mux_s10_v I__1496 (
            .O(N__13046),
            .I(N__13035));
    LocalMux I__1495 (
            .O(N__13043),
            .I(N__13032));
    InMux I__1494 (
            .O(N__13042),
            .I(N__13023));
    InMux I__1493 (
            .O(N__13041),
            .I(N__13023));
    InMux I__1492 (
            .O(N__13040),
            .I(N__13023));
    InMux I__1491 (
            .O(N__13039),
            .I(N__13023));
    InMux I__1490 (
            .O(N__13038),
            .I(N__13020));
    Odrv12 I__1489 (
            .O(N__13035),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    Odrv4 I__1488 (
            .O(N__13032),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1487 (
            .O(N__13023),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1486 (
            .O(N__13020),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    CascadeMux I__1485 (
            .O(N__13011),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_cascade_ ));
    InMux I__1484 (
            .O(N__13008),
            .I(N__13005));
    LocalMux I__1483 (
            .O(N__13005),
            .I(\this_vga_signals.mult1_un68_sum_axb1 ));
    CascadeMux I__1482 (
            .O(N__13002),
            .I(\this_vga_signals.if_i4_mux_0_cascade_ ));
    InMux I__1481 (
            .O(N__12999),
            .I(N__12994));
    InMux I__1480 (
            .O(N__12998),
            .I(N__12991));
    InMux I__1479 (
            .O(N__12997),
            .I(N__12988));
    LocalMux I__1478 (
            .O(N__12994),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    LocalMux I__1477 (
            .O(N__12991),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    LocalMux I__1476 (
            .O(N__12988),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    InMux I__1475 (
            .O(N__12981),
            .I(N__12978));
    LocalMux I__1474 (
            .O(N__12978),
            .I(\this_vga_signals.M_hcounter_q_RNIUULS4Z0Z_3 ));
    InMux I__1473 (
            .O(N__12975),
            .I(N__12971));
    InMux I__1472 (
            .O(N__12974),
            .I(N__12968));
    LocalMux I__1471 (
            .O(N__12971),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    LocalMux I__1470 (
            .O(N__12968),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    CascadeMux I__1469 (
            .O(N__12963),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ));
    CascadeMux I__1468 (
            .O(N__12960),
            .I(N__12957));
    InMux I__1467 (
            .O(N__12957),
            .I(N__12954));
    LocalMux I__1466 (
            .O(N__12954),
            .I(\this_vga_signals.if_m2_2 ));
    CascadeMux I__1465 (
            .O(N__12951),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_1_cascade_ ));
    InMux I__1464 (
            .O(N__12948),
            .I(N__12944));
    InMux I__1463 (
            .O(N__12947),
            .I(N__12941));
    LocalMux I__1462 (
            .O(N__12944),
            .I(\this_vga_signals.d_N_3_0_i ));
    LocalMux I__1461 (
            .O(N__12941),
            .I(\this_vga_signals.d_N_3_0_i ));
    InMux I__1460 (
            .O(N__12936),
            .I(N__12933));
    LocalMux I__1459 (
            .O(N__12933),
            .I(\this_vga_signals.mult1_un82_sum_c2_0 ));
    InMux I__1458 (
            .O(N__12930),
            .I(N__12927));
    LocalMux I__1457 (
            .O(N__12927),
            .I(N__12924));
    Odrv4 I__1456 (
            .O(N__12924),
            .I(M_this_data_tmp_qZ0Z_28));
    InMux I__1455 (
            .O(N__12921),
            .I(N__12918));
    LocalMux I__1454 (
            .O(N__12918),
            .I(N__12915));
    Span4Mux_h I__1453 (
            .O(N__12915),
            .I(N__12912));
    Odrv4 I__1452 (
            .O(N__12912),
            .I(N_833_0));
    InMux I__1451 (
            .O(N__12909),
            .I(N__12906));
    LocalMux I__1450 (
            .O(N__12906),
            .I(N__12903));
    Span4Mux_h I__1449 (
            .O(N__12903),
            .I(N__12899));
    InMux I__1448 (
            .O(N__12902),
            .I(N__12896));
    Odrv4 I__1447 (
            .O(N__12899),
            .I(M_this_oam_ram_read_data_16));
    LocalMux I__1446 (
            .O(N__12896),
            .I(M_this_oam_ram_read_data_16));
    CascadeMux I__1445 (
            .O(N__12891),
            .I(N__12888));
    CascadeBuf I__1444 (
            .O(N__12888),
            .I(N__12885));
    CascadeMux I__1443 (
            .O(N__12885),
            .I(N__12882));
    InMux I__1442 (
            .O(N__12882),
            .I(N__12879));
    LocalMux I__1441 (
            .O(N__12879),
            .I(N__12875));
    InMux I__1440 (
            .O(N__12878),
            .I(N__12872));
    Span4Mux_v I__1439 (
            .O(N__12875),
            .I(N__12869));
    LocalMux I__1438 (
            .O(N__12872),
            .I(N__12864));
    Span4Mux_v I__1437 (
            .O(N__12869),
            .I(N__12864));
    Odrv4 I__1436 (
            .O(N__12864),
            .I(M_this_ppu_vram_addr_i_6));
    InMux I__1435 (
            .O(N__12861),
            .I(N__12858));
    LocalMux I__1434 (
            .O(N__12858),
            .I(M_this_data_tmp_qZ0Z_18));
    InMux I__1433 (
            .O(N__12855),
            .I(N__12852));
    LocalMux I__1432 (
            .O(N__12852),
            .I(N__12849));
    Span4Mux_v I__1431 (
            .O(N__12849),
            .I(N__12846));
    Span4Mux_h I__1430 (
            .O(N__12846),
            .I(N__12843));
    Odrv4 I__1429 (
            .O(N__12843),
            .I(M_this_oam_ram_write_data_18));
    CascadeMux I__1428 (
            .O(N__12840),
            .I(N__12837));
    CascadeBuf I__1427 (
            .O(N__12837),
            .I(N__12834));
    CascadeMux I__1426 (
            .O(N__12834),
            .I(N__12831));
    InMux I__1425 (
            .O(N__12831),
            .I(N__12828));
    LocalMux I__1424 (
            .O(N__12828),
            .I(N__12824));
    InMux I__1423 (
            .O(N__12827),
            .I(N__12821));
    Span4Mux_v I__1422 (
            .O(N__12824),
            .I(N__12818));
    LocalMux I__1421 (
            .O(N__12821),
            .I(N__12813));
    Span4Mux_v I__1420 (
            .O(N__12818),
            .I(N__12813));
    Odrv4 I__1419 (
            .O(N__12813),
            .I(M_this_ppu_map_addr_4));
    InMux I__1418 (
            .O(N__12810),
            .I(N__12807));
    LocalMux I__1417 (
            .O(N__12807),
            .I(N__12804));
    Odrv4 I__1416 (
            .O(N__12804),
            .I(M_this_data_tmp_qZ0Z_30));
    InMux I__1415 (
            .O(N__12801),
            .I(N__12798));
    LocalMux I__1414 (
            .O(N__12798),
            .I(N__12795));
    Odrv4 I__1413 (
            .O(N__12795),
            .I(N_830_0));
    InMux I__1412 (
            .O(N__12792),
            .I(N__12789));
    LocalMux I__1411 (
            .O(N__12789),
            .I(M_this_data_tmp_qZ0Z_16));
    InMux I__1410 (
            .O(N__12786),
            .I(N__12783));
    LocalMux I__1409 (
            .O(N__12783),
            .I(N__12780));
    Span4Mux_h I__1408 (
            .O(N__12780),
            .I(N__12777));
    Odrv4 I__1407 (
            .O(N__12777),
            .I(M_this_oam_ram_write_data_16));
    InMux I__1406 (
            .O(N__12774),
            .I(N__12771));
    LocalMux I__1405 (
            .O(N__12771),
            .I(N__12768));
    Odrv4 I__1404 (
            .O(N__12768),
            .I(M_this_data_tmp_qZ0Z_14));
    InMux I__1403 (
            .O(N__12765),
            .I(N__12762));
    LocalMux I__1402 (
            .O(N__12762),
            .I(N__12759));
    Span4Mux_h I__1401 (
            .O(N__12759),
            .I(N__12756));
    Odrv4 I__1400 (
            .O(N__12756),
            .I(M_this_data_tmp_qZ0Z_27));
    InMux I__1399 (
            .O(N__12753),
            .I(N__12750));
    LocalMux I__1398 (
            .O(N__12750),
            .I(M_this_data_tmp_qZ0Z_3));
    InMux I__1397 (
            .O(N__12747),
            .I(N__12744));
    LocalMux I__1396 (
            .O(N__12744),
            .I(N__12741));
    Odrv12 I__1395 (
            .O(N__12741),
            .I(M_this_data_tmp_qZ0Z_7));
    InMux I__1394 (
            .O(N__12738),
            .I(N__12735));
    LocalMux I__1393 (
            .O(N__12735),
            .I(M_this_data_tmp_qZ0Z_2));
    InMux I__1392 (
            .O(N__12732),
            .I(N__12729));
    LocalMux I__1391 (
            .O(N__12729),
            .I(N__12726));
    Odrv4 I__1390 (
            .O(N__12726),
            .I(M_this_data_tmp_qZ0Z_4));
    InMux I__1389 (
            .O(N__12723),
            .I(N__12720));
    LocalMux I__1388 (
            .O(N__12720),
            .I(M_this_data_tmp_qZ0Z_25));
    InMux I__1387 (
            .O(N__12717),
            .I(N__12714));
    LocalMux I__1386 (
            .O(N__12714),
            .I(N__12711));
    Odrv4 I__1385 (
            .O(N__12711),
            .I(M_this_data_tmp_qZ0Z_31));
    InMux I__1384 (
            .O(N__12708),
            .I(N__12705));
    LocalMux I__1383 (
            .O(N__12705),
            .I(M_this_vga_signals_pixel_clk_0_0));
    CascadeMux I__1382 (
            .O(N__12702),
            .I(\this_vga_ramdac.i2_mux_0_cascade_ ));
    InMux I__1381 (
            .O(N__12699),
            .I(N__12696));
    LocalMux I__1380 (
            .O(N__12696),
            .I(N__12692));
    InMux I__1379 (
            .O(N__12695),
            .I(N__12689));
    Odrv4 I__1378 (
            .O(N__12692),
            .I(\this_vga_ramdac.N_2615_reto ));
    LocalMux I__1377 (
            .O(N__12689),
            .I(\this_vga_ramdac.N_2615_reto ));
    CascadeMux I__1376 (
            .O(N__12684),
            .I(\this_vga_ramdac.m16_cascade_ ));
    InMux I__1375 (
            .O(N__12681),
            .I(N__12676));
    InMux I__1374 (
            .O(N__12680),
            .I(N__12671));
    InMux I__1373 (
            .O(N__12679),
            .I(N__12671));
    LocalMux I__1372 (
            .O(N__12676),
            .I(N__12663));
    LocalMux I__1371 (
            .O(N__12671),
            .I(N__12663));
    InMux I__1370 (
            .O(N__12670),
            .I(N__12660));
    InMux I__1369 (
            .O(N__12669),
            .I(N__12655));
    InMux I__1368 (
            .O(N__12668),
            .I(N__12655));
    Odrv4 I__1367 (
            .O(N__12663),
            .I(G_480));
    LocalMux I__1366 (
            .O(N__12660),
            .I(G_480));
    LocalMux I__1365 (
            .O(N__12655),
            .I(G_480));
    InMux I__1364 (
            .O(N__12648),
            .I(N__12645));
    LocalMux I__1363 (
            .O(N__12645),
            .I(N__12641));
    InMux I__1362 (
            .O(N__12644),
            .I(N__12638));
    Odrv4 I__1361 (
            .O(N__12641),
            .I(\this_vga_ramdac.N_2613_reto ));
    LocalMux I__1360 (
            .O(N__12638),
            .I(\this_vga_ramdac.N_2613_reto ));
    InMux I__1359 (
            .O(N__12633),
            .I(N__12630));
    LocalMux I__1358 (
            .O(N__12630),
            .I(N__12627));
    Span4Mux_h I__1357 (
            .O(N__12627),
            .I(N__12624));
    Odrv4 I__1356 (
            .O(N__12624),
            .I(N_73_0));
    InMux I__1355 (
            .O(N__12621),
            .I(N__12618));
    LocalMux I__1354 (
            .O(N__12618),
            .I(N__12615));
    Odrv4 I__1353 (
            .O(N__12615),
            .I(\this_vga_ramdac.N_24_mux ));
    InMux I__1352 (
            .O(N__12612),
            .I(N__12609));
    LocalMux I__1351 (
            .O(N__12609),
            .I(N__12606));
    Odrv4 I__1350 (
            .O(N__12606),
            .I(\this_vga_ramdac.m19 ));
    InMux I__1349 (
            .O(N__12603),
            .I(N__12594));
    InMux I__1348 (
            .O(N__12602),
            .I(N__12594));
    InMux I__1347 (
            .O(N__12601),
            .I(N__12594));
    LocalMux I__1346 (
            .O(N__12594),
            .I(N__12589));
    InMux I__1345 (
            .O(N__12593),
            .I(N__12584));
    InMux I__1344 (
            .O(N__12592),
            .I(N__12584));
    Span4Mux_v I__1343 (
            .O(N__12589),
            .I(N__12578));
    LocalMux I__1342 (
            .O(N__12584),
            .I(N__12578));
    InMux I__1341 (
            .O(N__12583),
            .I(N__12575));
    Span4Mux_h I__1340 (
            .O(N__12578),
            .I(N__12572));
    LocalMux I__1339 (
            .O(N__12575),
            .I(N__12569));
    Span4Mux_v I__1338 (
            .O(N__12572),
            .I(N__12566));
    Span4Mux_v I__1337 (
            .O(N__12569),
            .I(N__12563));
    Odrv4 I__1336 (
            .O(N__12566),
            .I(M_this_vram_read_data_0));
    Odrv4 I__1335 (
            .O(N__12563),
            .I(M_this_vram_read_data_0));
    CascadeMux I__1334 (
            .O(N__12558),
            .I(N__12553));
    CascadeMux I__1333 (
            .O(N__12557),
            .I(N__12547));
    CascadeMux I__1332 (
            .O(N__12556),
            .I(N__12544));
    InMux I__1331 (
            .O(N__12553),
            .I(N__12537));
    InMux I__1330 (
            .O(N__12552),
            .I(N__12537));
    InMux I__1329 (
            .O(N__12551),
            .I(N__12537));
    InMux I__1328 (
            .O(N__12550),
            .I(N__12532));
    InMux I__1327 (
            .O(N__12547),
            .I(N__12532));
    InMux I__1326 (
            .O(N__12544),
            .I(N__12529));
    LocalMux I__1325 (
            .O(N__12537),
            .I(N__12526));
    LocalMux I__1324 (
            .O(N__12532),
            .I(N__12521));
    LocalMux I__1323 (
            .O(N__12529),
            .I(N__12521));
    Span4Mux_h I__1322 (
            .O(N__12526),
            .I(N__12518));
    Span4Mux_h I__1321 (
            .O(N__12521),
            .I(N__12515));
    Span4Mux_v I__1320 (
            .O(N__12518),
            .I(N__12512));
    Odrv4 I__1319 (
            .O(N__12515),
            .I(M_this_vram_read_data_3));
    Odrv4 I__1318 (
            .O(N__12512),
            .I(M_this_vram_read_data_3));
    CascadeMux I__1317 (
            .O(N__12507),
            .I(N__12502));
    CascadeMux I__1316 (
            .O(N__12506),
            .I(N__12498));
    InMux I__1315 (
            .O(N__12505),
            .I(N__12489));
    InMux I__1314 (
            .O(N__12502),
            .I(N__12489));
    InMux I__1313 (
            .O(N__12501),
            .I(N__12489));
    InMux I__1312 (
            .O(N__12498),
            .I(N__12484));
    InMux I__1311 (
            .O(N__12497),
            .I(N__12484));
    InMux I__1310 (
            .O(N__12496),
            .I(N__12481));
    LocalMux I__1309 (
            .O(N__12489),
            .I(N__12476));
    LocalMux I__1308 (
            .O(N__12484),
            .I(N__12476));
    LocalMux I__1307 (
            .O(N__12481),
            .I(N__12473));
    Span12Mux_v I__1306 (
            .O(N__12476),
            .I(N__12470));
    Span4Mux_v I__1305 (
            .O(N__12473),
            .I(N__12467));
    Odrv12 I__1304 (
            .O(N__12470),
            .I(M_this_vram_read_data_1));
    Odrv4 I__1303 (
            .O(N__12467),
            .I(M_this_vram_read_data_1));
    InMux I__1302 (
            .O(N__12462),
            .I(N__12456));
    InMux I__1301 (
            .O(N__12461),
            .I(N__12456));
    LocalMux I__1300 (
            .O(N__12456),
            .I(N__12450));
    InMux I__1299 (
            .O(N__12455),
            .I(N__12445));
    InMux I__1298 (
            .O(N__12454),
            .I(N__12445));
    InMux I__1297 (
            .O(N__12453),
            .I(N__12442));
    Span4Mux_h I__1296 (
            .O(N__12450),
            .I(N__12439));
    LocalMux I__1295 (
            .O(N__12445),
            .I(N__12434));
    LocalMux I__1294 (
            .O(N__12442),
            .I(N__12434));
    Span4Mux_v I__1293 (
            .O(N__12439),
            .I(N__12431));
    Span4Mux_h I__1292 (
            .O(N__12434),
            .I(N__12428));
    Odrv4 I__1291 (
            .O(N__12431),
            .I(M_this_vram_read_data_2));
    Odrv4 I__1290 (
            .O(N__12428),
            .I(M_this_vram_read_data_2));
    InMux I__1289 (
            .O(N__12423),
            .I(N__12420));
    LocalMux I__1288 (
            .O(N__12420),
            .I(N__12417));
    Odrv4 I__1287 (
            .O(N__12417),
            .I(\this_vga_ramdac.m6 ));
    CascadeMux I__1286 (
            .O(N__12414),
            .I(\this_vga_signals.mult1_un68_sum_axb1_cascade_ ));
    InMux I__1285 (
            .O(N__12411),
            .I(N__12408));
    LocalMux I__1284 (
            .O(N__12408),
            .I(\this_vga_signals.if_m2_0 ));
    InMux I__1283 (
            .O(N__12405),
            .I(N__12402));
    LocalMux I__1282 (
            .O(N__12402),
            .I(N__12399));
    Span4Mux_h I__1281 (
            .O(N__12399),
            .I(N__12396));
    Span4Mux_v I__1280 (
            .O(N__12396),
            .I(N__12393));
    Odrv4 I__1279 (
            .O(N__12393),
            .I(N_58_0));
    CascadeMux I__1278 (
            .O(N__12390),
            .I(N_3_0_cascade_));
    CascadeMux I__1277 (
            .O(N__12387),
            .I(G_480_cascade_));
    InMux I__1276 (
            .O(N__12384),
            .I(N__12381));
    LocalMux I__1275 (
            .O(N__12381),
            .I(N__12377));
    InMux I__1274 (
            .O(N__12380),
            .I(N__12374));
    Span4Mux_v I__1273 (
            .O(N__12377),
            .I(N__12371));
    LocalMux I__1272 (
            .O(N__12374),
            .I(N__12368));
    Odrv4 I__1271 (
            .O(N__12371),
            .I(\this_vga_ramdac.N_2614_reto ));
    Odrv4 I__1270 (
            .O(N__12368),
            .I(\this_vga_ramdac.N_2614_reto ));
    InMux I__1269 (
            .O(N__12363),
            .I(N__12359));
    InMux I__1268 (
            .O(N__12362),
            .I(N__12356));
    LocalMux I__1267 (
            .O(N__12359),
            .I(\this_vga_ramdac.N_2611_reto ));
    LocalMux I__1266 (
            .O(N__12356),
            .I(\this_vga_ramdac.N_2611_reto ));
    InMux I__1265 (
            .O(N__12351),
            .I(N__12348));
    LocalMux I__1264 (
            .O(N__12348),
            .I(N__12344));
    CascadeMux I__1263 (
            .O(N__12347),
            .I(N__12341));
    Span4Mux_h I__1262 (
            .O(N__12344),
            .I(N__12338));
    InMux I__1261 (
            .O(N__12341),
            .I(N__12335));
    Odrv4 I__1260 (
            .O(N__12338),
            .I(\this_vga_ramdac.N_2610_reto ));
    LocalMux I__1259 (
            .O(N__12335),
            .I(\this_vga_ramdac.N_2610_reto ));
    InMux I__1258 (
            .O(N__12330),
            .I(N__12327));
    LocalMux I__1257 (
            .O(N__12327),
            .I(N_2_0));
    CascadeMux I__1256 (
            .O(N__12324),
            .I(N_2_0_cascade_));
    InMux I__1255 (
            .O(N__12321),
            .I(N__12318));
    LocalMux I__1254 (
            .O(N__12318),
            .I(N__12315));
    Odrv4 I__1253 (
            .O(N__12315),
            .I(M_this_data_tmp_qZ0Z_20));
    InMux I__1252 (
            .O(N__12312),
            .I(N__12309));
    LocalMux I__1251 (
            .O(N__12309),
            .I(M_this_data_tmp_qZ0Z_21));
    InMux I__1250 (
            .O(N__12306),
            .I(N__12303));
    LocalMux I__1249 (
            .O(N__12303),
            .I(M_this_data_tmp_qZ0Z_22));
    InMux I__1248 (
            .O(N__12300),
            .I(N__12297));
    LocalMux I__1247 (
            .O(N__12297),
            .I(N__12294));
    Span4Mux_h I__1246 (
            .O(N__12294),
            .I(N__12291));
    Odrv4 I__1245 (
            .O(N__12291),
            .I(M_this_data_tmp_qZ0Z_23));
    InMux I__1244 (
            .O(N__12288),
            .I(N__12285));
    LocalMux I__1243 (
            .O(N__12285),
            .I(N__12282));
    Odrv4 I__1242 (
            .O(N__12282),
            .I(\this_oam_ram.M_this_oam_ram_read_data_22 ));
    CascadeMux I__1241 (
            .O(N__12279),
            .I(N__12276));
    InMux I__1240 (
            .O(N__12276),
            .I(N__12273));
    LocalMux I__1239 (
            .O(N__12273),
            .I(M_this_oam_ram_read_data_i_22));
    InMux I__1238 (
            .O(N__12270),
            .I(N__12267));
    LocalMux I__1237 (
            .O(N__12267),
            .I(N__12264));
    Span4Mux_h I__1236 (
            .O(N__12264),
            .I(N__12261));
    Odrv4 I__1235 (
            .O(N__12261),
            .I(N_890_0));
    InMux I__1234 (
            .O(N__12258),
            .I(N__12255));
    LocalMux I__1233 (
            .O(N__12255),
            .I(N__12252));
    Odrv4 I__1232 (
            .O(N__12252),
            .I(M_this_oam_ram_write_data_12));
    InMux I__1231 (
            .O(N__12249),
            .I(N__12246));
    LocalMux I__1230 (
            .O(N__12246),
            .I(N__12243));
    Span4Mux_h I__1229 (
            .O(N__12243),
            .I(N__12240));
    Odrv4 I__1228 (
            .O(N__12240),
            .I(N_831_0));
    InMux I__1227 (
            .O(N__12237),
            .I(N__12234));
    LocalMux I__1226 (
            .O(N__12234),
            .I(N__12231));
    Span4Mux_h I__1225 (
            .O(N__12231),
            .I(N__12228));
    Odrv4 I__1224 (
            .O(N__12228),
            .I(M_this_oam_ram_write_data_24));
    InMux I__1223 (
            .O(N__12225),
            .I(N__12222));
    LocalMux I__1222 (
            .O(N__12222),
            .I(N__12219));
    Span4Mux_h I__1221 (
            .O(N__12219),
            .I(N__12216));
    Odrv4 I__1220 (
            .O(N__12216),
            .I(N_832_0));
    InMux I__1219 (
            .O(N__12213),
            .I(N__12210));
    LocalMux I__1218 (
            .O(N__12210),
            .I(N__12207));
    Span4Mux_h I__1217 (
            .O(N__12207),
            .I(N__12204));
    Odrv4 I__1216 (
            .O(N__12204),
            .I(N_893_0));
    InMux I__1215 (
            .O(N__12201),
            .I(N__12198));
    LocalMux I__1214 (
            .O(N__12198),
            .I(M_this_data_tmp_qZ0Z_19));
    CascadeMux I__1213 (
            .O(N__12195),
            .I(N__12192));
    InMux I__1212 (
            .O(N__12192),
            .I(N__12189));
    LocalMux I__1211 (
            .O(N__12189),
            .I(M_this_vga_signals_address_4));
    InMux I__1210 (
            .O(N__12186),
            .I(N__12183));
    LocalMux I__1209 (
            .O(N__12183),
            .I(N__12180));
    Span4Mux_s3_v I__1208 (
            .O(N__12180),
            .I(N__12177));
    Odrv4 I__1207 (
            .O(N__12177),
            .I(M_this_map_ram_read_data_1));
    InMux I__1206 (
            .O(N__12174),
            .I(N__12171));
    LocalMux I__1205 (
            .O(N__12171),
            .I(N__12168));
    Span12Mux_s6_v I__1204 (
            .O(N__12168),
            .I(N__12165));
    Odrv12 I__1203 (
            .O(N__12165),
            .I(\this_ppu.un3_sprites_addr_cry_6_c_RNIP5LZ0Z8 ));
    CascadeMux I__1202 (
            .O(N__12162),
            .I(N__12159));
    CascadeBuf I__1201 (
            .O(N__12159),
            .I(N__12156));
    CascadeMux I__1200 (
            .O(N__12156),
            .I(N__12153));
    CascadeBuf I__1199 (
            .O(N__12153),
            .I(N__12150));
    CascadeMux I__1198 (
            .O(N__12150),
            .I(N__12147));
    CascadeBuf I__1197 (
            .O(N__12147),
            .I(N__12144));
    CascadeMux I__1196 (
            .O(N__12144),
            .I(N__12141));
    CascadeBuf I__1195 (
            .O(N__12141),
            .I(N__12138));
    CascadeMux I__1194 (
            .O(N__12138),
            .I(N__12135));
    CascadeBuf I__1193 (
            .O(N__12135),
            .I(N__12132));
    CascadeMux I__1192 (
            .O(N__12132),
            .I(N__12129));
    CascadeBuf I__1191 (
            .O(N__12129),
            .I(N__12126));
    CascadeMux I__1190 (
            .O(N__12126),
            .I(N__12123));
    CascadeBuf I__1189 (
            .O(N__12123),
            .I(N__12120));
    CascadeMux I__1188 (
            .O(N__12120),
            .I(N__12117));
    CascadeBuf I__1187 (
            .O(N__12117),
            .I(N__12114));
    CascadeMux I__1186 (
            .O(N__12114),
            .I(N__12111));
    CascadeBuf I__1185 (
            .O(N__12111),
            .I(N__12108));
    CascadeMux I__1184 (
            .O(N__12108),
            .I(N__12105));
    CascadeBuf I__1183 (
            .O(N__12105),
            .I(N__12102));
    CascadeMux I__1182 (
            .O(N__12102),
            .I(N__12099));
    CascadeBuf I__1181 (
            .O(N__12099),
            .I(N__12096));
    CascadeMux I__1180 (
            .O(N__12096),
            .I(N__12093));
    CascadeBuf I__1179 (
            .O(N__12093),
            .I(N__12090));
    CascadeMux I__1178 (
            .O(N__12090),
            .I(N__12087));
    CascadeBuf I__1177 (
            .O(N__12087),
            .I(N__12084));
    CascadeMux I__1176 (
            .O(N__12084),
            .I(N__12081));
    CascadeBuf I__1175 (
            .O(N__12081),
            .I(N__12078));
    CascadeMux I__1174 (
            .O(N__12078),
            .I(N__12075));
    CascadeBuf I__1173 (
            .O(N__12075),
            .I(N__12072));
    CascadeMux I__1172 (
            .O(N__12072),
            .I(N__12069));
    InMux I__1171 (
            .O(N__12069),
            .I(N__12066));
    LocalMux I__1170 (
            .O(N__12066),
            .I(N__12063));
    Span12Mux_h I__1169 (
            .O(N__12063),
            .I(N__12060));
    Odrv12 I__1168 (
            .O(N__12060),
            .I(M_this_ppu_sprites_addr_7));
    InMux I__1167 (
            .O(N__12057),
            .I(N__12054));
    LocalMux I__1166 (
            .O(N__12054),
            .I(M_this_data_tmp_qZ0Z_15));
    InMux I__1165 (
            .O(N__12051),
            .I(N__12048));
    LocalMux I__1164 (
            .O(N__12048),
            .I(M_this_data_tmp_qZ0Z_8));
    InMux I__1163 (
            .O(N__12045),
            .I(N__12042));
    LocalMux I__1162 (
            .O(N__12042),
            .I(M_this_data_tmp_qZ0Z_11));
    InMux I__1161 (
            .O(N__12039),
            .I(N__12036));
    LocalMux I__1160 (
            .O(N__12036),
            .I(N__12033));
    Odrv4 I__1159 (
            .O(N__12033),
            .I(N_835_0));
    InMux I__1158 (
            .O(N__12030),
            .I(N__12027));
    LocalMux I__1157 (
            .O(N__12027),
            .I(N__12024));
    Span4Mux_h I__1156 (
            .O(N__12024),
            .I(N__12021));
    Odrv4 I__1155 (
            .O(N__12021),
            .I(N_897_0));
    InMux I__1154 (
            .O(N__12018),
            .I(N__12015));
    LocalMux I__1153 (
            .O(N__12015),
            .I(N__12012));
    Span4Mux_h I__1152 (
            .O(N__12012),
            .I(N__12009));
    Odrv4 I__1151 (
            .O(N__12009),
            .I(N_53_0));
    InMux I__1150 (
            .O(N__12006),
            .I(N__12003));
    LocalMux I__1149 (
            .O(N__12003),
            .I(N__12000));
    Span4Mux_v I__1148 (
            .O(N__12000),
            .I(N__11997));
    Odrv4 I__1147 (
            .O(N__11997),
            .I(M_this_oam_ram_write_data_2));
    CascadeMux I__1146 (
            .O(N__11994),
            .I(N__11991));
    CascadeBuf I__1145 (
            .O(N__11991),
            .I(N__11988));
    CascadeMux I__1144 (
            .O(N__11988),
            .I(N__11985));
    InMux I__1143 (
            .O(N__11985),
            .I(N__11982));
    LocalMux I__1142 (
            .O(N__11982),
            .I(N__11978));
    InMux I__1141 (
            .O(N__11981),
            .I(N__11975));
    Span4Mux_v I__1140 (
            .O(N__11978),
            .I(N__11972));
    LocalMux I__1139 (
            .O(N__11975),
            .I(M_this_map_address_qZ0Z_7));
    Odrv4 I__1138 (
            .O(N__11972),
            .I(M_this_map_address_qZ0Z_7));
    InMux I__1137 (
            .O(N__11967),
            .I(un1_M_this_map_address_q_cry_6));
    CascadeMux I__1136 (
            .O(N__11964),
            .I(N__11961));
    CascadeBuf I__1135 (
            .O(N__11961),
            .I(N__11958));
    CascadeMux I__1134 (
            .O(N__11958),
            .I(N__11955));
    InMux I__1133 (
            .O(N__11955),
            .I(N__11952));
    LocalMux I__1132 (
            .O(N__11952),
            .I(N__11948));
    InMux I__1131 (
            .O(N__11951),
            .I(N__11945));
    Span4Mux_v I__1130 (
            .O(N__11948),
            .I(N__11942));
    LocalMux I__1129 (
            .O(N__11945),
            .I(M_this_map_address_qZ0Z_8));
    Odrv4 I__1128 (
            .O(N__11942),
            .I(M_this_map_address_qZ0Z_8));
    InMux I__1127 (
            .O(N__11937),
            .I(bfn_9_25_0_));
    InMux I__1126 (
            .O(N__11934),
            .I(un1_M_this_map_address_q_cry_8));
    CascadeMux I__1125 (
            .O(N__11931),
            .I(N__11928));
    CascadeBuf I__1124 (
            .O(N__11928),
            .I(N__11925));
    CascadeMux I__1123 (
            .O(N__11925),
            .I(N__11922));
    InMux I__1122 (
            .O(N__11922),
            .I(N__11919));
    LocalMux I__1121 (
            .O(N__11919),
            .I(N__11915));
    InMux I__1120 (
            .O(N__11918),
            .I(N__11912));
    Span4Mux_v I__1119 (
            .O(N__11915),
            .I(N__11909));
    LocalMux I__1118 (
            .O(N__11912),
            .I(M_this_map_address_qZ0Z_9));
    Odrv4 I__1117 (
            .O(N__11909),
            .I(M_this_map_address_qZ0Z_9));
    InMux I__1116 (
            .O(N__11904),
            .I(N__11901));
    LocalMux I__1115 (
            .O(N__11901),
            .I(N__11898));
    Odrv4 I__1114 (
            .O(N__11898),
            .I(\this_vga_ramdac.i2_mux ));
    InMux I__1113 (
            .O(N__11895),
            .I(N__11892));
    LocalMux I__1112 (
            .O(N__11892),
            .I(N__11888));
    InMux I__1111 (
            .O(N__11891),
            .I(N__11885));
    Span4Mux_v I__1110 (
            .O(N__11888),
            .I(N__11878));
    LocalMux I__1109 (
            .O(N__11885),
            .I(N__11878));
    InMux I__1108 (
            .O(N__11884),
            .I(N__11875));
    InMux I__1107 (
            .O(N__11883),
            .I(N__11870));
    Span4Mux_h I__1106 (
            .O(N__11878),
            .I(N__11865));
    LocalMux I__1105 (
            .O(N__11875),
            .I(N__11865));
    InMux I__1104 (
            .O(N__11874),
            .I(N__11862));
    CascadeMux I__1103 (
            .O(N__11873),
            .I(N__11858));
    LocalMux I__1102 (
            .O(N__11870),
            .I(N__11855));
    Span4Mux_v I__1101 (
            .O(N__11865),
            .I(N__11850));
    LocalMux I__1100 (
            .O(N__11862),
            .I(N__11850));
    InMux I__1099 (
            .O(N__11861),
            .I(N__11847));
    InMux I__1098 (
            .O(N__11858),
            .I(N__11844));
    Odrv12 I__1097 (
            .O(N__11855),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    Odrv4 I__1096 (
            .O(N__11850),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    LocalMux I__1095 (
            .O(N__11847),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    LocalMux I__1094 (
            .O(N__11844),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    IoInMux I__1093 (
            .O(N__11835),
            .I(N__11832));
    LocalMux I__1092 (
            .O(N__11832),
            .I(N__11829));
    Odrv12 I__1091 (
            .O(N__11829),
            .I(rgb_c_5));
    InMux I__1090 (
            .O(N__11826),
            .I(N__11823));
    LocalMux I__1089 (
            .O(N__11823),
            .I(N_60_0));
    CascadeMux I__1088 (
            .O(N__11820),
            .I(N__11817));
    InMux I__1087 (
            .O(N__11817),
            .I(N__11814));
    LocalMux I__1086 (
            .O(N__11814),
            .I(N__11811));
    Span4Mux_h I__1085 (
            .O(N__11811),
            .I(N__11808));
    Odrv4 I__1084 (
            .O(N__11808),
            .I(M_this_vga_signals_address_5));
    CascadeMux I__1083 (
            .O(N__11805),
            .I(N__11802));
    InMux I__1082 (
            .O(N__11802),
            .I(N__11799));
    LocalMux I__1081 (
            .O(N__11799),
            .I(M_this_vga_signals_address_2));
    InMux I__1080 (
            .O(N__11796),
            .I(N__11793));
    LocalMux I__1079 (
            .O(N__11793),
            .I(N__11790));
    Odrv4 I__1078 (
            .O(N__11790),
            .I(N_816_0));
    InMux I__1077 (
            .O(N__11787),
            .I(N__11784));
    LocalMux I__1076 (
            .O(N__11784),
            .I(N__11780));
    CascadeMux I__1075 (
            .O(N__11783),
            .I(N__11777));
    Span4Mux_v I__1074 (
            .O(N__11780),
            .I(N__11774));
    InMux I__1073 (
            .O(N__11777),
            .I(N__11771));
    Odrv4 I__1072 (
            .O(N__11774),
            .I(\this_vga_ramdac.N_2612_reto ));
    LocalMux I__1071 (
            .O(N__11771),
            .I(\this_vga_ramdac.N_2612_reto ));
    CascadeMux I__1070 (
            .O(N__11766),
            .I(N__11763));
    CascadeBuf I__1069 (
            .O(N__11763),
            .I(N__11760));
    CascadeMux I__1068 (
            .O(N__11760),
            .I(N__11757));
    InMux I__1067 (
            .O(N__11757),
            .I(N__11754));
    LocalMux I__1066 (
            .O(N__11754),
            .I(N__11750));
    InMux I__1065 (
            .O(N__11753),
            .I(N__11747));
    Span4Mux_v I__1064 (
            .O(N__11750),
            .I(N__11744));
    LocalMux I__1063 (
            .O(N__11747),
            .I(M_this_map_address_qZ0Z_0));
    Odrv4 I__1062 (
            .O(N__11744),
            .I(M_this_map_address_qZ0Z_0));
    CascadeMux I__1061 (
            .O(N__11739),
            .I(N__11736));
    CascadeBuf I__1060 (
            .O(N__11736),
            .I(N__11733));
    CascadeMux I__1059 (
            .O(N__11733),
            .I(N__11730));
    InMux I__1058 (
            .O(N__11730),
            .I(N__11727));
    LocalMux I__1057 (
            .O(N__11727),
            .I(N__11723));
    InMux I__1056 (
            .O(N__11726),
            .I(N__11720));
    Span4Mux_v I__1055 (
            .O(N__11723),
            .I(N__11717));
    LocalMux I__1054 (
            .O(N__11720),
            .I(M_this_map_address_qZ0Z_1));
    Odrv4 I__1053 (
            .O(N__11717),
            .I(M_this_map_address_qZ0Z_1));
    InMux I__1052 (
            .O(N__11712),
            .I(un1_M_this_map_address_q_cry_0));
    CascadeMux I__1051 (
            .O(N__11709),
            .I(N__11706));
    CascadeBuf I__1050 (
            .O(N__11706),
            .I(N__11703));
    CascadeMux I__1049 (
            .O(N__11703),
            .I(N__11700));
    InMux I__1048 (
            .O(N__11700),
            .I(N__11696));
    InMux I__1047 (
            .O(N__11699),
            .I(N__11693));
    LocalMux I__1046 (
            .O(N__11696),
            .I(N__11690));
    LocalMux I__1045 (
            .O(N__11693),
            .I(N__11685));
    Span4Mux_v I__1044 (
            .O(N__11690),
            .I(N__11685));
    Odrv4 I__1043 (
            .O(N__11685),
            .I(M_this_map_address_qZ0Z_2));
    InMux I__1042 (
            .O(N__11682),
            .I(un1_M_this_map_address_q_cry_1));
    CascadeMux I__1041 (
            .O(N__11679),
            .I(N__11676));
    CascadeBuf I__1040 (
            .O(N__11676),
            .I(N__11673));
    CascadeMux I__1039 (
            .O(N__11673),
            .I(N__11670));
    InMux I__1038 (
            .O(N__11670),
            .I(N__11666));
    InMux I__1037 (
            .O(N__11669),
            .I(N__11663));
    LocalMux I__1036 (
            .O(N__11666),
            .I(N__11660));
    LocalMux I__1035 (
            .O(N__11663),
            .I(N__11655));
    Span4Mux_v I__1034 (
            .O(N__11660),
            .I(N__11655));
    Odrv4 I__1033 (
            .O(N__11655),
            .I(M_this_map_address_qZ0Z_3));
    InMux I__1032 (
            .O(N__11652),
            .I(un1_M_this_map_address_q_cry_2));
    CascadeMux I__1031 (
            .O(N__11649),
            .I(N__11646));
    CascadeBuf I__1030 (
            .O(N__11646),
            .I(N__11643));
    CascadeMux I__1029 (
            .O(N__11643),
            .I(N__11640));
    InMux I__1028 (
            .O(N__11640),
            .I(N__11637));
    LocalMux I__1027 (
            .O(N__11637),
            .I(N__11633));
    InMux I__1026 (
            .O(N__11636),
            .I(N__11630));
    Span4Mux_v I__1025 (
            .O(N__11633),
            .I(N__11627));
    LocalMux I__1024 (
            .O(N__11630),
            .I(M_this_map_address_qZ0Z_4));
    Odrv4 I__1023 (
            .O(N__11627),
            .I(M_this_map_address_qZ0Z_4));
    InMux I__1022 (
            .O(N__11622),
            .I(un1_M_this_map_address_q_cry_3));
    CascadeMux I__1021 (
            .O(N__11619),
            .I(N__11616));
    CascadeBuf I__1020 (
            .O(N__11616),
            .I(N__11613));
    CascadeMux I__1019 (
            .O(N__11613),
            .I(N__11610));
    InMux I__1018 (
            .O(N__11610),
            .I(N__11607));
    LocalMux I__1017 (
            .O(N__11607),
            .I(N__11603));
    InMux I__1016 (
            .O(N__11606),
            .I(N__11600));
    Span4Mux_v I__1015 (
            .O(N__11603),
            .I(N__11597));
    LocalMux I__1014 (
            .O(N__11600),
            .I(M_this_map_address_qZ0Z_5));
    Odrv4 I__1013 (
            .O(N__11597),
            .I(M_this_map_address_qZ0Z_5));
    InMux I__1012 (
            .O(N__11592),
            .I(un1_M_this_map_address_q_cry_4));
    CascadeMux I__1011 (
            .O(N__11589),
            .I(N__11586));
    CascadeBuf I__1010 (
            .O(N__11586),
            .I(N__11583));
    CascadeMux I__1009 (
            .O(N__11583),
            .I(N__11580));
    InMux I__1008 (
            .O(N__11580),
            .I(N__11577));
    LocalMux I__1007 (
            .O(N__11577),
            .I(N__11573));
    InMux I__1006 (
            .O(N__11576),
            .I(N__11570));
    Span4Mux_v I__1005 (
            .O(N__11573),
            .I(N__11567));
    LocalMux I__1004 (
            .O(N__11570),
            .I(M_this_map_address_qZ0Z_6));
    Odrv4 I__1003 (
            .O(N__11567),
            .I(M_this_map_address_qZ0Z_6));
    InMux I__1002 (
            .O(N__11562),
            .I(un1_M_this_map_address_q_cry_5));
    InMux I__1001 (
            .O(N__11559),
            .I(N__11556));
    LocalMux I__1000 (
            .O(N__11556),
            .I(N__11553));
    Odrv4 I__999 (
            .O(N__11553),
            .I(M_this_oam_ram_write_data_0));
    InMux I__998 (
            .O(N__11550),
            .I(N__11547));
    LocalMux I__997 (
            .O(N__11547),
            .I(N__11544));
    Span4Mux_h I__996 (
            .O(N__11544),
            .I(N__11541));
    Odrv4 I__995 (
            .O(N__11541),
            .I(\this_oam_ram.M_this_oam_ram_read_data_12 ));
    InMux I__994 (
            .O(N__11538),
            .I(N__11535));
    LocalMux I__993 (
            .O(N__11535),
            .I(\this_oam_ram.M_this_oam_ram_read_data_17 ));
    InMux I__992 (
            .O(N__11532),
            .I(N__11529));
    LocalMux I__991 (
            .O(N__11529),
            .I(M_this_oam_ram_read_data_i_17));
    InMux I__990 (
            .O(N__11526),
            .I(N__11523));
    LocalMux I__989 (
            .O(N__11523),
            .I(\this_oam_ram.M_this_oam_ram_read_data_18 ));
    InMux I__988 (
            .O(N__11520),
            .I(N__11517));
    LocalMux I__987 (
            .O(N__11517),
            .I(M_this_oam_ram_read_data_i_18));
    InMux I__986 (
            .O(N__11514),
            .I(N__11511));
    LocalMux I__985 (
            .O(N__11511),
            .I(\this_oam_ram.M_this_oam_ram_read_data_20 ));
    InMux I__984 (
            .O(N__11508),
            .I(N__11505));
    LocalMux I__983 (
            .O(N__11505),
            .I(M_this_oam_ram_read_data_i_20));
    InMux I__982 (
            .O(N__11502),
            .I(N__11496));
    InMux I__981 (
            .O(N__11501),
            .I(N__11496));
    LocalMux I__980 (
            .O(N__11496),
            .I(this_pixel_clk_M_counter_q_i_1));
    InMux I__979 (
            .O(N__11493),
            .I(N__11486));
    InMux I__978 (
            .O(N__11492),
            .I(N__11486));
    InMux I__977 (
            .O(N__11491),
            .I(N__11483));
    LocalMux I__976 (
            .O(N__11486),
            .I(N__11480));
    LocalMux I__975 (
            .O(N__11483),
            .I(this_pixel_clk_M_counter_q_0));
    Odrv4 I__974 (
            .O(N__11480),
            .I(this_pixel_clk_M_counter_q_0));
    IoInMux I__973 (
            .O(N__11475),
            .I(N__11472));
    LocalMux I__972 (
            .O(N__11472),
            .I(N__11469));
    Span12Mux_s8_h I__971 (
            .O(N__11469),
            .I(N__11466));
    Odrv12 I__970 (
            .O(N__11466),
            .I(rgb_c_1));
    CascadeMux I__969 (
            .O(N__11463),
            .I(N__11460));
    InMux I__968 (
            .O(N__11460),
            .I(N__11457));
    LocalMux I__967 (
            .O(N__11457),
            .I(N__11454));
    Span4Mux_v I__966 (
            .O(N__11454),
            .I(N__11451));
    Odrv4 I__965 (
            .O(N__11451),
            .I(M_this_vga_signals_address_1));
    InMux I__964 (
            .O(N__11448),
            .I(\this_ppu.un3_sprites_addr_cry_0 ));
    InMux I__963 (
            .O(N__11445),
            .I(\this_ppu.un3_sprites_addr_cry_1 ));
    InMux I__962 (
            .O(N__11442),
            .I(N__11439));
    LocalMux I__961 (
            .O(N__11439),
            .I(N__11436));
    Odrv4 I__960 (
            .O(N__11436),
            .I(M_this_oam_ram_read_data_i_19));
    InMux I__959 (
            .O(N__11433),
            .I(\this_ppu.un3_sprites_addr_cry_2 ));
    InMux I__958 (
            .O(N__11430),
            .I(\this_ppu.un3_sprites_addr_cry_3 ));
    InMux I__957 (
            .O(N__11427),
            .I(\this_ppu.un3_sprites_addr_cry_4 ));
    InMux I__956 (
            .O(N__11424),
            .I(\this_ppu.un3_sprites_addr_cry_5 ));
    CascadeMux I__955 (
            .O(N__11421),
            .I(N__11418));
    InMux I__954 (
            .O(N__11418),
            .I(N__11415));
    LocalMux I__953 (
            .O(N__11415),
            .I(N__11412));
    Odrv4 I__952 (
            .O(N__11412),
            .I(M_this_oam_ram_read_data_23));
    InMux I__951 (
            .O(N__11409),
            .I(\this_ppu.un3_sprites_addr_cry_6 ));
    InMux I__950 (
            .O(N__11406),
            .I(N__11403));
    LocalMux I__949 (
            .O(N__11403),
            .I(\this_oam_ram.M_this_oam_ram_read_data_21 ));
    InMux I__948 (
            .O(N__11400),
            .I(N__11397));
    LocalMux I__947 (
            .O(N__11397),
            .I(M_this_oam_ram_read_data_i_21));
    InMux I__946 (
            .O(N__11394),
            .I(N__11391));
    LocalMux I__945 (
            .O(N__11391),
            .I(N__11388));
    Odrv4 I__944 (
            .O(N__11388),
            .I(M_this_oam_ram_write_data_4));
    InMux I__943 (
            .O(N__11385),
            .I(N__11382));
    LocalMux I__942 (
            .O(N__11382),
            .I(N__11379));
    Odrv4 I__941 (
            .O(N__11379),
            .I(N_895_0));
    InMux I__940 (
            .O(N__11376),
            .I(N__11373));
    LocalMux I__939 (
            .O(N__11373),
            .I(N__11370));
    Odrv4 I__938 (
            .O(N__11370),
            .I(N_891_0));
    InMux I__937 (
            .O(N__11367),
            .I(N__11364));
    LocalMux I__936 (
            .O(N__11364),
            .I(\this_oam_ram.M_this_oam_ram_read_data_10 ));
    InMux I__935 (
            .O(N__11361),
            .I(N__11358));
    LocalMux I__934 (
            .O(N__11358),
            .I(\this_oam_ram.M_this_oam_ram_read_data_11 ));
    InMux I__933 (
            .O(N__11355),
            .I(N__11352));
    LocalMux I__932 (
            .O(N__11352),
            .I(M_this_oam_ram_write_data_28));
    InMux I__931 (
            .O(N__11349),
            .I(N__11346));
    LocalMux I__930 (
            .O(N__11346),
            .I(N__11343));
    Odrv4 I__929 (
            .O(N__11343),
            .I(N_894_0));
    InMux I__928 (
            .O(N__11340),
            .I(N__11337));
    LocalMux I__927 (
            .O(N__11337),
            .I(N_889_0));
    InMux I__926 (
            .O(N__11334),
            .I(N__11331));
    LocalMux I__925 (
            .O(N__11331),
            .I(\this_ppu.M_this_oam_ram_read_data_i_16 ));
    IoInMux I__924 (
            .O(N__11328),
            .I(N__11325));
    LocalMux I__923 (
            .O(N__11325),
            .I(N__11322));
    Span12Mux_s2_h I__922 (
            .O(N__11322),
            .I(N__11319));
    Odrv12 I__921 (
            .O(N__11319),
            .I(rgb_c_3));
    IoInMux I__920 (
            .O(N__11316),
            .I(N__11313));
    LocalMux I__919 (
            .O(N__11313),
            .I(N__11310));
    Span4Mux_s3_h I__918 (
            .O(N__11310),
            .I(N__11307));
    Span4Mux_v I__917 (
            .O(N__11307),
            .I(N__11304));
    Odrv4 I__916 (
            .O(N__11304),
            .I(rgb_c_4));
    InMux I__915 (
            .O(N__11301),
            .I(N__11298));
    LocalMux I__914 (
            .O(N__11298),
            .I(N__11295));
    Span4Mux_h I__913 (
            .O(N__11295),
            .I(N__11292));
    Odrv4 I__912 (
            .O(N__11292),
            .I(N_834_0));
    InMux I__911 (
            .O(N__11289),
            .I(N__11286));
    LocalMux I__910 (
            .O(N__11286),
            .I(N__11283));
    Odrv4 I__909 (
            .O(N__11283),
            .I(N_818_0));
    InMux I__908 (
            .O(N__11280),
            .I(N__11277));
    LocalMux I__907 (
            .O(N__11277),
            .I(N__11274));
    Span4Mux_v I__906 (
            .O(N__11274),
            .I(N__11271));
    Odrv4 I__905 (
            .O(N__11271),
            .I(N_837_0));
    InMux I__904 (
            .O(N__11268),
            .I(N__11265));
    LocalMux I__903 (
            .O(N__11265),
            .I(N__11262));
    Odrv4 I__902 (
            .O(N__11262),
            .I(M_this_oam_ram_write_data_5));
    InMux I__901 (
            .O(N__11259),
            .I(N__11256));
    LocalMux I__900 (
            .O(N__11256),
            .I(M_this_oam_ram_write_data_8));
    InMux I__899 (
            .O(N__11253),
            .I(N__11250));
    LocalMux I__898 (
            .O(N__11250),
            .I(N_836_0));
    InMux I__897 (
            .O(N__11247),
            .I(N__11244));
    LocalMux I__896 (
            .O(N__11244),
            .I(N_896_0));
    CascadeMux I__895 (
            .O(N__11241),
            .I(N__11238));
    CascadeBuf I__894 (
            .O(N__11238),
            .I(N__11235));
    CascadeMux I__893 (
            .O(N__11235),
            .I(N__11232));
    InMux I__892 (
            .O(N__11232),
            .I(N__11228));
    InMux I__891 (
            .O(N__11231),
            .I(N__11225));
    LocalMux I__890 (
            .O(N__11228),
            .I(N__11222));
    LocalMux I__889 (
            .O(N__11225),
            .I(M_this_oam_address_qZ0Z_4));
    Odrv4 I__888 (
            .O(N__11222),
            .I(M_this_oam_address_qZ0Z_4));
    InMux I__887 (
            .O(N__11217),
            .I(un1_M_this_oam_address_q_cry_3));
    InMux I__886 (
            .O(N__11214),
            .I(un1_M_this_oam_address_q_cry_4));
    CascadeMux I__885 (
            .O(N__11211),
            .I(N__11208));
    CascadeBuf I__884 (
            .O(N__11208),
            .I(N__11205));
    CascadeMux I__883 (
            .O(N__11205),
            .I(N__11202));
    InMux I__882 (
            .O(N__11202),
            .I(N__11199));
    LocalMux I__881 (
            .O(N__11199),
            .I(N__11195));
    InMux I__880 (
            .O(N__11198),
            .I(N__11192));
    Span4Mux_h I__879 (
            .O(N__11195),
            .I(N__11189));
    LocalMux I__878 (
            .O(N__11192),
            .I(M_this_oam_address_qZ0Z_5));
    Odrv4 I__877 (
            .O(N__11189),
            .I(M_this_oam_address_qZ0Z_5));
    InMux I__876 (
            .O(N__11184),
            .I(N__11181));
    LocalMux I__875 (
            .O(N__11181),
            .I(\this_oam_ram.M_this_oam_ram_read_data_19 ));
    InMux I__874 (
            .O(N__11178),
            .I(N__11175));
    LocalMux I__873 (
            .O(N__11175),
            .I(M_this_data_tmp_qZ0Z_26));
    InMux I__872 (
            .O(N__11172),
            .I(N__11169));
    LocalMux I__871 (
            .O(N__11169),
            .I(M_this_oam_ram_write_data_26));
    InMux I__870 (
            .O(N__11166),
            .I(N__11163));
    LocalMux I__869 (
            .O(N__11163),
            .I(M_this_oam_ram_write_data_20));
    InMux I__868 (
            .O(N__11160),
            .I(N__11157));
    LocalMux I__867 (
            .O(N__11157),
            .I(N_892_0));
    IoInMux I__866 (
            .O(N__11154),
            .I(N__11151));
    LocalMux I__865 (
            .O(N__11151),
            .I(N__11148));
    Span12Mux_s6_h I__864 (
            .O(N__11148),
            .I(N__11145));
    Span12Mux_v I__863 (
            .O(N__11145),
            .I(N__11142));
    Odrv12 I__862 (
            .O(N__11142),
            .I(rgb_c_0));
    IoInMux I__861 (
            .O(N__11139),
            .I(N__11136));
    LocalMux I__860 (
            .O(N__11136),
            .I(N__11133));
    Odrv12 I__859 (
            .O(N__11133),
            .I(this_vga_signals_vvisibility_i));
    InMux I__858 (
            .O(N__11130),
            .I(N__11127));
    LocalMux I__857 (
            .O(N__11127),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    IoInMux I__856 (
            .O(N__11124),
            .I(N__11121));
    LocalMux I__855 (
            .O(N__11121),
            .I(N__11118));
    Span4Mux_s1_h I__854 (
            .O(N__11118),
            .I(N__11115));
    Span4Mux_h I__853 (
            .O(N__11115),
            .I(N__11112));
    Odrv4 I__852 (
            .O(N__11112),
            .I(rgb_c_2));
    InMux I__851 (
            .O(N__11109),
            .I(N__11106));
    LocalMux I__850 (
            .O(N__11106),
            .I(N__11103));
    Odrv12 I__849 (
            .O(N__11103),
            .I(port_clk_c));
    InMux I__848 (
            .O(N__11100),
            .I(N__11097));
    LocalMux I__847 (
            .O(N__11097),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    CascadeMux I__846 (
            .O(N__11094),
            .I(N__11091));
    CascadeBuf I__845 (
            .O(N__11091),
            .I(N__11088));
    CascadeMux I__844 (
            .O(N__11088),
            .I(N__11085));
    InMux I__843 (
            .O(N__11085),
            .I(N__11082));
    LocalMux I__842 (
            .O(N__11082),
            .I(N__11078));
    InMux I__841 (
            .O(N__11081),
            .I(N__11075));
    Span4Mux_v I__840 (
            .O(N__11078),
            .I(N__11072));
    LocalMux I__839 (
            .O(N__11075),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__838 (
            .O(N__11072),
            .I(M_this_oam_address_qZ0Z_0));
    CascadeMux I__837 (
            .O(N__11067),
            .I(N__11064));
    CascadeBuf I__836 (
            .O(N__11064),
            .I(N__11061));
    CascadeMux I__835 (
            .O(N__11061),
            .I(N__11058));
    InMux I__834 (
            .O(N__11058),
            .I(N__11055));
    LocalMux I__833 (
            .O(N__11055),
            .I(N__11051));
    InMux I__832 (
            .O(N__11054),
            .I(N__11048));
    Span4Mux_v I__831 (
            .O(N__11051),
            .I(N__11045));
    LocalMux I__830 (
            .O(N__11048),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__829 (
            .O(N__11045),
            .I(M_this_oam_address_qZ0Z_1));
    InMux I__828 (
            .O(N__11040),
            .I(un1_M_this_oam_address_q_cry_0));
    CascadeMux I__827 (
            .O(N__11037),
            .I(N__11034));
    CascadeBuf I__826 (
            .O(N__11034),
            .I(N__11031));
    CascadeMux I__825 (
            .O(N__11031),
            .I(N__11028));
    InMux I__824 (
            .O(N__11028),
            .I(N__11024));
    InMux I__823 (
            .O(N__11027),
            .I(N__11021));
    LocalMux I__822 (
            .O(N__11024),
            .I(N__11018));
    LocalMux I__821 (
            .O(N__11021),
            .I(M_this_oam_address_qZ0Z_2));
    Odrv4 I__820 (
            .O(N__11018),
            .I(M_this_oam_address_qZ0Z_2));
    InMux I__819 (
            .O(N__11013),
            .I(un1_M_this_oam_address_q_cry_1));
    CascadeMux I__818 (
            .O(N__11010),
            .I(N__11007));
    CascadeBuf I__817 (
            .O(N__11007),
            .I(N__11004));
    CascadeMux I__816 (
            .O(N__11004),
            .I(N__11001));
    InMux I__815 (
            .O(N__11001),
            .I(N__10998));
    LocalMux I__814 (
            .O(N__10998),
            .I(N__10994));
    InMux I__813 (
            .O(N__10997),
            .I(N__10991));
    Span4Mux_h I__812 (
            .O(N__10994),
            .I(N__10988));
    LocalMux I__811 (
            .O(N__10991),
            .I(M_this_oam_address_qZ0Z_3));
    Odrv4 I__810 (
            .O(N__10988),
            .I(M_this_oam_address_qZ0Z_3));
    InMux I__809 (
            .O(N__10983),
            .I(un1_M_this_oam_address_q_cry_2));
    IoInMux I__808 (
            .O(N__10980),
            .I(N__10977));
    LocalMux I__807 (
            .O(N__10977),
            .I(N__10974));
    Span4Mux_s3_h I__806 (
            .O(N__10974),
            .I(N__10971));
    Span4Mux_v I__805 (
            .O(N__10971),
            .I(N__10968));
    Odrv4 I__804 (
            .O(N__10968),
            .I(port_nmib_0_i));
    defparam IN_MUX_bfv_23_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_17_0_));
    defparam IN_MUX_bfv_23_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_18_0_ (
            .carryinitin(un1_M_this_sprites_address_q_cry_7),
            .carryinitout(bfn_23_18_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_24_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_21_0_));
    defparam IN_MUX_bfv_24_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_22_0_ (
            .carryinitin(M_this_data_count_q_cry_7),
            .carryinitout(bfn_24_22_0_));
    defparam IN_MUX_bfv_21_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_20_0_));
    defparam IN_MUX_bfv_21_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_21_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_21_21_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(un1_M_this_map_address_q_cry_7),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_26_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_26_23_0_));
    defparam IN_MUX_bfv_26_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_24_0_ (
            .carryinitin(M_this_external_address_q_cry_7),
            .carryinitout(bfn_26_24_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNI4KCU6_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__16548),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_1358_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_9  (
            .USERSIGNALTOGLOBALBUFFER(N__15809),
            .GLOBALBUFFEROUTPUT(M_this_reset_cond_out_g_0));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI0JAO7_9_LC_5_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI0JAO7_9_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI0JAO7_9_LC_5_15_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI0JAO7_9_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__17735),
            .in2(_gnd_net_),
            .in3(N__15879),
            .lcout(port_nmib_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_0_9_LC_5_27_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_0_9_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_0_9_LC_5_27_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_0_9_LC_5_27_1  (
            .in0(N__15872),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_vvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_6_19_0 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_6_19_0 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_6_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_6_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11100),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32633),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_6_19_2 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_6_19_2 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_6_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_6_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11130),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32633),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_6_20_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_6_20_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_6_20_0  (
            .in0(_gnd_net_),
            .in1(N__11787),
            .in2(_gnd_net_),
            .in3(N__11895),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_6_20_6 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_6_20_6 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_6_20_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_6_20_6  (
            .in0(N__11109),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32636),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_0_LC_7_17_0.C_ON=1'b1;
    defparam M_this_oam_address_q_0_LC_7_17_0.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_0_LC_7_17_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_oam_address_q_0_LC_7_17_0 (
            .in0(N__26788),
            .in1(N__11081),
            .in2(N__18624),
            .in3(N__18619),
            .lcout(M_this_oam_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(un1_M_this_oam_address_q_cry_0),
            .clk(N__32616),
            .ce(),
            .sr(N__26071));
    defparam M_this_oam_address_q_1_LC_7_17_1.C_ON=1'b1;
    defparam M_this_oam_address_q_1_LC_7_17_1.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_1_LC_7_17_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_oam_address_q_1_LC_7_17_1 (
            .in0(N__26792),
            .in1(N__11054),
            .in2(_gnd_net_),
            .in3(N__11040),
            .lcout(M_this_oam_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_oam_address_q_cry_0),
            .carryout(un1_M_this_oam_address_q_cry_1),
            .clk(N__32616),
            .ce(),
            .sr(N__26071));
    defparam M_this_oam_address_q_2_LC_7_17_2.C_ON=1'b1;
    defparam M_this_oam_address_q_2_LC_7_17_2.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_2_LC_7_17_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_oam_address_q_2_LC_7_17_2 (
            .in0(N__26789),
            .in1(N__11027),
            .in2(_gnd_net_),
            .in3(N__11013),
            .lcout(M_this_oam_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_oam_address_q_cry_1),
            .carryout(un1_M_this_oam_address_q_cry_2),
            .clk(N__32616),
            .ce(),
            .sr(N__26071));
    defparam M_this_oam_address_q_3_LC_7_17_3.C_ON=1'b1;
    defparam M_this_oam_address_q_3_LC_7_17_3.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_3_LC_7_17_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_oam_address_q_3_LC_7_17_3 (
            .in0(N__26793),
            .in1(N__10997),
            .in2(_gnd_net_),
            .in3(N__10983),
            .lcout(M_this_oam_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_oam_address_q_cry_2),
            .carryout(un1_M_this_oam_address_q_cry_3),
            .clk(N__32616),
            .ce(),
            .sr(N__26071));
    defparam M_this_oam_address_q_4_LC_7_17_4.C_ON=1'b1;
    defparam M_this_oam_address_q_4_LC_7_17_4.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_4_LC_7_17_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_oam_address_q_4_LC_7_17_4 (
            .in0(N__26790),
            .in1(N__11231),
            .in2(_gnd_net_),
            .in3(N__11217),
            .lcout(M_this_oam_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_oam_address_q_cry_3),
            .carryout(un1_M_this_oam_address_q_cry_4),
            .clk(N__32616),
            .ce(),
            .sr(N__26071));
    defparam M_this_oam_address_q_5_LC_7_17_5.C_ON=1'b0;
    defparam M_this_oam_address_q_5_LC_7_17_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_5_LC_7_17_5.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_5_LC_7_17_5 (
            .in0(N__11198),
            .in1(N__26791),
            .in2(_gnd_net_),
            .in3(N__11214),
            .lcout(M_this_oam_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32616),
            .ce(),
            .sr(N__26071));
    defparam M_this_data_tmp_q_esr_26_LC_7_18_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_26_LC_7_18_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_26_LC_7_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_26_LC_7_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32919),
            .lcout(M_this_data_tmp_qZ0Z_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32620),
            .ce(N__17664),
            .sr(N__26070));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_7_19_0 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_7_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11184),
            .lcout(M_this_oam_ram_read_data_i_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_26_LC_7_19_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_26_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_26_LC_7_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_26_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__11178),
            .in2(_gnd_net_),
            .in3(N__18618),
            .lcout(M_this_oam_ram_write_data_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_20_LC_7_19_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_20_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_20_LC_7_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_20_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__12321),
            .in2(_gnd_net_),
            .in3(N__18617),
            .lcout(M_this_oam_ram_write_data_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_23_LC_7_20_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_23_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_23_LC_7_20_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_23_LC_7_20_6  (
            .in0(N__18620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12300),
            .lcout(N_892_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_0_LC_7_21_5 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_0_LC_7_21_5 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_0_LC_7_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clk.M_counter_q_0_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11491),
            .lcout(this_pixel_clk_M_counter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32637),
            .ce(),
            .sr(N__26064));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_7_22_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_7_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__11891),
            .in2(_gnd_net_),
            .in3(N__12351),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_7_25_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_7_25_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_7_25_0  (
            .in0(N__11884),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12648),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_7_26_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_7_26_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_7_26_2  (
            .in0(N__11874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12384),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_15_LC_9_15_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_15_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_15_LC_9_15_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_15_LC_9_15_0  (
            .in0(N__18576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12057),
            .lcout(N_834_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_14_LC_9_15_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_14_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_14_LC_9_15_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_14_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__12774),
            .in2(_gnd_net_),
            .in3(N__18575),
            .lcout(N_818_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_1_LC_9_16_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_1_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_1_LC_9_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_1_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__13644),
            .in2(_gnd_net_),
            .in3(N__18592),
            .lcout(N_837_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_5_LC_9_16_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_5_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_5_LC_9_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_5_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__13296),
            .in2(_gnd_net_),
            .in3(N__18591),
            .lcout(M_this_oam_ram_write_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_8_LC_9_17_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_8_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_8_LC_9_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_8_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__12051),
            .in2(_gnd_net_),
            .in3(N__18597),
            .lcout(M_this_oam_ram_write_data_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_7_LC_9_17_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_7_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_7_LC_9_17_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_7_LC_9_17_1  (
            .in0(N__18601),
            .in1(N__12747),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_836_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_11_LC_9_17_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_11_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_11_LC_9_17_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_11_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__12045),
            .in2(_gnd_net_),
            .in3(N__18598),
            .lcout(N_896_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_4_LC_9_17_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_4_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_4_LC_9_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_4_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__12732),
            .in2(_gnd_net_),
            .in3(N__18596),
            .lcout(M_this_oam_ram_write_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_13_LC_9_17_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_13_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_13_LC_9_17_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_13_LC_9_17_5  (
            .in0(N__18599),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13497),
            .lcout(N_895_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_27_LC_9_17_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_27_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_27_LC_9_17_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_27_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(N__12765),
            .in2(_gnd_net_),
            .in3(N__18600),
            .lcout(N_891_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_9_17_7 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_9_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11367),
            .lcout(M_this_oam_ram_read_data_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_1_LC_9_18_2 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_1_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_1_LC_9_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_0_RNISG75_1_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11361),
            .lcout(M_this_oam_ram_read_data_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_28_LC_9_18_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_28_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_28_LC_9_18_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_28_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__12930),
            .in2(_gnd_net_),
            .in3(N__18608),
            .lcout(M_this_oam_ram_write_data_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_19_LC_9_18_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_19_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_19_LC_9_18_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_19_LC_9_18_5  (
            .in0(N__18609),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12201),
            .lcout(N_894_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_31_LC_9_18_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_31_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_31_LC_9_18_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_31_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__12717),
            .in2(_gnd_net_),
            .in3(N__18610),
            .lcout(N_889_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un3_sprites_addr_cry_0_c_inv_LC_9_19_0 .C_ON=1'b1;
    defparam \this_ppu.un3_sprites_addr_cry_0_c_inv_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un3_sprites_addr_cry_0_c_inv_LC_9_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un3_sprites_addr_cry_0_c_inv_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__11334),
            .in2(N__19318),
            .in3(N__12902),
            .lcout(\this_ppu.M_this_oam_ram_read_data_i_16 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\this_ppu.un3_sprites_addr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un3_sprites_addr_cry_0_c_RNIRLA8_LC_9_19_1 .C_ON=1'b1;
    defparam \this_ppu.un3_sprites_addr_cry_0_c_RNIRLA8_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un3_sprites_addr_cry_0_c_RNIRLA8_LC_9_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un3_sprites_addr_cry_0_c_RNIRLA8_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__11532),
            .in2(N__20926),
            .in3(N__11448),
            .lcout(\this_ppu.un3_sprites_addr_cry_0_c_RNIRLAZ0Z8 ),
            .ltout(),
            .carryin(\this_ppu.un3_sprites_addr_cry_0 ),
            .carryout(\this_ppu.un3_sprites_addr_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un3_sprites_addr_cry_1_c_RNITOB8_LC_9_19_2 .C_ON=1'b1;
    defparam \this_ppu.un3_sprites_addr_cry_1_c_RNITOB8_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un3_sprites_addr_cry_1_c_RNITOB8_LC_9_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un3_sprites_addr_cry_1_c_RNITOB8_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__11520),
            .in2(N__13880),
            .in3(N__11445),
            .lcout(\this_ppu.un3_sprites_addr_cry_1_c_RNITOBZ0Z8 ),
            .ltout(),
            .carryin(\this_ppu.un3_sprites_addr_cry_1 ),
            .carryout(\this_ppu.un3_sprites_addr_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un3_sprites_addr_cry_2_c_RNIVRC8_LC_9_19_3 .C_ON=1'b1;
    defparam \this_ppu.un3_sprites_addr_cry_2_c_RNIVRC8_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un3_sprites_addr_cry_2_c_RNIVRC8_LC_9_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un3_sprites_addr_cry_2_c_RNIVRC8_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__11442),
            .in2(N__13945),
            .in3(N__11433),
            .lcout(\this_ppu.un3_sprites_addr_cry_2_c_RNIVRCZ0Z8 ),
            .ltout(),
            .carryin(\this_ppu.un3_sprites_addr_cry_2 ),
            .carryout(\this_ppu.un3_sprites_addr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un3_sprites_addr_cry_3_c_RNI1VD8_LC_9_19_4 .C_ON=1'b1;
    defparam \this_ppu.un3_sprites_addr_cry_3_c_RNI1VD8_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un3_sprites_addr_cry_3_c_RNI1VD8_LC_9_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un3_sprites_addr_cry_3_c_RNI1VD8_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__11508),
            .in2(N__13813),
            .in3(N__11430),
            .lcout(\this_ppu.un3_sprites_addr_cry_3_c_RNI1VDZ0Z8 ),
            .ltout(),
            .carryin(\this_ppu.un3_sprites_addr_cry_3 ),
            .carryout(\this_ppu.un3_sprites_addr_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un3_sprites_addr_cry_4_c_RNI32F8_LC_9_19_5 .C_ON=1'b1;
    defparam \this_ppu.un3_sprites_addr_cry_4_c_RNI32F8_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un3_sprites_addr_cry_4_c_RNI32F8_LC_9_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un3_sprites_addr_cry_4_c_RNI32F8_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__11400),
            .in2(N__13576),
            .in3(N__11427),
            .lcout(\this_ppu.un3_sprites_addr_cry_4_c_RNI32FZ0Z8 ),
            .ltout(),
            .carryin(\this_ppu.un3_sprites_addr_cry_4 ),
            .carryout(\this_ppu.un3_sprites_addr_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un3_sprites_addr_cry_5_c_RNI55G8_LC_9_19_6 .C_ON=1'b1;
    defparam \this_ppu.un3_sprites_addr_cry_5_c_RNI55G8_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un3_sprites_addr_cry_5_c_RNI55G8_LC_9_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un3_sprites_addr_cry_5_c_RNI55G8_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__12878),
            .in2(N__12279),
            .in3(N__11424),
            .lcout(\this_ppu.un3_sprites_addr_cry_5_c_RNI55GZ0Z8 ),
            .ltout(),
            .carryin(\this_ppu.un3_sprites_addr_cry_5 ),
            .carryout(\this_ppu.un3_sprites_addr_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un3_sprites_addr_cry_6_c_RNIP5L8_LC_9_19_7 .C_ON=1'b0;
    defparam \this_ppu.un3_sprites_addr_cry_6_c_RNIP5L8_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un3_sprites_addr_cry_6_c_RNIP5L8_LC_9_19_7 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_ppu.un3_sprites_addr_cry_6_c_RNIP5L8_LC_9_19_7  (
            .in0(N__12827),
            .in1(_gnd_net_),
            .in2(N__11421),
            .in3(N__11409),
            .lcout(\this_ppu.un3_sprites_addr_cry_6_c_RNIP5LZ0Z8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m2_LC_9_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m2_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m2_LC_9_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m2_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__22928),
            .in2(_gnd_net_),
            .in3(N__21578),
            .lcout(\this_vga_signals.if_m2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_3_LC_9_20_1 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_3_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_3_LC_9_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_3_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11406),
            .lcout(M_this_oam_ram_read_data_i_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_0_LC_9_20_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_0_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_0_LC_9_20_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_0_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__13479),
            .in2(_gnd_net_),
            .in3(N__18623),
            .lcout(M_this_oam_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_2_LC_9_20_3 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_2_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_2_LC_9_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_0_RNISG75_2_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11550),
            .lcout(M_this_oam_ram_read_data_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_9_20_4 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_9_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11538),
            .lcout(M_this_oam_ram_read_data_i_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_9_20_5 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_9_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11526),
            .lcout(M_this_oam_ram_read_data_i_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_9_20_7 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_9_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11514),
            .lcout(M_this_oam_ram_read_data_i_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_1_LC_9_21_1 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_1_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_1_LC_9_21_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clk.M_counter_q_1_LC_9_21_1  (
            .in0(N__11502),
            .in1(N__11493),
            .in2(_gnd_net_),
            .in3(N__26181),
            .lcout(this_pixel_clk_M_counter_q_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32630),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.G_442_LC_9_21_5 .C_ON=1'b0;
    defparam \this_start_data_delay.G_442_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.G_442_LC_9_21_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_start_data_delay.G_442_LC_9_21_5  (
            .in0(N__11501),
            .in1(N__11492),
            .in2(_gnd_net_),
            .in3(N__26180),
            .lcout(G_442),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_9_22_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_9_22_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_9_22_0  (
            .in0(N__12363),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11883),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI946123_9_LC_9_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI946123_9_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI946123_9_LC_9_22_4 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI946123_9_LC_9_22_4  (
            .in0(N__13146),
            .in1(N__17129),
            .in2(_gnd_net_),
            .in3(N__13131),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI6B7F1_LC_9_22_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI6B7F1_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI6B7F1_LC_9_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI6B7F1_LC_9_22_6  (
            .in0(N__32896),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19891),
            .lcout(N_816_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_23_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_23_5 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_23_5  (
            .in0(N__11904),
            .in1(N__15822),
            .in2(N__11783),
            .in3(N__12670),
            .lcout(\this_vga_ramdac.N_2612_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32638),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_0_LC_9_24_0.C_ON=1'b1;
    defparam M_this_map_address_q_0_LC_9_24_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_0_LC_9_24_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_0_LC_9_24_0 (
            .in0(N__24041),
            .in1(N__11753),
            .in2(N__19896),
            .in3(N__19887),
            .lcout(M_this_map_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(un1_M_this_map_address_q_cry_0),
            .clk(N__32643),
            .ce(),
            .sr(N__26050));
    defparam M_this_map_address_q_1_LC_9_24_1.C_ON=1'b1;
    defparam M_this_map_address_q_1_LC_9_24_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_1_LC_9_24_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_1_LC_9_24_1 (
            .in0(N__24046),
            .in1(N__11726),
            .in2(_gnd_net_),
            .in3(N__11712),
            .lcout(M_this_map_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_0),
            .carryout(un1_M_this_map_address_q_cry_1),
            .clk(N__32643),
            .ce(),
            .sr(N__26050));
    defparam M_this_map_address_q_2_LC_9_24_2.C_ON=1'b1;
    defparam M_this_map_address_q_2_LC_9_24_2.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_2_LC_9_24_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_2_LC_9_24_2 (
            .in0(N__24042),
            .in1(N__11699),
            .in2(_gnd_net_),
            .in3(N__11682),
            .lcout(M_this_map_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_1),
            .carryout(un1_M_this_map_address_q_cry_2),
            .clk(N__32643),
            .ce(),
            .sr(N__26050));
    defparam M_this_map_address_q_3_LC_9_24_3.C_ON=1'b1;
    defparam M_this_map_address_q_3_LC_9_24_3.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_3_LC_9_24_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_3_LC_9_24_3 (
            .in0(N__24047),
            .in1(N__11669),
            .in2(_gnd_net_),
            .in3(N__11652),
            .lcout(M_this_map_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_2),
            .carryout(un1_M_this_map_address_q_cry_3),
            .clk(N__32643),
            .ce(),
            .sr(N__26050));
    defparam M_this_map_address_q_4_LC_9_24_4.C_ON=1'b1;
    defparam M_this_map_address_q_4_LC_9_24_4.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_4_LC_9_24_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_4_LC_9_24_4 (
            .in0(N__24043),
            .in1(N__11636),
            .in2(_gnd_net_),
            .in3(N__11622),
            .lcout(M_this_map_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_3),
            .carryout(un1_M_this_map_address_q_cry_4),
            .clk(N__32643),
            .ce(),
            .sr(N__26050));
    defparam M_this_map_address_q_5_LC_9_24_5.C_ON=1'b1;
    defparam M_this_map_address_q_5_LC_9_24_5.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_5_LC_9_24_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_5_LC_9_24_5 (
            .in0(N__24048),
            .in1(N__11606),
            .in2(_gnd_net_),
            .in3(N__11592),
            .lcout(M_this_map_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_4),
            .carryout(un1_M_this_map_address_q_cry_5),
            .clk(N__32643),
            .ce(),
            .sr(N__26050));
    defparam M_this_map_address_q_6_LC_9_24_6.C_ON=1'b1;
    defparam M_this_map_address_q_6_LC_9_24_6.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_6_LC_9_24_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_6_LC_9_24_6 (
            .in0(N__24044),
            .in1(N__11576),
            .in2(_gnd_net_),
            .in3(N__11562),
            .lcout(M_this_map_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_5),
            .carryout(un1_M_this_map_address_q_cry_6),
            .clk(N__32643),
            .ce(),
            .sr(N__26050));
    defparam M_this_map_address_q_7_LC_9_24_7.C_ON=1'b1;
    defparam M_this_map_address_q_7_LC_9_24_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_7_LC_9_24_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_7_LC_9_24_7 (
            .in0(N__24045),
            .in1(N__11981),
            .in2(_gnd_net_),
            .in3(N__11967),
            .lcout(M_this_map_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_6),
            .carryout(un1_M_this_map_address_q_cry_7),
            .clk(N__32643),
            .ce(),
            .sr(N__26050));
    defparam M_this_map_address_q_8_LC_9_25_0.C_ON=1'b1;
    defparam M_this_map_address_q_8_LC_9_25_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_8_LC_9_25_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_8_LC_9_25_0 (
            .in0(N__24038),
            .in1(N__11951),
            .in2(_gnd_net_),
            .in3(N__11937),
            .lcout(M_this_map_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(un1_M_this_map_address_q_cry_8),
            .clk(N__32647),
            .ce(),
            .sr(N__26047));
    defparam M_this_map_address_q_9_LC_9_25_1.C_ON=1'b0;
    defparam M_this_map_address_q_9_LC_9_25_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_9_LC_9_25_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_map_address_q_9_LC_9_25_1 (
            .in0(N__11918),
            .in1(N__24039),
            .in2(_gnd_net_),
            .in3(N__11934),
            .lcout(M_this_map_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32647),
            .ce(),
            .sr(N__26047));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_26_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_26_2 .LUT_INIT=16'b0001010100111101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_26_2  (
            .in0(N__12453),
            .in1(N__12496),
            .in2(N__12556),
            .in3(N__12583),
            .lcout(\this_vga_ramdac.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_26_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_26_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_26_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_q_ret_LC_9_26_5  (
            .in0(N__15817),
            .in1(N__17128),
            .in2(N__11873),
            .in3(N__12681),
            .lcout(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32651),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_9_27_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_9_27_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_9_27_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_9_27_6  (
            .in0(N__12699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11861),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIAF7F1_LC_9_28_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIAF7F1_LC_9_28_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIAF7F1_LC_9_28_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIAF7F1_LC_9_28_2  (
            .in0(N__28191),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19897),
            .lcout(N_60_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIT1827_9_LC_9_28_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIT1827_9_LC_9_28_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIT1827_9_LC_9_28_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIT1827_9_LC_9_28_3  (
            .in0(_gnd_net_),
            .in1(N__17119),
            .in2(_gnd_net_),
            .in3(N__13104),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI0MGR61_9_LC_9_28_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI0MGR61_9_LC_9_28_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI0MGR61_9_LC_9_28_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI0MGR61_9_LC_9_28_5  (
            .in0(_gnd_net_),
            .in1(N__17118),
            .in2(_gnd_net_),
            .in3(N__13179),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI7CFM8_9_LC_9_29_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI7CFM8_9_LC_9_29_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI7CFM8_9_LC_9_29_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI7CFM8_9_LC_9_29_0  (
            .in0(_gnd_net_),
            .in1(N__17121),
            .in2(_gnd_net_),
            .in3(N__13053),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIPFB21_2_LC_9_31_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIPFB21_2_LC_9_31_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIPFB21_2_LC_9_31_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \this_ppu.M_state_q_RNIPFB21_2_LC_9_31_7  (
            .in0(N__12186),
            .in1(N__32119),
            .in2(N__31971),
            .in3(N__12174),
            .lcout(M_this_ppu_sprites_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_15_LC_10_15_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_15_LC_10_15_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_15_LC_10_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_15_LC_10_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27907),
            .lcout(M_this_data_tmp_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32560),
            .ce(N__17357),
            .sr(N__26069));
    defparam M_this_data_tmp_q_esr_8_LC_10_16_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_8_LC_10_16_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_8_LC_10_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_8_LC_10_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28469),
            .lcout(M_this_data_tmp_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32569),
            .ce(N__17353),
            .sr(N__26067));
    defparam M_this_data_tmp_q_esr_11_LC_10_16_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_11_LC_10_16_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_11_LC_10_16_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_11_LC_10_16_6 (
            .in0(N__31356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32569),
            .ce(N__17353),
            .sr(N__26067));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_9_LC_10_17_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_9_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_9_LC_10_17_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_9_LC_10_17_0  (
            .in0(N__13488),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18582),
            .lcout(N_835_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_3_LC_10_17_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_3_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_3_LC_10_17_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_3_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__12753),
            .in2(_gnd_net_),
            .in3(N__18580),
            .lcout(N_897_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_6_LC_10_17_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_6_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_6_LC_10_17_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_6_LC_10_17_3  (
            .in0(N__18581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14142),
            .lcout(N_53_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_2_LC_10_17_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_2_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_2_LC_10_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_2_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__12738),
            .in2(_gnd_net_),
            .in3(N__18578),
            .lcout(M_this_oam_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_29_LC_10_17_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_29_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_29_LC_10_17_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_29_LC_10_17_5  (
            .in0(N__18579),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13308),
            .lcout(N_890_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_12_LC_10_17_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_12_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_12_LC_10_17_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_12_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__13287),
            .in2(_gnd_net_),
            .in3(N__18577),
            .lcout(M_this_oam_ram_write_data_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_25_LC_10_18_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_25_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_25_LC_10_18_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_25_LC_10_18_1  (
            .in0(N__18590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12723),
            .lcout(N_831_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_24_LC_10_18_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_24_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_24_LC_10_18_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_24_LC_10_18_3  (
            .in0(N__18587),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13635),
            .lcout(M_this_oam_ram_write_data_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_22_LC_10_18_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_22_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_22_LC_10_18_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_22_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__12306),
            .in2(_gnd_net_),
            .in3(N__18589),
            .lcout(N_832_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_21_LC_10_18_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_21_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_21_LC_10_18_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_21_LC_10_18_7  (
            .in0(N__18588),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12312),
            .lcout(N_893_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_16_LC_10_19_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_16_LC_10_19_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_16_LC_10_19_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_16_LC_10_19_0 (
            .in0(N__28468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32597),
            .ce(N__15957),
            .sr(N__26058));
    defparam M_this_data_tmp_q_esr_18_LC_10_19_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_18_LC_10_19_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_18_LC_10_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_18_LC_10_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32908),
            .lcout(M_this_data_tmp_qZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32597),
            .ce(N__15957),
            .sr(N__26058));
    defparam M_this_data_tmp_q_esr_19_LC_10_19_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_19_LC_10_19_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_19_LC_10_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_19_LC_10_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31357),
            .lcout(M_this_data_tmp_qZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32597),
            .ce(N__15957),
            .sr(N__26058));
    defparam M_this_data_tmp_q_esr_20_LC_10_19_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_20_LC_10_19_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_20_LC_10_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_20_LC_10_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28266),
            .lcout(M_this_data_tmp_qZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32597),
            .ce(N__15957),
            .sr(N__26058));
    defparam M_this_data_tmp_q_esr_21_LC_10_19_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_21_LC_10_19_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_21_LC_10_19_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_21_LC_10_19_5 (
            .in0(N__24463),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32597),
            .ce(N__15957),
            .sr(N__26058));
    defparam M_this_data_tmp_q_esr_22_LC_10_19_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_22_LC_10_19_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_22_LC_10_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_22_LC_10_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28190),
            .lcout(M_this_data_tmp_qZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32597),
            .ce(N__15957),
            .sr(N__26058));
    defparam M_this_data_tmp_q_esr_23_LC_10_19_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_23_LC_10_19_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_23_LC_10_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_23_LC_10_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27911),
            .lcout(M_this_data_tmp_qZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32597),
            .ce(N__15957),
            .sr(N__26058));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_2_LC_10_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_2_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_2_LC_10_20_3 .LUT_INIT=16'b1010011010010101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_2_LC_10_20_3  (
            .in0(N__12998),
            .in1(N__12411),
            .in2(N__14622),
            .in3(N__12974),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_4_LC_10_20_7 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_4_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_4_LC_10_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_4_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12288),
            .lcout(M_this_oam_ram_read_data_i_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIUULS4_3_LC_10_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIUULS4_3_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIUULS4_3_LC_10_21_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIUULS4_3_LC_10_21_0  (
            .in0(N__14480),
            .in1(_gnd_net_),
            .in2(N__14550),
            .in3(N__13041),
            .lcout(\this_vga_signals.M_hcounter_q_RNIUULS4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_10_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_10_21_2 .LUT_INIT=16'b1001001111001001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_10_21_2  (
            .in0(N__14481),
            .in1(N__13083),
            .in2(N__14551),
            .in3(N__13042),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_21_4 .LUT_INIT=16'b1001101110001001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_21_4  (
            .in0(N__14478),
            .in1(N__13082),
            .in2(N__14549),
            .in3(N__13039),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_21_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_21_5  (
            .in0(N__13040),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14479),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_10_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_10_21_6 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \this_vga_signals.un4_haddress_if_m2_0_LC_10_21_6  (
            .in0(N__14535),
            .in1(N__13390),
            .in2(N__12414),
            .in3(N__13364),
            .lcout(\this_vga_signals.if_m2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBG7F1_LC_10_22_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBG7F1_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBG7F1_LC_10_22_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBG7F1_LC_10_22_1  (
            .in0(N__27912),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19868),
            .lcout(N_58_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIR5V44_0_LC_10_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIR5V44_0_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIR5V44_0_LC_10_23_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNIR5V44_0_LC_10_23_1  (
            .in0(N__21497),
            .in1(N__13708),
            .in2(_gnd_net_),
            .in3(N__13248),
            .lcout(N_3_0),
            .ltout(N_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.G_480_LC_10_23_2 .C_ON=1'b0;
    defparam \this_start_data_delay.G_480_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.G_480_LC_10_23_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \this_start_data_delay.G_480_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__12708),
            .in2(N__12390),
            .in3(N__12330),
            .lcout(G_480),
            .ltout(G_480_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_10_23_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_10_23_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_10_23_3 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_10_23_3  (
            .in0(N__12380),
            .in1(N__12612),
            .in2(N__12387),
            .in3(N__15814),
            .lcout(\this_vga_ramdac.N_2614_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32631),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_10_23_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_10_23_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_10_23_4 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_10_23_4  (
            .in0(N__12669),
            .in1(N__12362),
            .in2(N__15821),
            .in3(N__12423),
            .lcout(\this_vga_ramdac.N_2611_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32631),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_10_23_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_10_23_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_10_23_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_10_23_5  (
            .in0(N__12621),
            .in1(N__15810),
            .in2(N__12347),
            .in3(N__12668),
            .lcout(\this_vga_ramdac.N_2610_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32631),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_RNIIQFU3_1_LC_10_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_RNIIQFU3_1_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_RNIIQFU3_1_LC_10_23_6 .LUT_INIT=16'b0001000010101010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_RNIIQFU3_1_LC_10_23_6  (
            .in0(N__13732),
            .in1(N__21663),
            .in2(N__13710),
            .in3(N__21496),
            .lcout(N_2_0),
            .ltout(N_2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_10_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_10_23_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_10_23_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_2_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12324),
            .in3(N__13260),
            .lcout(M_this_vga_signals_pixel_clk_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32631),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_10_25_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_10_25_1 .LUT_INIT=16'b0100011100100101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_10_25_1  (
            .in0(N__12462),
            .in1(N__12505),
            .in2(N__12558),
            .in3(N__12603),
            .lcout(),
            .ltout(\this_vga_ramdac.i2_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_10_25_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_10_25_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_10_25_2 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_10_25_2  (
            .in0(N__12680),
            .in1(N__15816),
            .in2(N__12702),
            .in3(N__12695),
            .lcout(\this_vga_ramdac.N_2615_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32639),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_10_25_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_10_25_4 .LUT_INIT=16'b0100101100010111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_10_25_4  (
            .in0(N__12602),
            .in1(N__12552),
            .in2(N__12507),
            .in3(N__12461),
            .lcout(),
            .ltout(\this_vga_ramdac.m16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_10_25_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_10_25_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_10_25_5 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_10_25_5  (
            .in0(N__12644),
            .in1(N__15815),
            .in2(N__12684),
            .in3(N__12679),
            .lcout(\this_vga_ramdac.N_2613_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32639),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI497F1_LC_10_25_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI497F1_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI497F1_LC_10_25_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI497F1_LC_10_25_6  (
            .in0(_gnd_net_),
            .in1(N__28395),
            .in2(_gnd_net_),
            .in3(N__19883),
            .lcout(N_73_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_10_25_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_10_25_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_10_25_7 .LUT_INIT=16'b0101010100100010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_10_25_7  (
            .in0(N__12551),
            .in1(N__12501),
            .in2(_gnd_net_),
            .in3(N__12601),
            .lcout(\this_vga_ramdac.N_24_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_10_26_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_10_26_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_10_26_0 .LUT_INIT=16'b0110010100101011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_10_26_0  (
            .in0(N__12454),
            .in1(N__12497),
            .in2(N__12557),
            .in3(N__12592),
            .lcout(\this_vga_ramdac.m19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_10_26_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_10_26_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_10_26_3 .LUT_INIT=16'b0000001111101111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_10_26_3  (
            .in0(N__12593),
            .in1(N__12550),
            .in2(N__12506),
            .in3(N__12455),
            .lcout(\this_vga_ramdac.m6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_14_LC_11_15_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_14_LC_11_15_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_14_LC_11_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_14_LC_11_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28179),
            .lcout(M_this_data_tmp_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32549),
            .ce(N__17361),
            .sr(N__26068));
    defparam M_this_data_tmp_q_esr_27_LC_11_16_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_27_LC_11_16_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_27_LC_11_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_27_LC_11_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31359),
            .lcout(M_this_data_tmp_qZ0Z_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32561),
            .ce(N__17645),
            .sr(N__26065));
    defparam M_this_data_tmp_q_esr_30_LC_11_16_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_30_LC_11_16_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_30_LC_11_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_30_LC_11_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28189),
            .lcout(M_this_data_tmp_qZ0Z_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32561),
            .ce(N__17645),
            .sr(N__26065));
    defparam M_this_data_tmp_q_esr_3_LC_11_17_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_3_LC_11_17_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_3_LC_11_17_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_3_LC_11_17_1 (
            .in0(N__31358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32570),
            .ce(N__16521),
            .sr(N__26062));
    defparam M_this_data_tmp_q_esr_7_LC_11_17_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_7_LC_11_17_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_7_LC_11_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_7_LC_11_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27945),
            .lcout(M_this_data_tmp_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32570),
            .ce(N__16521),
            .sr(N__26062));
    defparam M_this_data_tmp_q_esr_2_LC_11_17_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_2_LC_11_17_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_2_LC_11_17_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_2_LC_11_17_4 (
            .in0(N__32915),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32570),
            .ce(N__16521),
            .sr(N__26062));
    defparam M_this_data_tmp_q_esr_4_LC_11_17_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_4_LC_11_17_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_4_LC_11_17_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_4_LC_11_17_5 (
            .in0(N__28325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32570),
            .ce(N__16521),
            .sr(N__26062));
    defparam M_this_data_tmp_q_esr_25_LC_11_18_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_25_LC_11_18_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_25_LC_11_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_25_LC_11_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30928),
            .lcout(M_this_data_tmp_qZ0Z_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32580),
            .ce(N__17659),
            .sr(N__26059));
    defparam M_this_data_tmp_q_esr_31_LC_11_18_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_31_LC_11_18_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_31_LC_11_18_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 M_this_data_tmp_q_esr_31_LC_11_18_6 (
            .in0(_gnd_net_),
            .in1(N__27937),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32580),
            .ce(N__17659),
            .sr(N__26059));
    defparam M_this_data_tmp_q_esr_28_LC_11_18_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_28_LC_11_18_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_28_LC_11_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_28_LC_11_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28326),
            .lcout(M_this_data_tmp_qZ0Z_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32580),
            .ce(N__17659),
            .sr(N__26059));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_17_LC_11_19_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_17_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_17_LC_11_19_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_17_LC_11_19_0  (
            .in0(N__18585),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15396),
            .lcout(N_833_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI98B5_0_LC_11_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI98B5_0_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI98B5_0_LC_11_19_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_ppu.M_haddress_q_RNI98B5_0_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__19311),
            .in2(_gnd_net_),
            .in3(N__12909),
            .lcout(\this_ppu.un3_sprites_addr_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIIT3_6_LC_11_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIIT3_6_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIIT3_6_LC_11_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.M_haddress_q_RNIIT3_6_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13604),
            .lcout(M_this_ppu_vram_addr_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_18_LC_11_19_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_18_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_18_LC_11_19_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_18_LC_11_19_4  (
            .in0(N__18584),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12861),
            .lcout(M_this_oam_ram_write_data_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI5S7_7_LC_11_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI5S7_7_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI5S7_7_LC_11_19_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_ppu.M_haddress_q_RNI5S7_7_LC_11_19_5  (
            .in0(N__13605),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13526),
            .lcout(M_this_ppu_map_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_30_LC_11_19_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_30_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_i_30_LC_11_19_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_i_30_LC_11_19_6  (
            .in0(N__18586),
            .in1(N__12810),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_830_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_16_LC_11_19_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_16_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_16_LC_11_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_16_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__12792),
            .in2(_gnd_net_),
            .in3(N__18583),
            .lcout(M_this_oam_ram_write_data_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIB0ACH_2_LC_11_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIB0ACH_2_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIB0ACH_2_LC_11_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIB0ACH_2_LC_11_20_0  (
            .in0(N__13363),
            .in1(N__14612),
            .in2(N__13394),
            .in3(N__14552),
            .lcout(\this_vga_signals.d_N_3_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_11_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_11_20_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__13386),
            .in2(_gnd_net_),
            .in3(N__13362),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m4_LC_11_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m4_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m4_LC_11_20_2 .LUT_INIT=16'b0000011001100000;
    LogicCell40 \this_vga_signals.un4_haddress_if_m4_LC_11_20_2  (
            .in0(N__14599),
            .in1(N__14798),
            .in2(N__13011),
            .in3(N__14553),
            .lcout(),
            .ltout(\this_vga_signals.if_i4_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_LC_11_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_LC_11_20_3 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_LC_11_20_3  (
            .in0(N__12997),
            .in1(N__13008),
            .in2(N__13002),
            .in3(N__12947),
            .lcout(\this_vga_signals.mult1_un82_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_11_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_11_20_4 .LUT_INIT=16'b1010100110100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_11_20_4  (
            .in0(N__12999),
            .in1(N__12981),
            .in2(N__12960),
            .in3(N__12975),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c2_LC_11_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c2_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c2_LC_11_20_5 .LUT_INIT=16'b0101111100000101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c2_LC_11_20_5  (
            .in0(N__14799),
            .in1(_gnd_net_),
            .in2(N__12963),
            .in3(N__14600),
            .lcout(\this_vga_signals.mult1_un82_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m2_2_LC_11_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m2_2_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m2_2_LC_11_20_6 .LUT_INIT=16'b0001001001001000;
    LogicCell40 \this_vga_signals.un4_haddress_if_m2_2_LC_11_20_6  (
            .in0(N__14547),
            .in1(N__14473),
            .in2(N__14613),
            .in3(N__13049),
            .lcout(\this_vga_signals.if_m2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_1_LC_11_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_1_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_1_LC_11_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_1_LC_11_21_0  (
            .in0(N__13278),
            .in1(N__14351),
            .in2(N__14419),
            .in3(N__13038),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_LC_11_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_LC_11_21_1 .LUT_INIT=16'b0010110101001011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_LC_11_21_1  (
            .in0(N__13094),
            .in1(N__14475),
            .in2(N__12951),
            .in3(N__14410),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_ac0_3_0_LC_11_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_ac0_3_0_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_ac0_3_0_LC_11_21_2 .LUT_INIT=16'b1101001111000001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_ac0_3_0_LC_11_21_2  (
            .in0(N__14848),
            .in1(N__13152),
            .in2(N__14807),
            .in3(N__13112),
            .lcout(\this_vga_signals.mult1_un89_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_11_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_11_21_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_11_21_3  (
            .in0(N__13113),
            .in1(N__12948),
            .in2(N__13172),
            .in3(N__12936),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un89_sum_axbxc3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI6DOUP9_9_LC_11_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI6DOUP9_9_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI6DOUP9_9_LC_11_21_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI6DOUP9_9_LC_11_21_4  (
            .in0(N__17120),
            .in1(_gnd_net_),
            .in2(N__13206),
            .in3(N__13203),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axb1_LC_11_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axb1_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axb1_LC_11_21_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axb1_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__14607),
            .in2(_gnd_net_),
            .in3(N__13165),
            .lcout(\this_vga_signals.mult1_un82_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_11_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_11_21_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__13142),
            .in2(_gnd_net_),
            .in3(N__13124),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_11_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_11_22_0 .LUT_INIT=16'b1100111010001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_11_22_0  (
            .in0(N__13276),
            .in1(N__13064),
            .in2(N__14418),
            .in3(N__14349),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_11_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_11_22_3 .LUT_INIT=16'b1100000110000011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_11_22_3  (
            .in0(N__14350),
            .in1(N__14406),
            .in2(N__13068),
            .in3(N__13277),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_11_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_11_22_4 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_11_22_4  (
            .in0(N__14225),
            .in1(N__14170),
            .in2(N__14291),
            .in3(N__14346),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9 ),
            .ltout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_1_LC_11_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_1_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_1_LC_11_22_5 .LUT_INIT=16'b0101010110101110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_1_LC_11_22_5  (
            .in0(N__14348),
            .in1(N__14401),
            .in2(N__13074),
            .in3(N__13275),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_11_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_11_22_6 .LUT_INIT=16'b0111101000011010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_11_22_6  (
            .in0(N__14402),
            .in1(N__14454),
            .in2(N__13071),
            .in3(N__13063),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_11_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_11_22_7 .LUT_INIT=16'b1100000101111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_11_22_7  (
            .in0(N__14347),
            .in1(N__14274),
            .in2(N__14181),
            .in3(N__14224),
            .lcout(\this_vga_signals.SUM_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_LC_11_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_11_23_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_11_23_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(N__13259),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_pcounter_q_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32623),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_RNIC95C3_LC_11_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIC95C3_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIC95C3_LC_11_23_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_RNIC95C3_LC_11_23_4  (
            .in0(N__13745),
            .in1(N__13728),
            .in2(_gnd_net_),
            .in3(N__21661),
            .lcout(\this_vga_signals.M_pcounter_q_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI3O9R_1_LC_11_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI3O9R_1_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI3O9R_1_LC_11_23_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI3O9R_1_LC_11_23_5  (
            .in0(N__14806),
            .in1(N__14618),
            .in2(_gnd_net_),
            .in3(N__14548),
            .lcout(\this_vga_signals.N_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_1_LC_11_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_1_LC_11_23_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_1_LC_11_23_7 .LUT_INIT=16'b0000010011110000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_1_LC_11_23_7  (
            .in0(N__21662),
            .in1(N__13709),
            .in2(N__13734),
            .in3(N__21525),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32623),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI9JJM1_0_LC_11_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI9JJM1_0_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI9JJM1_0_LC_11_24_1 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI9JJM1_0_LC_11_24_1  (
            .in0(N__13241),
            .in1(N__14476),
            .in2(N__14853),
            .in3(N__14420),
            .lcout(\this_vga_signals.M_hcounter_q_RNI9JJM1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_5_LC_11_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_5_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_5_LC_11_24_3 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIADGD1_5_LC_11_24_3  (
            .in0(N__13242),
            .in1(N__14477),
            .in2(_gnd_net_),
            .in3(N__14421),
            .lcout(),
            .ltout(\this_vga_signals.M_hcounter_q_RNIADGD1Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIOC7D3_6_LC_11_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIOC7D3_6_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIOC7D3_6_LC_11_24_4 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIOC7D3_6_LC_11_24_4  (
            .in0(N__14363),
            .in1(N__13233),
            .in2(N__13227),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.i5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_11_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_11_24_7 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_11_24_7  (
            .in0(N__14247),
            .in1(_gnd_net_),
            .in2(N__14196),
            .in3(N__14305),
            .lcout(this_vga_signals_hvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_11_25_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_11_25_2 .LUT_INIT=16'b1101010111010111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_11_25_2  (
            .in0(N__14245),
            .in1(N__14191),
            .in2(N__14309),
            .in3(N__14364),
            .lcout(\this_vga_signals.SUM_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIML464_9_LC_11_25_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIML464_9_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIML464_9_LC_11_25_5 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIML464_9_LC_11_25_5  (
            .in0(N__14192),
            .in1(N__13449),
            .in2(N__14310),
            .in3(N__14246),
            .lcout(this_vga_signals_hsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNI1DAA_7_LC_11_25_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNI1DAA_7_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNI1DAA_7_LC_11_25_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_vaddress_q_RNI1DAA_7_LC_11_25_7  (
            .in0(_gnd_net_),
            .in1(N__16158),
            .in2(_gnd_net_),
            .in3(N__16205),
            .lcout(M_this_ppu_map_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI9E7F1_LC_11_26_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI9E7F1_LC_11_26_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI9E7F1_LC_11_26_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI9E7F1_LC_11_26_2  (
            .in0(N__24507),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19892),
            .lcout(N_63_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIMF36L_9_LC_11_26_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIMF36L_9_LC_11_26_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIMF36L_9_LC_11_26_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIMF36L_9_LC_11_26_4  (
            .in0(N__17079),
            .in1(N__13398),
            .in2(_gnd_net_),
            .in3(N__13368),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHL0E5_9_LC_11_26_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHL0E5_9_LC_11_26_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHL0E5_9_LC_11_26_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIHL0E5_9_LC_11_26_5  (
            .in0(_gnd_net_),
            .in1(N__13329),
            .in2(_gnd_net_),
            .in3(N__17078),
            .lcout(M_this_vga_signals_address_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_29_LC_12_15_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_29_LC_12_15_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_29_LC_12_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_29_LC_12_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24502),
            .lcout(M_this_data_tmp_qZ0Z_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32541),
            .ce(N__17663),
            .sr(N__26066));
    defparam M_this_data_tmp_q_esr_5_LC_12_16_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_5_LC_12_16_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_5_LC_12_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_5_LC_12_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24490),
            .lcout(M_this_data_tmp_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32550),
            .ce(N__16520),
            .sr(N__26063));
    defparam M_this_data_tmp_q_esr_12_LC_12_17_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_12_LC_12_17_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_12_LC_12_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_12_LC_12_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28324),
            .lcout(M_this_data_tmp_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32562),
            .ce(N__17352),
            .sr(N__26060));
    defparam M_this_data_tmp_q_esr_13_LC_12_17_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_13_LC_12_17_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_13_LC_12_17_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_13_LC_12_17_3 (
            .in0(N__24489),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32562),
            .ce(N__17352),
            .sr(N__26060));
    defparam M_this_data_tmp_q_esr_9_LC_12_17_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_9_LC_12_17_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_9_LC_12_17_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_9_LC_12_17_6 (
            .in0(N__30929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32562),
            .ce(N__17352),
            .sr(N__26060));
    defparam M_this_data_tmp_q_esr_0_LC_12_18_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_0_LC_12_18_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_0_LC_12_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_0_LC_12_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28447),
            .lcout(M_this_data_tmp_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32571),
            .ce(N__16512),
            .sr(N__26056));
    defparam \this_ppu.M_haddress_q_5_LC_12_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_5_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_5_LC_12_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_haddress_q_5_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__13558),
            .in2(_gnd_net_),
            .in3(N__13457),
            .lcout(M_this_ppu_map_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32581),
            .ce(),
            .sr(N__14922));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_12_19_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_12_19_1 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_12_19_1  (
            .in0(N__28527),
            .in1(N__26991),
            .in2(N__28677),
            .in3(N__28626),
            .lcout(M_this_ppu_vram_data_0),
            .ltout(M_this_ppu_vram_data_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.vram_en_i_a2_0_LC_12_19_2 .C_ON=1'b0;
    defparam \this_ppu.vram_en_i_a2_0_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.vram_en_i_a2_0_LC_12_19_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.vram_en_i_a2_0_LC_12_19_2  (
            .in0(N__28783),
            .in1(N__17182),
            .in2(N__13467),
            .in3(N__21160),
            .lcout(\this_ppu.N_134 ),
            .ltout(\this_ppu.N_134_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIUTM1G_5_LC_12_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIUTM1G_5_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIUTM1G_5_LC_12_19_3 .LUT_INIT=16'b1100111111001100;
    LogicCell40 \this_ppu.M_state_q_RNIUTM1G_5_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__14640),
            .in2(N__13464),
            .in3(N__32123),
            .lcout(M_this_ppu_vram_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_6_LC_12_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_6_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_6_LC_12_19_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_haddress_q_6_LC_12_19_4  (
            .in0(N__13559),
            .in1(N__13606),
            .in2(_gnd_net_),
            .in3(N__13458),
            .lcout(M_this_ppu_vram_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32581),
            .ce(),
            .sr(N__14922));
    defparam \this_ppu.M_haddress_q_RNINDU1G_1_LC_12_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNINDU1G_1_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNINDU1G_1_LC_12_19_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNINDU1G_1_LC_12_19_5  (
            .in0(N__20910),
            .in1(N__19285),
            .in2(_gnd_net_),
            .in3(N__13995),
            .lcout(\this_ppu.un1_M_haddress_q_c2 ),
            .ltout(\this_ppu.un1_M_haddress_q_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI4T92G_4_LC_12_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI4T92G_4_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI4T92G_4_LC_12_19_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNI4T92G_4_LC_12_19_6  (
            .in0(N__13796),
            .in1(N__13927),
            .in2(N__13461),
            .in3(N__13873),
            .lcout(\this_ppu.un1_M_haddress_q_c5 ),
            .ltout(\this_ppu.un1_M_haddress_q_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_7_LC_12_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_7_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_7_LC_12_19_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \this_ppu.M_haddress_q_7_LC_12_19_7  (
            .in0(N__13607),
            .in1(N__13560),
            .in2(N__13530),
            .in3(N__13527),
            .lcout(\this_ppu.M_haddress_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32581),
            .ce(),
            .sr(N__14922));
    defparam \this_ppu.M_state_q_1_LC_12_20_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_1_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_1_LC_12_20_1 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \this_ppu.M_state_q_1_LC_12_20_1  (
            .in0(N__32140),
            .in1(N__13977),
            .in2(N__14694),
            .in3(N__13758),
            .lcout(\this_ppu.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32590),
            .ce(),
            .sr(N__26051));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_21_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__14849),
            .in2(N__14808),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_21_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_21_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_21_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_12_21_1  (
            .in0(N__21491),
            .in1(N__14617),
            .in2(_gnd_net_),
            .in3(N__13515),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__32598),
            .ce(),
            .sr(N__14750));
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_21_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_21_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_21_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_12_21_2  (
            .in0(N__21488),
            .in1(N__14528),
            .in2(_gnd_net_),
            .in3(N__13512),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__32598),
            .ce(),
            .sr(N__14750));
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_21_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_21_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_21_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_12_21_3  (
            .in0(N__21492),
            .in1(N__14474),
            .in2(_gnd_net_),
            .in3(N__13509),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__32598),
            .ce(),
            .sr(N__14750));
    defparam \this_vga_signals.M_hcounter_q_5_LC_12_21_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_12_21_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_12_21_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_12_21_4  (
            .in0(N__21489),
            .in1(N__14412),
            .in2(_gnd_net_),
            .in3(N__13506),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__32598),
            .ce(),
            .sr(N__14750));
    defparam \this_vga_signals.M_hcounter_q_6_LC_12_21_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_12_21_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_12_21_5  (
            .in0(N__21493),
            .in1(N__14359),
            .in2(_gnd_net_),
            .in3(N__13503),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__32598),
            .ce(),
            .sr(N__14750));
    defparam \this_vga_signals.M_hcounter_q_7_LC_12_21_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_12_21_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_12_21_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_12_21_6  (
            .in0(N__21490),
            .in1(N__14180),
            .in2(_gnd_net_),
            .in3(N__13500),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__32598),
            .ce(),
            .sr(N__14750));
    defparam \this_vga_signals.M_hcounter_q_8_LC_12_21_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_12_21_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_12_21_7  (
            .in0(N__21494),
            .in1(N__14235),
            .in2(_gnd_net_),
            .in3(N__13752),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__32598),
            .ce(),
            .sr(N__14750));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_12_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_12_22_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_12_22_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__14290),
            .in2(_gnd_net_),
            .in3(N__13749),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32607),
            .ce(N__14862),
            .sr(N__14749));
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_12_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_12_23_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_12_23_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_0_LC_12_23_0  (
            .in0(N__13746),
            .in1(N__13733),
            .in2(_gnd_net_),
            .in3(N__21638),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32617),
            .ce(N__21524),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI7C7F1_LC_12_24_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI7C7F1_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI7C7F1_LC_12_24_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI7C7F1_LC_12_24_5  (
            .in0(_gnd_net_),
            .in1(N__31330),
            .in2(_gnd_net_),
            .in3(N__19876),
            .lcout(N_815_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIE00C4_9_LC_12_26_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIE00C4_9_LC_12_26_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIE00C4_9_LC_12_26_6 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIE00C4_9_LC_12_26_6  (
            .in0(N__14292),
            .in1(N__14236),
            .in2(N__15865),
            .in3(N__14182),
            .lcout(M_this_vga_ramdac_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI8D7F1_LC_12_27_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI8D7F1_LC_12_27_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI8D7F1_LC_12_27_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI8D7F1_LC_12_27_1  (
            .in0(N__28245),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19823),
            .lcout(N_814_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNI0655_6_LC_12_27_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNI0655_6_LC_12_27_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNI0655_6_LC_12_27_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.M_vaddress_q_RNI0655_6_LC_12_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16206),
            .lcout(this_ppu_M_vaddress_q_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_1_LC_13_16_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_1_LC_13_16_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_1_LC_13_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_1_LC_13_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30846),
            .lcout(M_this_data_tmp_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32542),
            .ce(N__16516),
            .sr(N__26061));
    defparam M_this_data_tmp_q_esr_24_LC_13_17_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_24_LC_13_17_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_24_LC_13_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_24_LC_13_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28454),
            .lcout(M_this_data_tmp_qZ0Z_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32551),
            .ce(N__17649),
            .sr(N__26057));
    defparam M_this_data_tmp_q_esr_6_LC_13_18_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_6_LC_13_18_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_6_LC_13_18_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_6_LC_13_18_1 (
            .in0(N__28148),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32563),
            .ce(N__16499),
            .sr(N__26054));
    defparam \this_ppu.M_haddress_q_RNIEV7R_2_LC_13_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIEV7R_2_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIEV7R_2_LC_13_19_0 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_ppu.M_haddress_q_RNIEV7R_2_LC_13_19_0  (
            .in0(N__32134),
            .in1(N__13863),
            .in2(N__31935),
            .in3(N__14130),
            .lcout(M_this_ppu_sprites_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_2_LC_13_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_2_LC_13_19_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_2_LC_13_19_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_haddress_q_2_LC_13_19_1  (
            .in0(N__13997),
            .in1(N__13865),
            .in2(N__19307),
            .in3(N__20912),
            .lcout(M_this_ppu_vram_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32572),
            .ce(),
            .sr(N__14918));
    defparam \this_ppu.M_haddress_q_RNO_0_3_LC_13_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNO_0_3_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNO_0_3_LC_13_19_2 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \this_ppu.M_haddress_q_RNO_0_3_LC_13_19_2  (
            .in0(N__32133),
            .in1(N__19286),
            .in2(N__14649),
            .in3(N__13975),
            .lcout(),
            .ltout(\this_ppu.un1_M_haddress_q_c1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_3_LC_13_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_3_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_3_LC_13_19_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \this_ppu.M_haddress_q_3_LC_13_19_3  (
            .in0(N__13928),
            .in1(N__13866),
            .in2(N__14013),
            .in3(N__20913),
            .lcout(M_this_ppu_map_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32572),
            .ce(),
            .sr(N__14918));
    defparam \this_ppu.M_haddress_q_1_LC_13_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_1_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_1_LC_13_19_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_haddress_q_1_LC_13_19_4  (
            .in0(N__20911),
            .in1(N__19290),
            .in2(_gnd_net_),
            .in3(N__13996),
            .lcout(M_this_ppu_vram_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32572),
            .ce(),
            .sr(N__14918));
    defparam \this_ppu.M_haddress_q_0_LC_13_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_0_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_0_LC_13_19_5 .LUT_INIT=16'b0010110100111100;
    LogicCell40 \this_ppu.M_haddress_q_0_LC_13_19_5  (
            .in0(N__13976),
            .in1(N__14647),
            .in2(N__19306),
            .in3(N__32135),
            .lcout(M_this_ppu_vram_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32572),
            .ce(),
            .sr(N__14918));
    defparam \this_ppu.M_haddress_q_4_LC_13_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_4_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_4_LC_13_19_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_haddress_q_4_LC_13_19_6  (
            .in0(N__13929),
            .in1(N__13864),
            .in2(N__13797),
            .in3(N__13833),
            .lcout(M_this_ppu_map_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32572),
            .ce(),
            .sr(N__14918));
    defparam \this_ppu.M_state_q_RNO_1_1_LC_13_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_1_1_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_1_1_LC_13_20_2 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \this_ppu.M_state_q_RNO_1_1_LC_13_20_2  (
            .in0(N__16982),
            .in1(N__32132),
            .in2(N__14648),
            .in3(N__16917),
            .lcout(\this_ppu.N_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_1_LC_13_20_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_13_20_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.M_state_q_RNO_0_1_LC_13_20_4  (
            .in0(N__14657),
            .in1(N__31883),
            .in2(_gnd_net_),
            .in3(N__17459),
            .lcout(\this_ppu.M_state_qc_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_4_LC_13_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_4_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_4_LC_13_20_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_state_q_RNO_0_4_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__14672),
            .in2(_gnd_net_),
            .in3(N__28791),
            .lcout(),
            .ltout(\this_ppu.M_state_qc_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_4_LC_13_20_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_4_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_4_LC_13_20_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_ppu.M_state_q_4_LC_13_20_6  (
            .in0(N__32136),
            .in1(N__17189),
            .in2(N__14661),
            .in3(N__21161),
            .lcout(\this_ppu.M_state_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32582),
            .ce(),
            .sr(N__26048));
    defparam \this_ppu.M_state_q_5_LC_13_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_5_LC_13_20_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_5_LC_13_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.M_state_q_5_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14658),
            .lcout(\this_ppu.M_state_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32582),
            .ce(),
            .sr(N__26048));
    defparam \this_start_data_delay.G_464_LC_13_21_4 .C_ON=1'b0;
    defparam \this_start_data_delay.G_464_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.G_464_LC_13_21_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.G_464_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(N__21478),
            .in2(_gnd_net_),
            .in3(N__21637),
            .lcout(G_464),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_13_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_13_22_1 .LUT_INIT=16'b0001111111111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_13_22_1  (
            .in0(N__14772),
            .in1(N__14828),
            .in2(N__14611),
            .in3(N__14521),
            .lcout(),
            .ltout(\this_vga_signals.N_18_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_5_LC_13_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_5_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_5_LC_13_22_2 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIEVMV1_5_LC_13_22_2  (
            .in0(N__14472),
            .in1(N__14411),
            .in2(N__14367),
            .in3(N__14352),
            .lcout(),
            .ltout(\this_vga_signals.m23_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_13_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_13_22_3 .LUT_INIT=16'b1000100000001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_13_22_3  (
            .in0(N__14278),
            .in1(N__14226),
            .in2(N__14199),
            .in3(N__14171),
            .lcout(this_vga_signals_M_hcounter_d7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_22_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_22_7  (
            .in0(N__21521),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14742),
            .lcout(\this_vga_signals.N_1090_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_0_LC_13_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_13_23_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_13_23_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_13_23_2  (
            .in0(N__21522),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14838),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32608),
            .ce(),
            .sr(N__14751));
    defparam \this_vga_signals.M_hcounter_q_1_LC_13_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_13_23_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_13_23_3 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_13_23_3  (
            .in0(N__14837),
            .in1(N__21523),
            .in2(_gnd_net_),
            .in3(N__14783),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32608),
            .ce(),
            .sr(N__14751));
    defparam \this_reset_cond.M_stage_q_1_LC_14_15_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_14_15_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_14_15_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__16303),
            .in2(_gnd_net_),
            .in3(N__14997),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32534),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_14_15_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_14_15_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_14_15_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__16304),
            .in2(_gnd_net_),
            .in3(N__14721),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32534),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_14_16_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_14_16_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_14_16_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_14_16_1  (
            .in0(N__16302),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14715),
            .lcout(\this_reset_cond.M_stage_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32537),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_0_LC_14_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_0_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_0_LC_14_17_3 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \this_ppu.M_count_q_0_LC_14_17_3  (
            .in0(N__15357),
            .in1(N__15171),
            .in2(_gnd_net_),
            .in3(N__15120),
            .lcout(\this_ppu.M_count_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32543),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_oam_ram_write_data_10_LC_14_17_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_10_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_oam_ram_write_data_10_LC_14_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_this_oam_ram_write_data_10_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__15402),
            .in2(_gnd_net_),
            .in3(N__18527),
            .lcout(M_this_oam_ram_write_data_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_14_18_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_14_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__15356),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\this_ppu.un1_M_count_q_1_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_14_18_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_14_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__14937),
            .in2(N__29676),
            .in3(N__14697),
            .lcout(\this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_0_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_14_18_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_14_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__29569),
            .in2(N__15330),
            .in3(N__14892),
            .lcout(\this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_1_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_14_18_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_14_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__15374),
            .in2(N__29677),
            .in3(N__14889),
            .lcout(\this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_2_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_14_18_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_14_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__29573),
            .in2(N__14955),
            .in3(N__14886),
            .lcout(\this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_3_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_14_18_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_14_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__14972),
            .in2(N__29678),
            .in3(N__14883),
            .lcout(\this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_4_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_14_18_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_14_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__29577),
            .in2(N__15087),
            .in3(N__14880),
            .lcout(\this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_5_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_7_LC_14_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_14_18_7 .LUT_INIT=16'b1100110000110110;
    LogicCell40 \this_ppu.M_count_q_RNO_0_7_LC_14_18_7  (
            .in0(N__17467),
            .in1(N__15434),
            .in2(N__16887),
            .in3(N__14877),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIKRC91_1_LC_14_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIKRC91_1_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIKRC91_1_LC_14_19_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_state_q_RNIKRC91_1_LC_14_19_0  (
            .in0(N__17466),
            .in1(N__17420),
            .in2(_gnd_net_),
            .in3(N__17402),
            .lcout(\this_ppu.M_state_d_0_sqmuxa_1 ),
            .ltout(\this_ppu.M_state_d_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI2UC86_1_LC_14_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI2UC86_1_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI2UC86_1_LC_14_19_1 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \this_ppu.M_state_q_RNI2UC86_1_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__15773),
            .in2(N__14874),
            .in3(N__16876),
            .lcout(\this_ppu.N_1456_0 ),
            .ltout(\this_ppu.N_1456_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_4_LC_14_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_4_LC_14_19_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_4_LC_14_19_2 .LUT_INIT=16'b1110000000010000;
    LogicCell40 \this_ppu.M_count_q_4_LC_14_19_2  (
            .in0(N__15161),
            .in1(N__14871),
            .in2(N__14865),
            .in3(N__14951),
            .lcout(\this_ppu.M_count_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32564),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_5_LC_14_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_5_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_5_LC_14_19_4 .LUT_INIT=16'b1010100000000010;
    LogicCell40 \this_ppu.M_count_q_5_LC_14_19_4  (
            .in0(N__15116),
            .in1(N__14991),
            .in2(N__15172),
            .in3(N__14973),
            .lcout(\this_ppu.M_count_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32564),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_1_LC_14_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_1_LC_14_19_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_1_LC_14_19_5 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_1_LC_14_19_5  (
            .in0(N__14936),
            .in1(N__15160),
            .in2(N__14985),
            .in3(N__15115),
            .lcout(\this_ppu.M_count_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32564),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNICD0G_1_LC_14_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNICD0G_1_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNICD0G_1_LC_14_19_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_count_q_RNICD0G_1_LC_14_19_6  (
            .in0(N__14971),
            .in1(N__14950),
            .in2(N__15086),
            .in3(N__14935),
            .lcout(\this_ppu.M_state_q_srsts_i_a3_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIE20V4_0_LC_14_20_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIE20V4_0_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIE20V4_0_LC_14_20_0 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \this_ppu.M_state_q_RNIE20V4_0_LC_14_20_0  (
            .in0(N__16974),
            .in1(N__15772),
            .in2(N__16922),
            .in3(N__16944),
            .lcout(\this_ppu.M_state_q_RNIE20V4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNIAUKV3_0_LC_14_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNIAUKV3_0_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNIAUKV3_0_LC_14_20_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNIAUKV3_0_LC_14_20_1  (
            .in0(N__15030),
            .in1(N__15051),
            .in2(_gnd_net_),
            .in3(N__15902),
            .lcout(M_this_vga_signals_line_clk_0),
            .ltout(M_this_vga_signals_line_clk_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI2TJN4_0_LC_14_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI2TJN4_0_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI2TJN4_0_LC_14_20_2 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \this_ppu.M_state_q_RNI2TJN4_0_LC_14_20_2  (
            .in0(N__16972),
            .in1(_gnd_net_),
            .in2(N__14901),
            .in3(N__16943),
            .lcout(\this_ppu.M_state_d_0_sqmuxa ),
            .ltout(\this_ppu.M_state_d_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIJV275_2_LC_14_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIJV275_2_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIJV275_2_LC_14_20_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIJV275_2_LC_14_20_3  (
            .in0(N__30281),
            .in1(N__16833),
            .in2(N__14898),
            .in3(N__32177),
            .lcout(\this_ppu.un1_M_vaddress_q_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_14_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_14_20_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_0_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__15031),
            .in2(_gnd_net_),
            .in3(N__15932),
            .lcout(),
            .ltout(\this_vga_signals.N_1000_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_0_LC_14_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_0_LC_14_20_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_0_LC_14_20_5 .LUT_INIT=16'b0111010011001100;
    LogicCell40 \this_vga_signals.M_lcounter_q_0_LC_14_20_5  (
            .in0(N__21660),
            .in1(N__15052),
            .in2(N__14895),
            .in3(N__21536),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32573),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI22015_0_LC_14_20_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI22015_0_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI22015_0_LC_14_20_6 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \this_ppu.M_state_q_RNI22015_0_LC_14_20_6  (
            .in0(N__16973),
            .in1(N__16945),
            .in2(N__17468),
            .in3(N__16916),
            .lcout(\this_ppu.un10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_4_LC_14_21_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_4_LC_14_21_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_4_LC_14_21_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_4_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__16280),
            .in2(_gnd_net_),
            .in3(N__15063),
            .lcout(\this_reset_cond.M_stage_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32583),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_LC_14_21_1 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_LC_14_21_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.line_clk.M_last_q_LC_14_21_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_LC_14_21_1  (
            .in0(N__15054),
            .in1(N__15032),
            .in2(_gnd_net_),
            .in3(N__15903),
            .lcout(\this_ppu.M_last_q ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32583),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIE6DH5_4_LC_14_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIE6DH5_4_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIE6DH5_4_LC_14_21_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIE6DH5_4_LC_14_21_5  (
            .in0(N__16625),
            .in1(N__16691),
            .in2(_gnd_net_),
            .in3(N__16712),
            .lcout(\this_ppu.un1_M_vaddress_q_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_14_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_14_21_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_1_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__15053),
            .in2(_gnd_net_),
            .in3(N__15933),
            .lcout(),
            .ltout(\this_vga_signals.i21_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_1_LC_14_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_1_LC_14_21_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_1_LC_14_21_7 .LUT_INIT=16'b0110001011101010;
    LogicCell40 \this_vga_signals.M_lcounter_q_1_LC_14_21_7  (
            .in0(N__15033),
            .in1(N__21495),
            .in2(N__15036),
            .in3(N__21639),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32583),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGB2A6_6_LC_14_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGB2A6_6_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGB2A6_6_LC_14_22_0 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGB2A6_6_LC_14_22_0  (
            .in0(N__21622),
            .in1(N__15408),
            .in2(_gnd_net_),
            .in3(N__22400),
            .lcout(\this_vga_signals.N_129_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_6_LC_14_24_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_6_LC_14_24_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_6_LC_14_24_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_vaddress_q_6_LC_14_24_4  (
            .in0(N__16197),
            .in1(N__16775),
            .in2(_gnd_net_),
            .in3(N__16175),
            .lcout(\this_ppu.M_vaddress_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32609),
            .ce(),
            .sr(N__16584));
    defparam \this_start_data_delay.M_last_q_RNI5A7F1_LC_14_25_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI5A7F1_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI5A7F1_LC_14_25_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI5A7F1_LC_14_25_1  (
            .in0(N__30863),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19872),
            .lcout(N_817_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_15_14_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_15_14_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_15_14_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_15_14_4  (
            .in0(N__16293),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32531),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_10_LC_15_16_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_10_LC_15_16_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_10_LC_15_16_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_10_LC_15_16_2 (
            .in0(N__32826),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32535),
            .ce(N__17339),
            .sr(N__26055));
    defparam M_this_data_tmp_q_esr_17_LC_15_17_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_17_LC_15_17_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_17_LC_15_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_17_LC_15_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30913),
            .lcout(M_this_data_tmp_qZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32538),
            .ce(N__15947),
            .sr(N__26052));
    defparam \this_ppu.M_count_q_3_LC_15_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_3_LC_15_18_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_3_LC_15_18_0 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_3_LC_15_18_0  (
            .in0(N__15375),
            .in1(N__15174),
            .in2(N__15384),
            .in3(N__15119),
            .lcout(\this_ppu.M_count_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32544),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNI890G_7_LC_15_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNI890G_7_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNI890G_7_LC_15_18_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_count_q_RNI890G_7_LC_15_18_1  (
            .in0(N__15373),
            .in1(N__15325),
            .in2(N__15435),
            .in3(N__15355),
            .lcout(\this_ppu.M_state_q_srsts_i_a3_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_2_LC_15_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_2_LC_15_18_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_2_LC_15_18_4 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_2_LC_15_18_4  (
            .in0(N__15326),
            .in1(N__15173),
            .in2(N__15339),
            .in3(N__15118),
            .lcout(\this_ppu.M_count_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32544),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIMGCA_0_LC_15_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIMGCA_0_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIMGCA_0_LC_15_19_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_ppu.M_vaddress_q_RNIMGCA_0_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__16820),
            .in2(_gnd_net_),
            .in3(N__16449),
            .lcout(),
            .ltout(\this_ppu.un10_sprites_addr_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIMQ241_2_LC_15_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIMQ241_2_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIMQ241_2_LC_15_19_2 .LUT_INIT=16'b0000111101001110;
    LogicCell40 \this_ppu.M_state_q_RNIMQ241_2_LC_15_19_2  (
            .in0(N__31884),
            .in1(N__15312),
            .in2(N__15294),
            .in3(N__32076),
            .lcout(M_this_ppu_sprites_addr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_6_LC_15_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_6_LC_15_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_6_LC_15_19_3 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_6_LC_15_19_3  (
            .in0(N__15085),
            .in1(N__15165),
            .in2(N__15132),
            .in3(N__15117),
            .lcout(\this_ppu.M_count_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32552),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIS8A01_0_LC_15_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIS8A01_0_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIS8A01_0_LC_15_19_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \this_ppu.M_vaddress_q_RNIS8A01_0_LC_15_19_4  (
            .in0(N__16821),
            .in1(N__32078),
            .in2(N__31912),
            .in3(N__15726),
            .lcout(M_this_ppu_sprites_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_15_19_5 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_15_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_0_RNISG75_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15606),
            .lcout(M_this_oam_ram_read_data_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIMTR41_2_LC_15_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIMTR41_2_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIMTR41_2_LC_15_19_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \this_ppu.M_state_q_RNIMTR41_2_LC_15_19_7  (
            .in0(N__32077),
            .in1(N__31885),
            .in2(N__15591),
            .in3(N__16416),
            .lcout(M_this_ppu_sprites_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.dmalto4_0_o2_LC_15_20_1 .C_ON=1'b0;
    defparam \this_start_data_delay.dmalto4_0_o2_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.dmalto4_0_o2_LC_15_20_1 .LUT_INIT=16'b1111001110100010;
    LogicCell40 \this_start_data_delay.dmalto4_0_o2_LC_15_20_1  (
            .in0(N__17775),
            .in1(N__19046),
            .in2(N__24318),
            .in3(N__22178),
            .lcout(\this_start_data_delay.N_43_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIELANC_0_LC_15_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIELANC_0_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIELANC_0_LC_15_20_3 .LUT_INIT=16'b1011111110101010;
    LogicCell40 \this_ppu.M_state_q_RNIELANC_0_LC_15_20_3  (
            .in0(N__15771),
            .in1(N__15850),
            .in2(N__17724),
            .in3(N__16871),
            .lcout(\this_ppu.M_state_q_RNIELANCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_0_LC_15_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_0_LC_15_20_5 .SEQ_MODE=4'b1001;
    defparam \this_ppu.M_state_q_0_LC_15_20_5 .LUT_INIT=16'b1111100011111100;
    LogicCell40 \this_ppu.M_state_q_0_LC_15_20_5  (
            .in0(N__16978),
            .in1(N__16946),
            .in2(N__15456),
            .in3(N__16921),
            .lcout(\this_ppu.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32565),
            .ce(),
            .sr(N__26045));
    defparam \this_ppu.M_count_q_7_LC_15_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_7_LC_15_20_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_7_LC_15_20_7 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \this_ppu.M_count_q_7_LC_15_20_7  (
            .in0(N__15452),
            .in1(N__15444),
            .in2(_gnd_net_),
            .in3(N__16872),
            .lcout(\this_ppu.M_count_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32565),
            .ce(),
            .sr(N__26045));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI4KCU6_9_LC_15_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI4KCU6_9_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI4KCU6_9_LC_15_21_0 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI4KCU6_9_LC_15_21_0  (
            .in0(N__22580),
            .in1(_gnd_net_),
            .in2(N__15417),
            .in3(N__21476),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNI4KCU6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI8O063_8_LC_15_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI8O063_8_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI8O063_8_LC_15_21_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI8O063_8_LC_15_21_2  (
            .in0(N__21990),
            .in1(N__23091),
            .in2(N__15918),
            .in3(N__21893),
            .lcout(\this_vga_signals.N_1028 ),
            .ltout(\this_vga_signals.N_1028_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFPFL6_9_LC_15_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFPFL6_9_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFPFL6_9_LC_15_21_3 .LUT_INIT=16'b0100000011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIFPFL6_9_LC_15_21_3  (
            .in0(N__22403),
            .in1(N__21670),
            .in2(N__15936),
            .in3(N__22581),
            .lcout(\this_vga_signals.N_999 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_15_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_15_21_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__22929),
            .in2(_gnd_net_),
            .in3(N__21579),
            .lcout(),
            .ltout(\this_vga_signals.N_1004_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIILO32_LC_15_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIILO32_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIILO32_LC_15_21_5 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIILO32_LC_15_21_5  (
            .in0(N__22859),
            .in1(N__22704),
            .in2(N__15921),
            .in3(N__20518),
            .lcout(\this_vga_signals.N_1013 ),
            .ltout(\this_vga_signals.N_1013_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9AJQ2_5_LC_15_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9AJQ2_5_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9AJQ2_5_LC_15_21_6 .LUT_INIT=16'b0101000101010001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI9AJQ2_5_LC_15_21_6  (
            .in0(N__22401),
            .in1(N__23090),
            .in2(N__15909),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\this_vga_signals.N_105_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3HRS3_8_LC_15_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3HRS3_8_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3HRS3_8_LC_15_21_7 .LUT_INIT=16'b0000000011100111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI3HRS3_8_LC_15_21_7  (
            .in0(N__21892),
            .in1(N__21989),
            .in2(N__15906),
            .in3(N__22579),
            .lcout(\this_vga_signals.N_113_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_6_LC_15_22_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_6_LC_15_22_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_6_LC_15_22_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_6_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__16317),
            .in2(_gnd_net_),
            .in3(N__15885),
            .lcout(\this_reset_cond.M_stage_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32584),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_5_LC_15_22_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_5_LC_15_22_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_5_LC_15_22_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_5_LC_15_22_1  (
            .in0(N__16316),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15891),
            .lcout(\this_reset_cond.M_stage_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32584),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_9_LC_15_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_9_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_9_LC_15_22_2 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_9_LC_15_22_2  (
            .in0(N__17025),
            .in1(N__20255),
            .in2(N__16215),
            .in3(N__22584),
            .lcout(this_vga_signals_vvisibility),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_9_LC_15_22_5 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_9_LC_15_22_5 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_9_LC_15_22_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_9_LC_15_22_5  (
            .in0(N__16320),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16221),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32584),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_7_LC_15_22_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_7_LC_15_22_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_7_LC_15_22_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_7_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__16318),
            .in2(_gnd_net_),
            .in3(N__16326),
            .lcout(\this_reset_cond.M_stage_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32584),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_8_LC_15_22_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_8_LC_15_22_7 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_8_LC_15_22_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_8_LC_15_22_7  (
            .in0(N__16319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16227),
            .lcout(\this_reset_cond.M_stage_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32584),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_8_LC_15_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_8_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_8_LC_15_23_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_8_LC_15_23_4  (
            .in0(N__21902),
            .in1(N__22000),
            .in2(N__22402),
            .in3(N__22583),
            .lcout(\this_vga_signals.vaddress_ac0_9_0_a0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_7_LC_15_24_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_7_LC_15_24_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_7_LC_15_24_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_vaddress_q_7_LC_15_24_6  (
            .in0(N__16198),
            .in1(N__16771),
            .in2(N__16157),
            .in3(N__16176),
            .lcout(\this_ppu.M_vaddress_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32599),
            .ce(),
            .sr(N__16583));
    defparam \this_ppu.M_state_q_3_LC_15_30_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_3_LC_15_30_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_3_LC_15_30_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.M_state_q_3_LC_15_30_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31965),
            .lcout(\this_ppu.M_state_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32640),
            .ce(),
            .sr(N__26044));
    defparam M_this_state_q_17_LC_16_15_0.C_ON=1'b0;
    defparam M_this_state_q_17_LC_16_15_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_17_LC_16_15_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 M_this_state_q_17_LC_16_15_0 (
            .in0(N__19404),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24243),
            .lcout(led23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32530),
            .ce(),
            .sr(N__26053));
    defparam dma_0_sbtinv_LC_16_16_6.C_ON=1'b0;
    defparam dma_0_sbtinv_LC_16_16_6.SEQ_MODE=4'b0000;
    defparam dma_0_sbtinv_LC_16_16_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 dma_0_sbtinv_LC_16_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17734),
            .lcout(dma_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI8G791_14_LC_16_17_3.C_ON=1'b0;
    defparam M_this_state_q_RNI8G791_14_LC_16_17_3.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI8G791_14_LC_16_17_3.LUT_INIT=16'b1110111010101010;
    LogicCell40 M_this_state_q_RNI8G791_14_LC_16_17_3 (
            .in0(N__26204),
            .in1(N__19119),
            .in2(_gnd_net_),
            .in3(N__24235),
            .lcout(N_1430_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.port_data_rw_0_a2_1_LC_16_17_7 .C_ON=1'b0;
    defparam \this_start_data_delay.port_data_rw_0_a2_1_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.port_data_rw_0_a2_1_LC_16_17_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_start_data_delay.port_data_rw_0_a2_1_LC_16_17_7  (
            .in0(N__31649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23913),
            .lcout(\this_start_data_delay.port_data_rw_0_a2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIUCR11_LC_16_18_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIUCR11_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIUCR11_LC_16_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIUCR11_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__19403),
            .in2(_gnd_net_),
            .in3(N__24242),
            .lcout(),
            .ltout(M_this_state_q_ns_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_RNIAI791_9_LC_16_18_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_RNIAI791_9_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \this_reset_cond.M_stage_q_RNIAI791_9_LC_16_18_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \this_reset_cond.M_stage_q_RNIAI791_9_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16524),
            .in3(N__26203),
            .lcout(M_this_state_q_ns_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_12_LC_16_18_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_12_LC_16_18_7 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_12_LC_16_18_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \this_sprites_ram.mem_radreg_12_LC_16_18_7  (
            .in0(N__31856),
            .in1(N__32142),
            .in2(N__16470),
            .in3(N__16353),
            .lcout(\this_sprites_ram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32536),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un10_sprites_addr_cry_0_c_inv_LC_16_19_0 .C_ON=1'b1;
    defparam \this_ppu.un10_sprites_addr_cry_0_c_inv_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un10_sprites_addr_cry_0_c_inv_LC_16_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un10_sprites_addr_cry_0_c_inv_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__16428),
            .in2(N__16832),
            .in3(N__16448),
            .lcout(\this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\this_ppu.un10_sprites_addr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5B_LC_16_19_1 .C_ON=1'b1;
    defparam \this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5B_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5B_LC_16_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5B_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__16422),
            .in2(N__32176),
            .in3(N__16410),
            .lcout(\this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5BZ0 ),
            .ltout(),
            .carryin(\this_ppu.un10_sprites_addr_cry_0 ),
            .carryout(\this_ppu.un10_sprites_addr_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un10_sprites_addr_cry_1_c_RNIOM6B_LC_16_19_2 .C_ON=1'b1;
    defparam \this_ppu.un10_sprites_addr_cry_1_c_RNIOM6B_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un10_sprites_addr_cry_1_c_RNIOM6B_LC_16_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un10_sprites_addr_cry_1_c_RNIOM6B_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__16407),
            .in2(N__30280),
            .in3(N__16392),
            .lcout(\this_ppu.un10_sprites_addr_cry_1_c_RNIOM6BZ0 ),
            .ltout(),
            .carryin(\this_ppu.un10_sprites_addr_cry_1 ),
            .carryout(\this_ppu.un10_sprites_addr_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un10_sprites_addr_cry_2_c_RNIQP7B_LC_16_19_3 .C_ON=1'b1;
    defparam \this_ppu.un10_sprites_addr_cry_2_c_RNIQP7B_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un10_sprites_addr_cry_2_c_RNIQP7B_LC_16_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un10_sprites_addr_cry_2_c_RNIQP7B_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__16389),
            .in2(N__16682),
            .in3(N__16374),
            .lcout(\this_ppu.un10_sprites_addr_cry_2_c_RNIQP7BZ0 ),
            .ltout(),
            .carryin(\this_ppu.un10_sprites_addr_cry_2 ),
            .carryout(\this_ppu.un10_sprites_addr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un10_sprites_addr_cry_3_c_RNISS8B_LC_16_19_4 .C_ON=1'b1;
    defparam \this_ppu.un10_sprites_addr_cry_3_c_RNISS8B_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un10_sprites_addr_cry_3_c_RNISS8B_LC_16_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un10_sprites_addr_cry_3_c_RNISS8B_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__16610),
            .in2(N__16371),
            .in3(N__16347),
            .lcout(\this_ppu.un10_sprites_addr_cry_3_c_RNISS8BZ0 ),
            .ltout(),
            .carryin(\this_ppu.un10_sprites_addr_cry_3 ),
            .carryout(\this_ppu.un10_sprites_addr_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un10_sprites_addr_cry_4_c_RNIUV9B_LC_16_19_5 .C_ON=1'b0;
    defparam \this_ppu.un10_sprites_addr_cry_4_c_RNIUV9B_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un10_sprites_addr_cry_4_c_RNIUV9B_LC_16_19_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_ppu.un10_sprites_addr_cry_4_c_RNIUV9B_LC_16_19_5  (
            .in0(N__16751),
            .in1(N__16344),
            .in2(_gnd_net_),
            .in3(N__16329),
            .lcout(\this_ppu.un10_sprites_addr_cry_4_c_RNIUV9BZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_0_LC_16_20_0 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_0_LC_16_20_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_0_LC_16_20_0 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \this_ppu.M_vaddress_q_0_LC_16_20_0  (
            .in0(N__16986),
            .in1(N__16947),
            .in2(N__16834),
            .in3(N__16923),
            .lcout(M_this_ppu_vram_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32548),
            .ce(),
            .sr(N__16582));
    defparam \this_ppu.M_vaddress_q_1_LC_16_20_1 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_1_LC_16_20_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_1_LC_16_20_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_vaddress_q_1_LC_16_20_1  (
            .in0(N__32174),
            .in1(N__16825),
            .in2(_gnd_net_),
            .in3(N__16886),
            .lcout(\this_ppu.M_vaddress_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32548),
            .ce(),
            .sr(N__16582));
    defparam \this_ppu.M_vaddress_q_2_LC_16_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_2_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_2_LC_16_20_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \this_ppu.M_vaddress_q_2_LC_16_20_2  (
            .in0(N__16885),
            .in1(N__32175),
            .in2(N__16835),
            .in3(N__30279),
            .lcout(\this_ppu.M_vaddress_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32548),
            .ce(),
            .sr(N__16582));
    defparam \this_ppu.M_vaddress_q_5_LC_16_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_5_LC_16_20_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_5_LC_16_20_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_vaddress_q_5_LC_16_20_3  (
            .in0(N__16722),
            .in1(N__16755),
            .in2(N__16687),
            .in3(N__16615),
            .lcout(M_this_ppu_map_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32548),
            .ce(),
            .sr(N__16582));
    defparam \this_ppu.M_vaddress_q_3_LC_16_20_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_3_LC_16_20_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_3_LC_16_20_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_vaddress_q_3_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__16672),
            .in2(_gnd_net_),
            .in3(N__16720),
            .lcout(M_this_ppu_map_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32548),
            .ce(),
            .sr(N__16582));
    defparam \this_ppu.M_vaddress_q_4_LC_16_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_4_LC_16_20_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_4_LC_16_20_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \this_ppu.M_vaddress_q_4_LC_16_20_5  (
            .in0(N__16721),
            .in1(_gnd_net_),
            .in2(N__16686),
            .in3(N__16614),
            .lcout(M_this_ppu_map_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32548),
            .ce(),
            .sr(N__16582));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIPE977_9_LC_16_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIPE977_9_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIPE977_9_LC_16_21_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIPE977_9_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(N__21477),
            .in2(_gnd_net_),
            .in3(N__16541),
            .lcout(\this_vga_signals.N_1090_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_16_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_16_22_0 .LUT_INIT=16'b0001101101110010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_LC_16_22_0  (
            .in0(N__17019),
            .in1(N__17673),
            .in2(N__17580),
            .in3(N__17562),
            .lcout(),
            .ltout(\this_vga_signals.g1_2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_16_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_16_22_1 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_LC_16_22_1  (
            .in0(N__17373),
            .in1(N__22935),
            .in2(N__16527),
            .in3(N__17007),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_c3_0_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI3KH3P1_1_LC_16_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI3KH3P1_1_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI3KH3P1_1_LC_16_22_2 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI3KH3P1_1_LC_16_22_2  (
            .in0(N__17130),
            .in1(N__17385),
            .in2(N__17049),
            .in3(N__17523),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_5_LC_16_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_5_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_5_LC_16_22_3 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICM2P1_5_LC_16_22_3  (
            .in0(N__23087),
            .in1(N__23248),
            .in2(N__22437),
            .in3(N__22386),
            .lcout(\this_vga_signals.un6_vvisibilitylt9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_LC_16_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_LC_16_22_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_LC_16_22_5  (
            .in0(N__16992),
            .in1(N__17967),
            .in2(N__18057),
            .in3(N__17571),
            .lcout(\this_vga_signals.g2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_8_LC_16_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_8_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_8_LC_16_23_0 .LUT_INIT=16'b1000101011100111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_8_LC_16_23_0  (
            .in0(N__21903),
            .in1(N__22001),
            .in2(N__20187),
            .in3(N__22582),
            .lcout(),
            .ltout(\this_vga_signals.SUM_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_16_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_16_23_1 .LUT_INIT=16'b1001011010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_13_LC_16_23_1  (
            .in0(N__22002),
            .in1(N__22391),
            .in2(N__17013),
            .in3(N__20256),
            .lcout(\this_vga_signals.g3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_2_LC_16_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_2_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_2_LC_16_23_3 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_2_LC_16_23_3  (
            .in0(N__22861),
            .in1(N__20286),
            .in2(N__23286),
            .in3(N__18260),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c2_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_16_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_16_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_8_LC_16_23_4  (
            .in0(N__18261),
            .in1(N__18702),
            .in2(N__17010),
            .in3(N__17586),
            .lcout(\this_vga_signals.N_4_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_a3_LC_16_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_a3_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_a3_LC_16_23_5 .LUT_INIT=16'b1111011111111101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_a3_LC_16_23_5  (
            .in0(N__23278),
            .in1(N__22392),
            .in2(N__23100),
            .in3(N__20424),
            .lcout(),
            .ltout(\this_vga_signals.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g4_LC_16_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g4_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g4_LC_16_23_6 .LUT_INIT=16'b1110110011111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g4_LC_16_23_6  (
            .in0(N__22393),
            .in1(N__17001),
            .in2(N__16995),
            .in3(N__18885),
            .lcout(\this_vga_signals.g4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI9H791_15_LC_17_16_6.C_ON=1'b0;
    defparam M_this_state_q_RNI9H791_15_LC_17_16_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI9H791_15_LC_17_16_6.LUT_INIT=16'b1110111010101010;
    LogicCell40 M_this_state_q_RNI9H791_15_LC_17_16_6 (
            .in0(N__26205),
            .in1(N__19146),
            .in2(_gnd_net_),
            .in3(N__24241),
            .lcout(N_1438_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.port_data_rw_0_i_LC_17_17_3 .C_ON=1'b0;
    defparam \this_start_data_delay.port_data_rw_0_i_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.port_data_rw_0_i_LC_17_17_3 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \this_start_data_delay.port_data_rw_0_i_LC_17_17_3  (
            .in0(N__23576),
            .in1(N__17304),
            .in2(N__18153),
            .in3(N__17766),
            .lcout(port_data_rw_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_17_18_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_17_18_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_17_18_0  (
            .in0(N__17274),
            .in1(N__17262),
            .in2(_gnd_net_),
            .in3(N__30108),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_17_18_4 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_17_18_4 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_17_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17250),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32545),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_17_19_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_17_19_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_17_19_1  (
            .in0(N__30100),
            .in1(N__17232),
            .in2(_gnd_net_),
            .in3(N__17217),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_17_19_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_17_19_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_17_19_2  (
            .in0(N__28719),
            .in1(N__28661),
            .in2(N__17202),
            .in3(N__28587),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_17_19_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_17_19_3 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_17_19_3  (
            .in0(N__28662),
            .in1(N__17199),
            .in2(N__17193),
            .in3(N__17475),
            .lcout(M_this_ppu_vram_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_11_LC_17_19_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_11_LC_17_19_5 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_11_LC_17_19_5 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \this_sprites_ram.mem_radreg_11_LC_17_19_5  (
            .in0(N__17157),
            .in1(N__17151),
            .in2(N__31882),
            .in3(N__32124),
            .lcout(\this_sprites_ram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32553),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_17_19_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_17_19_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_17_19_7  (
            .in0(N__30101),
            .in1(N__17505),
            .in2(_gnd_net_),
            .in3(N__17490),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_2_LC_17_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_2_LC_17_20_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_2_LC_17_20_5 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \this_ppu.M_state_q_2_LC_17_20_5  (
            .in0(N__17469),
            .in1(N__17427),
            .in2(_gnd_net_),
            .in3(N__17409),
            .lcout(\this_ppu.M_state_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32566),
            .ce(),
            .sr(N__26046));
    defparam m1_LC_17_21_0.C_ON=1'b0;
    defparam m1_LC_17_21_0.SEQ_MODE=4'b0000;
    defparam m1_LC_17_21_0.LUT_INIT=16'b1100110001100110;
    LogicCell40 m1_LC_17_21_0 (
            .in0(N__17886),
            .in1(N__17929),
            .in2(_gnd_net_),
            .in3(N__18078),
            .lcout(),
            .ltout(N_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIRPN94A_2_LC_17_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIRPN94A_2_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIRPN94A_2_LC_17_21_1 .LUT_INIT=16'b1101101100100100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIRPN94A_2_LC_17_21_1  (
            .in0(N__22840),
            .in1(N__22715),
            .in2(N__17391),
            .in3(N__17514),
            .lcout(),
            .ltout(\this_vga_signals.N_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI75QSCH1_2_LC_17_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI75QSCH1_2_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI75QSCH1_2_LC_17_21_2 .LUT_INIT=16'b1000101101000111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI75QSCH1_2_LC_17_21_2  (
            .in0(N__17367),
            .in1(N__17826),
            .in2(N__17388),
            .in3(N__17379),
            .lcout(\this_vga_signals.vaddress_N_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_17_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_17_21_3 .LUT_INIT=16'b1011010001001011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_17_21_3  (
            .in0(N__18080),
            .in1(N__17885),
            .in2(N__18009),
            .in3(N__17838),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_17_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_17_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_11_LC_17_21_4  (
            .in0(N__17871),
            .in1(N__17547),
            .in2(N__17910),
            .in3(N__18007),
            .lcout(\this_vga_signals.mult1_un75_sum_axb1_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIDON0D8_3_LC_17_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIDON0D8_3_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIDON0D8_3_LC_17_21_5 .LUT_INIT=16'b1001011011000011;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIDON0D8_3_LC_17_21_5  (
            .in0(N__18079),
            .in1(N__22839),
            .in2(N__17934),
            .in3(N__17884),
            .lcout(\this_vga_signals.N_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_m2_LC_17_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_m2_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_m2_LC_17_21_6 .LUT_INIT=16'b1011001000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_m2_LC_17_21_6  (
            .in0(N__22714),
            .in1(N__18324),
            .in2(N__22865),
            .in3(N__17597),
            .lcout(\this_vga_signals.mult1_un68_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIKLMK17_2_LC_17_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIKLMK17_2_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIKLMK17_2_LC_17_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIKLMK17_2_LC_17_21_7  (
            .in0(N__18027),
            .in1(N__17953),
            .in2(N__17553),
            .in3(N__17820),
            .lcout(\this_vga_signals.g0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_0_LC_17_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_0_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_0_LC_17_22_0 .LUT_INIT=16'b1010101001011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_0_LC_17_22_0  (
            .in0(N__18297),
            .in1(N__18099),
            .in2(N__23277),
            .in3(N__19008),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_17_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_17_22_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_17_22_1  (
            .in0(N__18230),
            .in1(_gnd_net_),
            .in2(N__17550),
            .in3(N__18767),
            .lcout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_17_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_17_22_2 .LUT_INIT=16'b0001011100101011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_17_22_2  (
            .in0(N__18766),
            .in1(N__23266),
            .in2(N__22868),
            .in3(N__18231),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m2_3_1_LC_17_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m2_3_1_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m2_3_1_LC_17_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m2_3_1_LC_17_22_3  (
            .in0(N__18232),
            .in1(N__17546),
            .in2(N__17958),
            .in3(N__17928),
            .lcout(\this_vga_signals.if_m2_3_1 ),
            .ltout(\this_vga_signals.if_m2_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIBALLEF_2_LC_17_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIBALLEF_2_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIBALLEF_2_LC_17_22_4 .LUT_INIT=16'b0001010001000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIBALLEF_2_LC_17_22_4  (
            .in0(N__22706),
            .in1(N__18033),
            .in2(N__17535),
            .in3(N__18008),
            .lcout(),
            .ltout(\this_vga_signals.g2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIOP5EV51_1_LC_17_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIOP5EV51_1_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIOP5EV51_1_LC_17_22_5 .LUT_INIT=16'b0000101111110100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIOP5EV51_1_LC_17_22_5  (
            .in0(N__17985),
            .in1(N__22934),
            .in2(N__17532),
            .in3(N__17529),
            .lcout(\this_vga_signals.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m1_0_LC_17_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m1_0_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m1_0_LC_17_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m1_0_LC_17_22_6  (
            .in0(N__18768),
            .in1(N__23267),
            .in2(_gnd_net_),
            .in3(N__18229),
            .lcout(\this_vga_signals.if_m1_0 ),
            .ltout(\this_vga_signals.if_m1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m1_9_0_LC_17_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m1_9_0_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m1_9_0_LC_17_22_7 .LUT_INIT=16'b1101001110111100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m1_9_0_LC_17_22_7  (
            .in0(N__18323),
            .in1(N__22854),
            .in2(N__17517),
            .in3(N__22705),
            .lcout(\this_vga_signals.if_m1_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIVGRQM1_1_LC_17_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIVGRQM1_1_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIVGRQM1_1_LC_17_23_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIVGRQM1_1_LC_17_23_0  (
            .in0(N__18249),
            .in1(N__22933),
            .in2(_gnd_net_),
            .in3(N__18120),
            .lcout(\this_vga_signals.N_129_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_17_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_17_23_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_17_23_1  (
            .in0(_gnd_net_),
            .in1(N__23259),
            .in2(_gnd_net_),
            .in3(N__18762),
            .lcout(\this_vga_signals.if_m1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_17_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_17_23_2 .LUT_INIT=16'b1011001000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_LC_17_23_2  (
            .in0(N__22707),
            .in1(N__18316),
            .in2(N__22869),
            .in3(N__17598),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_LC_17_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_LC_17_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_0_a3_LC_17_23_3  (
            .in0(N__18114),
            .in1(N__18763),
            .in2(N__18108),
            .in3(N__18251),
            .lcout(\this_vga_signals.g0_3_0_a3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_17_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_17_23_4 .LUT_INIT=16'b0001011100101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_LC_17_23_4  (
            .in0(N__18250),
            .in1(N__22857),
            .in2(N__23282),
            .in3(N__18781),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_17_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_17_23_5 .LUT_INIT=16'b1001111111111001;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_LC_17_23_5  (
            .in0(N__18782),
            .in1(N__18247),
            .in2(N__23099),
            .in3(N__20667),
            .lcout(\this_vga_signals.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_1_LC_17_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_1_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_1_LC_17_23_6 .LUT_INIT=16'b0001011100101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_1_LC_17_23_6  (
            .in0(N__18248),
            .in1(N__22856),
            .in2(N__23283),
            .in3(N__18783),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c2_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_17_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_17_23_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_LC_17_23_7  (
            .in0(N__22361),
            .in1(N__18126),
            .in2(N__17565),
            .in3(N__18138),
            .lcout(\this_vga_signals.g0_i_x4_7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_9_N_2L1_LC_17_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_9_N_2L1_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_9_N_2L1_LC_17_24_0 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_9_N_2L1_LC_17_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23284),
            .in3(N__18772),
            .lcout(),
            .ltout(\this_vga_signals.g0_9_N_2L1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_9_N_3L3_LC_17_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_9_N_3L3_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_9_N_3L3_LC_17_24_1 .LUT_INIT=16'b0101100010000101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_9_N_3L3_LC_17_24_1  (
            .in0(N__22866),
            .in1(N__18636),
            .in2(N__17556),
            .in3(N__18242),
            .lcout(\this_vga_signals.g0_9_N_3L3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_1_LC_17_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_1_LC_17_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_1_LC_17_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_1_LC_17_24_2  (
            .in0(N__18924),
            .in1(N__18270),
            .in2(_gnd_net_),
            .in3(N__20372),
            .lcout(),
            .ltout(\this_vga_signals.g0_i_x4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_3_LC_17_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_3_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_3_LC_17_24_3 .LUT_INIT=16'b0001011101110001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_3_LC_17_24_3  (
            .in0(N__22867),
            .in1(N__23272),
            .in2(N__17685),
            .in3(N__18243),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c2_0_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_17_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_17_24_4 .LUT_INIT=16'b0001010001000001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_9_LC_17_24_4  (
            .in0(N__22708),
            .in1(N__18168),
            .in2(N__17682),
            .in3(N__17679),
            .lcout(\this_vga_signals.g0_i_a4_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_a0_LC_17_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_a0_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_a0_LC_17_24_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_a0_LC_17_24_6  (
            .in0(_gnd_net_),
            .in1(N__20580),
            .in2(_gnd_net_),
            .in3(N__20520),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI7F791_13_LC_18_16_6.C_ON=1'b0;
    defparam M_this_state_q_RNI7F791_13_LC_18_16_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI7F791_13_LC_18_16_6.LUT_INIT=16'b1110111010101010;
    LogicCell40 M_this_state_q_RNI7F791_13_LC_18_16_6 (
            .in0(N__26206),
            .in1(N__19092),
            .in2(_gnd_net_),
            .in3(N__24227),
            .lcout(N_1422_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_3_LC_18_17_0.C_ON=1'b0;
    defparam M_this_data_count_q_3_LC_18_17_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_18_17_0.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_3_LC_18_17_0 (
            .in0(N__28965),
            .in1(N__29212),
            .in2(_gnd_net_),
            .in3(N__28979),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32546),
            .ce(N__29108),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_14_LC_18_18_3.C_ON=1'b0;
    defparam M_this_data_count_q_14_LC_18_18_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_14_LC_18_18_3.LUT_INIT=16'b1100000010101010;
    LogicCell40 M_this_data_count_q_14_LC_18_18_3 (
            .in0(N__29295),
            .in1(N__26963),
            .in2(N__28167),
            .in3(N__29188),
            .lcout(M_this_data_count_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32554),
            .ce(N__29103),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIICAO1_0_LC_18_19_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIICAO1_0_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIICAO1_0_LC_18_19_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIICAO1_0_LC_18_19_0  (
            .in0(N__19628),
            .in1(N__18673),
            .in2(N__19705),
            .in3(N__18684),
            .lcout(M_this_state_d_0_sqmuxa_2),
            .ltout(M_this_state_d_0_sqmuxa_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_LC_18_19_1.C_ON=1'b0;
    defparam M_this_substate_q_LC_18_19_1.SEQ_MODE=4'b1000;
    defparam M_this_substate_q_LC_18_19_1.LUT_INIT=16'b1111000011111010;
    LogicCell40 M_this_substate_q_LC_18_19_1 (
            .in0(N__18674),
            .in1(_gnd_net_),
            .in2(N__17601),
            .in3(N__18690),
            .lcout(M_this_substate_qZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32567),
            .ce(),
            .sr(N__26049));
    defparam \this_start_data_delay.M_last_q_RNILCRA6_LC_18_19_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNILCRA6_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNILCRA6_LC_18_19_4 .LUT_INIT=16'b0100111001011111;
    LogicCell40 \this_start_data_delay.M_last_q_RNILCRA6_LC_18_19_4  (
            .in0(N__26967),
            .in1(N__26196),
            .in2(N__24462),
            .in3(N__24624),
            .lcout(M_this_data_count_q_3_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_3_LC_18_20_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_3_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_3_LC_18_20_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIK0EI1_3_LC_18_20_0  (
            .in0(N__19704),
            .in1(N__19627),
            .in2(N__19569),
            .in3(N__19490),
            .lcout(\this_start_data_delay.N_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.dmalto4_0_a2_0_1_LC_18_20_1 .C_ON=1'b0;
    defparam \this_start_data_delay.dmalto4_0_a2_0_1_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.dmalto4_0_a2_0_1_LC_18_20_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_start_data_delay.dmalto4_0_a2_0_1_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__21262),
            .in2(_gnd_net_),
            .in3(N__23780),
            .lcout(\this_start_data_delay.N_76_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_1_LC_18_20_2.C_ON=1'b0;
    defparam M_this_state_q_1_LC_18_20_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_18_20_2.LUT_INIT=16'b0101000001010100;
    LogicCell40 M_this_state_q_1_LC_18_20_2 (
            .in0(N__26207),
            .in1(N__21319),
            .in2(N__17787),
            .in3(N__24224),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32574),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_2_LC_18_20_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_2_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_2_LC_18_20_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIK0EI1_2_LC_18_20_4  (
            .in0(N__19703),
            .in1(N__19626),
            .in2(N__19568),
            .in3(N__19491),
            .lcout(),
            .ltout(\this_start_data_delay.N_65_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_18_20_5.C_ON=1'b0;
    defparam M_this_state_q_4_LC_18_20_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_18_20_5.LUT_INIT=16'b0000000011110100;
    LogicCell40 M_this_state_q_4_LC_18_20_5 (
            .in0(N__24225),
            .in1(N__21263),
            .in2(N__17778),
            .in3(N__26208),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32574),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.dmalto4_0_o2_0_LC_18_20_6 .C_ON=1'b0;
    defparam \this_start_data_delay.dmalto4_0_o2_0_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.dmalto4_0_o2_0_LC_18_20_6 .LUT_INIT=16'b1110111011100000;
    LogicCell40 \this_start_data_delay.dmalto4_0_o2_0_LC_18_20_6  (
            .in0(N__23781),
            .in1(N__21100),
            .in2(N__24313),
            .in3(N__21318),
            .lcout(\this_start_data_delay.N_42_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.dmalto4_0_a2_LC_18_20_7 .C_ON=1'b0;
    defparam \this_start_data_delay.dmalto4_0_a2_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.dmalto4_0_a2_LC_18_20_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_start_data_delay.dmalto4_0_a2_LC_18_20_7  (
            .in0(N__17762),
            .in1(N__23571),
            .in2(N__18399),
            .in3(N__19431),
            .lcout(dma_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_2_LC_18_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_2_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_2_LC_18_21_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_2_LC_18_21_0  (
            .in0(N__22270),
            .in1(N__20245),
            .in2(N__20373),
            .in3(N__18884),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2 ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_LC_18_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_LC_18_21_1 .LUT_INIT=16'b0000111100000110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_LC_18_21_1  (
            .in0(N__20371),
            .in1(N__22272),
            .in2(N__17688),
            .in3(N__17799),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_LC_18_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_LC_18_21_2 .LUT_INIT=16'b1101000001110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_LC_18_21_2  (
            .in0(N__18797),
            .in1(N__18785),
            .in2(N__17889),
            .in3(N__18257),
            .lcout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3),
            .ltout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_18_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_18_21_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_18_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17874),
            .in3(N__18081),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m4_LC_18_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m4_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m4_LC_18_21_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m4_LC_18_21_4  (
            .in0(N__17865),
            .in1(N__17847),
            .in2(N__17841),
            .in3(N__17837),
            .lcout(\this_vga_signals.if_i4_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIKL00E1_2_LC_18_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIKL00E1_2_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIKL00E1_2_LC_18_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIKL00E1_2_LC_18_21_5  (
            .in0(N__18258),
            .in1(N__22858),
            .in2(_gnd_net_),
            .in3(N__22713),
            .lcout(\this_vga_signals.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_1_LC_18_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_1_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_1_LC_18_21_6 .LUT_INIT=16'b0001101110101011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_1_LC_18_21_6  (
            .in0(N__22269),
            .in1(N__18883),
            .in2(N__17814),
            .in3(N__20423),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_0_2_1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_0_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_18_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_18_21_7 .LUT_INIT=16'b1111001111111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_0_LC_18_21_7  (
            .in0(_gnd_net_),
            .in1(N__20370),
            .in2(N__17793),
            .in3(N__22271),
            .lcout(\this_vga_signals.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_18_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_18_22_0 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_18_22_0  (
            .in0(N__20660),
            .in1(N__23000),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_0_LC_18_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_0_LC_18_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_0_LC_18_22_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_0_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17790),
            .in3(N__18764),
            .lcout(\this_vga_signals.mult1_un61_sum_axb2_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axb2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_LC_18_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_LC_18_22_2 .LUT_INIT=16'b0000100000100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_LC_18_22_2  (
            .in0(N__22849),
            .in1(N__18233),
            .in2(N__18084),
            .in3(N__17975),
            .lcout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d),
            .ltout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_18_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_18_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_18_22_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_LC_18_22_3  (
            .in0(N__18063),
            .in1(N__18047),
            .in2(N__18036),
            .in3(N__18132),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_18_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_18_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_LC_18_22_4  (
            .in0(N__17906),
            .in1(N__18026),
            .in2(N__18012),
            .in3(N__18003),
            .lcout(\this_vga_signals.mult1_un75_sum_axb1_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_18_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_18_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_19_LC_18_22_5  (
            .in0(_gnd_net_),
            .in1(N__20661),
            .in2(N__23039),
            .in3(N__18765),
            .lcout(),
            .ltout(\this_vga_signals.N_4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_18_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_18_22_6 .LUT_INIT=16'b1000000000000010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_12_LC_18_22_6  (
            .in0(N__22850),
            .in1(N__18234),
            .in2(N__17979),
            .in3(N__17976),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_d_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_1_LC_18_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_1_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_1_LC_18_22_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_1_LC_18_22_7  (
            .in0(N__18235),
            .in1(N__17957),
            .in2(N__22716),
            .in3(N__17933),
            .lcout(\this_vga_signals.mult1_un75_sum_axb1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_ns_LC_18_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_ns_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_ns_LC_18_23_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_ns_LC_18_23_0  (
            .in0(N__19023),
            .in1(N__20366),
            .in2(_gnd_net_),
            .in3(N__18930),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_18_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_18_23_1 .LUT_INIT=16'b0000111100000001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_18_23_1  (
            .in0(N__19014),
            .in1(N__19000),
            .in2(N__17895),
            .in3(N__18292),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_18_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_18_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_18_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_28_LC_18_23_2  (
            .in0(_gnd_net_),
            .in1(N__23202),
            .in2(N__17892),
            .in3(N__18777),
            .lcout(),
            .ltout(\this_vga_signals.N_4_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_18_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_18_23_3 .LUT_INIT=16'b0001101001111010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_25_LC_18_23_3  (
            .in0(N__22855),
            .in1(N__22702),
            .in2(N__18141),
            .in3(N__20610),
            .lcout(\this_vga_signals.N_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_LC_18_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_LC_18_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_LC_18_23_5 .LUT_INIT=16'b1011111001111101;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_LC_18_23_5  (
            .in0(N__18776),
            .in1(N__20589),
            .in2(N__23092),
            .in3(N__18236),
            .lcout(\this_vga_signals.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_1_LC_18_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_1_LC_18_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_1_LC_18_23_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_1_LC_18_23_6  (
            .in0(N__20656),
            .in1(N__23069),
            .in2(_gnd_net_),
            .in3(N__20691),
            .lcout(\this_vga_signals.g0_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_18_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_18_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_18_23_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_18_23_7  (
            .in0(_gnd_net_),
            .in1(N__20297),
            .in2(_gnd_net_),
            .in3(N__20655),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_0_8_LC_18_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_0_8_LC_18_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_0_8_LC_18_24_0 .LUT_INIT=16'b1101100101001101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_0_8_LC_18_24_0  (
            .in0(N__22578),
            .in1(N__21901),
            .in2(N__20183),
            .in3(N__21985),
            .lcout(\this_vga_signals.SUM_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNISDV89_4_LC_18_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNISDV89_4_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNISDV89_4_LC_18_24_1 .LUT_INIT=16'b0010110110000111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNISDV89_4_LC_18_24_1  (
            .in0(N__18984),
            .in1(N__18162),
            .in2(N__23203),
            .in3(N__20151),
            .lcout(\this_vga_signals.N_24_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_18_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_18_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_18_24_2 .LUT_INIT=16'b1011101100011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_2_LC_18_24_2  (
            .in0(N__23268),
            .in1(N__18098),
            .in2(N__23097),
            .in3(N__20654),
            .lcout(\this_vga_signals.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_3_LC_18_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_3_LC_18_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_3_LC_18_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_0_a3_3_LC_18_24_3  (
            .in0(N__20653),
            .in1(N__18828),
            .in2(N__20274),
            .in3(N__22387),
            .lcout(\this_vga_signals.g0_3_0_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_18_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_18_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_18_24_4  (
            .in0(N__23077),
            .in1(N__23158),
            .in2(_gnd_net_),
            .in3(N__20652),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_x4_LC_18_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_x4_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_x4_LC_18_24_5 .LUT_INIT=16'b0010110011010011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_x4_LC_18_24_5  (
            .in0(N__23159),
            .in1(N__19004),
            .in2(N__18327),
            .in3(N__18293),
            .lcout(\this_vga_signals.if_N_9_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_18_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_18_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_18_24_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_18_24_6  (
            .in0(N__18978),
            .in1(_gnd_net_),
            .in2(N__18882),
            .in3(N__20651),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_m2_LC_18_25_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_m2_LC_18_25_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_m2_LC_18_25_3 .LUT_INIT=16'b0110111100001001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_m2_LC_18_25_3  (
            .in0(N__18660),
            .in1(N__18276),
            .in2(N__18909),
            .in3(N__18920),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_1_0 ),
            .ltout(\this_vga_signals.mult1_un47_sum_c3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_4_LC_18_25_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_4_LC_18_25_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_4_LC_18_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_4_LC_18_25_4  (
            .in0(N__18897),
            .in1(N__18784),
            .in2(N__18264),
            .in3(N__18259),
            .lcout(\this_vga_signals.g2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_7_LC_18_26_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_7_LC_18_26_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_7_LC_18_26_3 .LUT_INIT=16'b0001001111101100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_7_LC_18_26_3  (
            .in0(N__23183),
            .in1(N__22362),
            .in2(N__23098),
            .in3(N__21999),
            .lcout(\this_vga_signals.m12_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_19_16_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_19_16_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_19_16_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_19_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_16_LC_19_16_1.C_ON=1'b0;
    defparam M_this_state_q_16_LC_19_16_1.SEQ_MODE=4'b1000;
    defparam M_this_state_q_16_LC_19_16_1.LUT_INIT=16'b0000110000001010;
    LogicCell40 M_this_state_q_16_LC_19_16_1 (
            .in0(N__19394),
            .in1(N__19144),
            .in2(N__26226),
            .in3(N__24231),
            .lcout(M_this_state_qZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32547),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_14_LC_19_17_0.C_ON=1'b0;
    defparam M_this_state_q_14_LC_19_17_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_14_LC_19_17_0.LUT_INIT=16'b0000110000001010;
    LogicCell40 M_this_state_q_14_LC_19_17_0 (
            .in0(N__19115),
            .in1(N__19091),
            .in2(N__26225),
            .in3(N__24239),
            .lcout(M_this_state_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32555),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un25_i_a2_3_a2_2_a3_3_LC_19_17_5 .C_ON=1'b0;
    defparam \this_start_data_delay.un25_i_a2_3_a2_2_a3_3_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un25_i_a2_3_a2_2_a3_3_LC_19_17_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_start_data_delay.un25_i_a2_3_a2_2_a3_3_LC_19_17_5  (
            .in0(N__23489),
            .in1(N__19764),
            .in2(N__20741),
            .in3(N__19427),
            .lcout(\this_start_data_delay.N_400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_12_LC_19_17_7.C_ON=1'b0;
    defparam M_this_state_q_12_LC_19_17_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_12_LC_19_17_7.LUT_INIT=16'b0011001100110010;
    LogicCell40 M_this_state_q_12_LC_19_17_7 (
            .in0(N__18387),
            .in1(N__26214),
            .in2(N__26786),
            .in3(N__18483),
            .lcout(M_this_state_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32555),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un25_i_a2_i_o2_4_LC_19_18_2 .C_ON=1'b0;
    defparam \this_start_data_delay.un25_i_a2_i_o2_4_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un25_i_a2_i_o2_4_LC_19_18_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_start_data_delay.un25_i_a2_i_o2_4_LC_19_18_2  (
            .in0(_gnd_net_),
            .in1(N__18482),
            .in2(_gnd_net_),
            .in3(N__19395),
            .lcout(\this_start_data_delay.N_55_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_ns_0_i_o2_0_LC_19_18_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_ns_0_i_o2_0_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_ns_0_i_o2_0_LC_19_18_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.M_this_state_q_ns_0_i_o2_0_LC_19_18_4  (
            .in0(N__22167),
            .in1(N__21093),
            .in2(N__24317),
            .in3(N__21320),
            .lcout(\this_start_data_delay.N_112_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.dmalto4_0_a2_1_LC_19_18_5 .C_ON=1'b0;
    defparam \this_start_data_delay.dmalto4_0_a2_1_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.dmalto4_0_a2_1_LC_19_18_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.dmalto4_0_a2_1_LC_19_18_5  (
            .in0(N__23906),
            .in1(N__19755),
            .in2(N__23496),
            .in3(N__20730),
            .lcout(\this_start_data_delay.dmalto4_0_a2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_data_count_qlde_i_o2_1_LC_19_18_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_data_count_qlde_i_o2_1_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_data_count_qlde_i_o2_1_LC_19_18_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_start_data_delay.M_this_data_count_qlde_i_o2_1_LC_19_18_6  (
            .in0(N__20729),
            .in1(N__19754),
            .in2(_gnd_net_),
            .in3(N__23905),
            .lcout(\this_start_data_delay.N_90_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNICA9G3_0_LC_19_18_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNICA9G3_0_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNICA9G3_0_LC_19_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNICA9G3_0_LC_19_18_7  (
            .in0(_gnd_net_),
            .in1(N__20731),
            .in2(_gnd_net_),
            .in3(N__23663),
            .lcout(\this_start_data_delay.N_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_3_LC_19_19_0.C_ON=1'b0;
    defparam M_this_state_q_3_LC_19_19_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_19_19_0.LUT_INIT=16'b0101000001010100;
    LogicCell40 M_this_state_q_3_LC_19_19_0 (
            .in0(N__26211),
            .in1(N__22171),
            .in2(N__18381),
            .in3(N__24240),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32575),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI3MH61_LC_19_19_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI3MH61_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI3MH61_LC_19_19_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI3MH61_LC_19_19_2  (
            .in0(N__18372),
            .in1(N__31596),
            .in2(N__18354),
            .in3(N__23733),
            .lcout(\this_start_data_delay.N_47_0 ),
            .ltout(\this_start_data_delay.N_47_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIVMHD1_LC_19_19_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIVMHD1_LC_19_19_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIVMHD1_LC_19_19_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIVMHD1_LC_19_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18333),
            .in3(N__19932),
            .lcout(\this_start_data_delay.N_48_0 ),
            .ltout(\this_start_data_delay.N_48_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_LC_19_19_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_LC_19_19_4 .LUT_INIT=16'b0111000001100000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIK0EI1_LC_19_19_4  (
            .in0(N__19687),
            .in1(N__19550),
            .in2(N__18330),
            .in3(N__19620),
            .lcout(N_28_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI7R5F1_LC_19_19_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI7R5F1_LC_19_19_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI7R5F1_LC_19_19_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI7R5F1_LC_19_19_6  (
            .in0(N__19933),
            .in1(N__19549),
            .in2(_gnd_net_),
            .in3(N__19967),
            .lcout(\this_start_data_delay.N_82 ),
            .ltout(\this_start_data_delay.N_82_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIICAO1_LC_19_19_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIICAO1_LC_19_19_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIICAO1_LC_19_19_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIICAO1_LC_19_19_7  (
            .in0(N__19619),
            .in1(N__19686),
            .in2(N__18678),
            .in3(N__18675),
            .lcout(\this_start_data_delay.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_x4_LC_19_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_x4_LC_19_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_x4_LC_19_20_0 .LUT_INIT=16'b1110110000010011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_x4_LC_19_20_0  (
            .in0(N__20504),
            .in1(N__22265),
            .in2(N__20579),
            .in3(N__21951),
            .lcout(\this_vga_signals.g0_0_x4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_19_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_19_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_19_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_19_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21715),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32585),
            .ce(N__23407),
            .sr(N__23313));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_0_LC_19_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_0_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_0_LC_19_20_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_0_LC_19_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20130),
            .in3(N__20028),
            .lcout(\this_vga_signals.vaddress_c2 ),
            .ltout(\this_vga_signals.vaddress_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_19_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_19_20_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_24_LC_19_20_3  (
            .in0(N__21949),
            .in1(N__20084),
            .in2(N__18648),
            .in3(N__22570),
            .lcout(),
            .ltout(\this_vga_signals.N_5_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_1_LC_19_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_1_LC_19_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_1_LC_19_20_4 .LUT_INIT=16'b0000110100001011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_1_LC_19_20_4  (
            .in0(N__22571),
            .in1(N__21897),
            .in2(N__18645),
            .in3(N__21950),
            .lcout(),
            .ltout(\this_vga_signals.g0_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_19_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_19_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_19_20_5 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_1_LC_19_20_5  (
            .in0(N__18804),
            .in1(N__19992),
            .in2(N__18642),
            .in3(N__19986),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_19_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_19_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_19_20_6 .LUT_INIT=16'b0111100010110100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_21_LC_19_20_6  (
            .in0(N__23221),
            .in1(N__23065),
            .in2(N__18639),
            .in3(N__20666),
            .lcout(\this_vga_signals.N_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_19_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_19_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_19_20_7 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_0_LC_19_20_7  (
            .in0(N__22264),
            .in1(N__20572),
            .in2(_gnd_net_),
            .in3(N__20503),
            .lcout(\this_vga_signals.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_19_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_19_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_0_LC_19_21_0  (
            .in0(N__22703),
            .in1(N__18798),
            .in2(N__22860),
            .in3(N__18786),
            .lcout(\this_vga_signals.g0_5_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_19_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_19_21_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_19_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_19_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21385),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32591),
            .ce(N__23360),
            .sr(N__23315));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_19_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_19_21_4 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_19_21_4  (
            .in0(N__20552),
            .in1(N__20502),
            .in2(_gnd_net_),
            .in3(N__20073),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_19_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_19_21_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_19_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_19_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21720),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32591),
            .ce(N__23360),
            .sr(N__23315));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_a4_LC_19_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_a4_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_a4_LC_19_21_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_a4_LC_19_21_6  (
            .in0(N__21775),
            .in1(N__20072),
            .in2(N__20247),
            .in3(N__22545),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_0_a4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_1_LC_19_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_1_LC_19_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_1_LC_19_21_7 .LUT_INIT=16'b1101111111111011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_1_LC_19_21_7  (
            .in0(N__22544),
            .in1(N__21819),
            .in2(N__20086),
            .in3(N__20233),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_19_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_19_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_19_22_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_19_22_2  (
            .in0(N__22994),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23201),
            .lcout(\this_vga_signals.vaddress_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_19_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_19_22_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_19_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_19_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21353),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32600),
            .ce(N__23397),
            .sr(N__23318));
    defparam \this_vga_signals.un5_vaddress_g2_1_0_LC_19_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_1_0_LC_19_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_1_0_LC_19_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_1_0_LC_19_22_4  (
            .in0(N__22995),
            .in1(N__22843),
            .in2(_gnd_net_),
            .in3(N__22672),
            .lcout(\this_vga_signals.g2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_19_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_19_22_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_19_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_19_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21354),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32600),
            .ce(N__23397),
            .sr(N__23318));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_ns_LC_19_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_ns_LC_19_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_ns_LC_19_22_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_ns_LC_19_22_6  (
            .in0(_gnd_net_),
            .in1(N__20126),
            .in2(N__20007),
            .in3(N__20262),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_602_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_22_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21352),
            .lcout(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32600),
            .ce(N__23397),
            .sr(N__23318));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_LC_19_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_LC_19_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_LC_19_23_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_LC_19_23_0  (
            .in0(N__18839),
            .in1(N__21735),
            .in2(N__18855),
            .in3(N__18818),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_19_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_19_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_19_23_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_LC_19_23_1  (
            .in0(N__18819),
            .in1(N__18854),
            .in2(N__22020),
            .in3(N__18840),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_2_LC_19_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_2_LC_19_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_2_LC_19_23_2 .LUT_INIT=16'b0110110000110110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_2_LC_19_23_2  (
            .in0(N__18953),
            .in1(N__20334),
            .in2(N__20456),
            .in3(N__20414),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_3_ns_LC_19_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_3_ns_LC_19_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_3_ns_LC_19_23_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_3_ns_LC_19_23_3  (
            .in0(_gnd_net_),
            .in1(N__20697),
            .in2(_gnd_net_),
            .in3(N__20246),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_19_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_19_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_19_23_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_19_23_4  (
            .in0(N__20100),
            .in1(N__21734),
            .in2(N__18822),
            .in3(N__18817),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_x1_LC_19_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_x1_LC_19_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_x1_LC_19_23_5 .LUT_INIT=16'b0000111010000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_x1_LC_19_23_5  (
            .in0(N__20450),
            .in1(N__18952),
            .in2(N__18807),
            .in3(N__18977),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_4_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_19_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_19_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_19_23_6 .LUT_INIT=16'b1001000111011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_19_23_6  (
            .in0(N__18951),
            .in1(N__20333),
            .in2(N__20455),
            .in3(N__20413),
            .lcout(\this_vga_signals.mult1_un47_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un47_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_19_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_19_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_19_23_7 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_19_23_7  (
            .in0(N__20514),
            .in1(_gnd_net_),
            .in2(N__19017),
            .in3(N__20565),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_19_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_19_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_19_24_0 .LUT_INIT=16'b0000111000000110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_19_24_0  (
            .in0(N__20351),
            .in1(N__18962),
            .in2(N__20457),
            .in3(N__20410),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI6FO86_LC_19_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI6FO86_LC_19_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI6FO86_LC_19_24_1 .LUT_INIT=16'b0000010110100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI6FO86_LC_19_24_1  (
            .in0(N__20412),
            .in1(_gnd_net_),
            .in2(N__18966),
            .in3(N__20454),
            .lcout(\this_vga_signals.i1_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_0_LC_19_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_0_LC_19_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_0_LC_19_24_3 .LUT_INIT=16'b0001000111101110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_0_LC_19_24_3  (
            .in0(N__20509),
            .in1(N__20569),
            .in2(_gnd_net_),
            .in3(N__20087),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc1_0 ),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_x0_LC_19_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_x0_LC_19_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_x0_LC_19_24_4 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_x0_LC_19_24_4  (
            .in0(_gnd_net_),
            .in1(N__18961),
            .in2(N__18933),
            .in3(N__20409),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_4_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_6_LC_19_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_6_LC_19_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_6_LC_19_24_5 .LUT_INIT=16'b0100011101110001;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_6_LC_19_24_5  (
            .in0(N__20411),
            .in1(N__22334),
            .in2(N__20519),
            .in3(N__20570),
            .lcout(\this_vga_signals.g1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_19_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_19_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_19_24_6 .LUT_INIT=16'b1010010100001111;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_19_24_6  (
            .in0(N__20571),
            .in1(_gnd_net_),
            .in2(N__22363),
            .in3(N__20513),
            .lcout(\this_vga_signals.vaddress_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_19_25_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_19_25_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_19_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_19_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21390),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32624),
            .ce(N__23409),
            .sr(N__23319));
    defparam \this_ppu.M_haddress_q_RNIOC7O_0_LC_19_31_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIOC7O_0_LC_19_31_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIOC7O_0_LC_19_31_2 .LUT_INIT=16'b0101011101010100;
    LogicCell40 \this_ppu.M_haddress_q_RNIOC7O_0_LC_19_31_2  (
            .in0(N__19353),
            .in1(N__32075),
            .in2(N__31939),
            .in3(N__19334),
            .lcout(M_this_ppu_sprites_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNILR691_LC_20_16_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNILR691_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNILR691_LC_20_16_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNILR691_LC_20_16_1  (
            .in0(N__26187),
            .in1(N__21099),
            .in2(_gnd_net_),
            .in3(N__24158),
            .lcout(\this_start_data_delay.N_993 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_13_LC_20_16_2.C_ON=1'b0;
    defparam M_this_state_q_13_LC_20_16_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_13_LC_20_16_2.LUT_INIT=16'b0011000100110000;
    LogicCell40 M_this_state_q_13_LC_20_16_2 (
            .in0(N__24159),
            .in1(N__26188),
            .in2(N__20709),
            .in3(N__19087),
            .lcout(M_this_state_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32556),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_15_LC_20_16_4.C_ON=1'b0;
    defparam M_this_state_q_15_LC_20_16_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_15_LC_20_16_4.LUT_INIT=16'b0011001000010000;
    LogicCell40 M_this_state_q_15_LC_20_16_4 (
            .in0(N__24160),
            .in1(N__26189),
            .in2(N__19145),
            .in3(N__19111),
            .lcout(M_this_state_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32556),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_o2_LC_20_16_6 .C_ON=1'b0;
    defparam \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_o2_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_o2_LC_20_16_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_o2_LC_20_16_6  (
            .in0(N__19137),
            .in1(N__19110),
            .in2(_gnd_net_),
            .in3(N__19086),
            .lcout(\this_start_data_delay.N_80_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIHQLO2_LC_20_16_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIHQLO2_LC_20_16_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIHQLO2_LC_20_16_7 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \this_start_data_delay.M_last_q_RNIHQLO2_LC_20_16_7  (
            .in0(N__19068),
            .in1(N__26255),
            .in2(_gnd_net_),
            .in3(N__24157),
            .lcout(\this_start_data_delay.M_this_state_q_ns_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_o2_0_LC_20_17_0 .C_ON=1'b0;
    defparam \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_o2_0_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_o2_0_LC_20_17_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_o2_0_LC_20_17_0  (
            .in0(N__19455),
            .in1(N__19058),
            .in2(_gnd_net_),
            .in3(N__23955),
            .lcout(\this_start_data_delay.N_89_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_a2_LC_20_17_2 .C_ON=1'b0;
    defparam \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_a2_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_a2_LC_20_17_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_a2_LC_20_17_2  (
            .in0(_gnd_net_),
            .in1(N__19390),
            .in2(_gnd_net_),
            .in3(N__19059),
            .lcout(),
            .ltout(\this_start_data_delay.un1_M_this_state_q_1_i_a2_0_aZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_external_address_qlde_i_a3_0_LC_20_17_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_external_address_qlde_i_a3_0_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_external_address_qlde_i_a3_0_LC_20_17_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_start_data_delay.M_this_external_address_qlde_i_a3_0_LC_20_17_3  (
            .in0(N__23956),
            .in1(N__19456),
            .in2(N__19050),
            .in3(N__19047),
            .lcout(\this_start_data_delay.N_122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIA89G3_LC_20_17_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIA89G3_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIA89G3_LC_20_17_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIA89G3_LC_20_17_4  (
            .in0(N__23727),
            .in1(N__19763),
            .in2(_gnd_net_),
            .in3(N__26877),
            .lcout(),
            .ltout(\this_start_data_delay.N_127_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_11_LC_20_17_5.C_ON=1'b0;
    defparam M_this_state_q_11_LC_20_17_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_11_LC_20_17_5.LUT_INIT=16'b0011000000110010;
    LogicCell40 M_this_state_q_11_LC_20_17_5 (
            .in0(N__19458),
            .in1(N__26218),
            .in2(N__19461),
            .in3(N__24217),
            .lcout(M_this_state_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32568),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIP7R11_LC_20_18_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIP7R11_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIP7R11_LC_20_18_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIP7R11_LC_20_18_1  (
            .in0(N__19457),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24126),
            .lcout(N_822_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un30_3_0_o2_1_LC_20_18_2 .C_ON=1'b0;
    defparam \this_start_data_delay.un30_3_0_o2_1_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un30_3_0_o2_1_LC_20_18_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_start_data_delay.un30_3_0_o2_1_LC_20_18_2  (
            .in0(N__23958),
            .in1(N__21089),
            .in2(_gnd_net_),
            .in3(N__21321),
            .lcout(),
            .ltout(\this_start_data_delay.N_844_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIEFRT1_LC_20_18_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIEFRT1_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIEFRT1_LC_20_18_3 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \this_start_data_delay.M_last_q_RNIEFRT1_LC_20_18_3  (
            .in0(N__23490),
            .in1(N__22163),
            .in2(N__19437),
            .in3(N__24125),
            .lcout(\this_start_data_delay.N_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un1_M_this_substate_q4_2_i_0_303_i_a2_i_a2_LC_20_18_4 .C_ON=1'b0;
    defparam \this_start_data_delay.un1_M_this_substate_q4_2_i_0_303_i_a2_i_a2_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un1_M_this_substate_q4_2_i_0_303_i_a2_i_a2_LC_20_18_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_start_data_delay.un1_M_this_substate_q4_2_i_0_303_i_a2_i_a2_LC_20_18_4  (
            .in0(N__19423),
            .in1(N__19723),
            .in2(_gnd_net_),
            .in3(N__23491),
            .lcout(\this_start_data_delay.N_151 ),
            .ltout(\this_start_data_delay.N_151_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un1_M_this_substate_q4_2_i_0_303_i_a2_i_i_LC_20_18_5 .C_ON=1'b0;
    defparam \this_start_data_delay.un1_M_this_substate_q4_2_i_0_303_i_a2_i_i_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un1_M_this_substate_q4_2_i_0_303_i_a2_i_i_LC_20_18_5 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \this_start_data_delay.un1_M_this_substate_q4_2_i_0_303_i_a2_i_i_LC_20_18_5  (
            .in0(N__26183),
            .in1(_gnd_net_),
            .in2(N__19434),
            .in3(N__26867),
            .lcout(N_33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIOU691_LC_20_18_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIOU691_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIOU691_LC_20_18_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIOU691_LC_20_18_6  (
            .in0(N__24127),
            .in1(N__24309),
            .in2(_gnd_net_),
            .in3(N__26182),
            .lcout(N_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_o2_LC_20_18_7 .C_ON=1'b0;
    defparam \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_o2_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_o2_LC_20_18_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_o2_LC_20_18_7  (
            .in0(_gnd_net_),
            .in1(N__19422),
            .in2(_gnd_net_),
            .in3(N__19399),
            .lcout(\this_start_data_delay.N_93_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_0_LC_20_19_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_0_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_0_LC_20_19_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIK0EI1_0_LC_20_19_0  (
            .in0(N__19624),
            .in1(N__19559),
            .in2(N__19706),
            .in3(N__19488),
            .lcout(\this_start_data_delay.N_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIOVDB1_LC_20_19_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIOVDB1_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIOVDB1_LC_20_19_2 .LUT_INIT=16'b0011111000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIOVDB1_LC_20_19_2  (
            .in0(N__19625),
            .in1(N__19560),
            .in2(N__19707),
            .in3(N__19968),
            .lcout(),
            .ltout(\this_start_data_delay.N_909_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_0_LC_20_19_3.C_ON=1'b0;
    defparam M_this_state_q_0_LC_20_19_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_0_LC_20_19_3.LUT_INIT=16'b1111111100111011;
    LogicCell40 M_this_state_q_0_LC_20_19_3 (
            .in0(N__19934),
            .in1(N__19905),
            .in2(N__19956),
            .in3(N__26212),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32586),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI3F19A_LC_20_19_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI3F19A_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI3F19A_LC_20_19_5 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \this_start_data_delay.M_last_q_RNI3F19A_LC_20_19_5  (
            .in0(N__19727),
            .in1(N__19914),
            .in2(N__21117),
            .in3(N__26875),
            .lcout(\this_start_data_delay.M_this_state_q_ns_0_i_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIA89G3_0_LC_20_19_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIA89G3_0_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIA89G3_0_LC_20_19_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIA89G3_0_LC_20_19_6  (
            .in0(_gnd_net_),
            .in1(N__19756),
            .in2(_gnd_net_),
            .in3(N__23664),
            .lcout(),
            .ltout(\this_start_data_delay.N_910_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_10_LC_20_19_7.C_ON=1'b0;
    defparam M_this_state_q_10_LC_20_19_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_10_LC_20_19_7.LUT_INIT=16'b0000000011111110;
    LogicCell40 M_this_state_q_10_LC_20_19_7 (
            .in0(N__24040),
            .in1(N__19794),
            .in2(N__19767),
            .in3(N__26213),
            .lcout(M_this_state_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32586),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIDHST1_LC_20_20_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIDHST1_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIDHST1_LC_20_20_1 .LUT_INIT=16'b0010001100000001;
    LogicCell40 \this_start_data_delay.M_last_q_RNIDHST1_LC_20_20_1  (
            .in0(N__24308),
            .in1(N__23776),
            .in2(N__19731),
            .in3(N__24221),
            .lcout(\this_start_data_delay.M_this_data_count_qlde_i_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_1_LC_20_20_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_1_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIK0EI1_1_LC_20_20_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIK0EI1_1_LC_20_20_3  (
            .in0(N__19696),
            .in1(N__19629),
            .in2(N__19567),
            .in3(N__19489),
            .lcout(\this_start_data_delay.N_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_2_LC_20_20_4.C_ON=1'b0;
    defparam M_this_state_q_2_LC_20_20_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_20_20_4.LUT_INIT=16'b0011000100110000;
    LogicCell40 M_this_state_q_2_LC_20_20_4 (
            .in0(N__24222),
            .in1(N__26209),
            .in2(N__19470),
            .in3(N__21088),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32592),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_6_LC_20_20_6.C_ON=1'b0;
    defparam M_this_state_q_6_LC_20_20_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_20_20_6.LUT_INIT=16'b0000000011011100;
    LogicCell40 M_this_state_q_6_LC_20_20_6 (
            .in0(N__24223),
            .in1(N__19998),
            .in2(N__23795),
            .in3(N__26210),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32592),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_20_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_20_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_20_20_7 .LUT_INIT=16'b1011111111111101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_22_LC_20_20_7  (
            .in0(N__21871),
            .in1(N__20237),
            .in2(N__22316),
            .in3(N__22533),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_20_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_20_21_0 .LUT_INIT=16'b1101111111111011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_23_LC_20_21_0  (
            .in0(N__20238),
            .in1(N__21862),
            .in2(N__22327),
            .in3(N__21948),
            .lcout(\this_vga_signals.N_4558_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_20_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_20_21_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_20_21_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_20_21_1  (
            .in0(N__23429),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32601),
            .ce(N__23401),
            .sr(N__23314));
    defparam \this_vga_signals.un5_vaddress_g0_4_i_a3_1_0_LC_20_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_i_a3_1_0_LC_20_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_i_a3_1_0_LC_20_21_2 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_i_a3_1_0_LC_20_21_2  (
            .in0(N__22531),
            .in1(N__21860),
            .in2(N__20088),
            .in3(N__21946),
            .lcout(),
            .ltout(\this_vga_signals.g0_4_i_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_i_1_LC_20_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_i_1_LC_20_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_i_1_LC_20_21_3 .LUT_INIT=16'b0100011111001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_i_1_LC_20_21_3  (
            .in0(N__19974),
            .in1(N__20239),
            .in2(N__19980),
            .in3(N__20083),
            .lcout(),
            .ltout(\this_vga_signals.g0_4_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_i_LC_20_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_i_LC_20_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_i_LC_20_21_4 .LUT_INIT=16'b0010111101001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_i_LC_20_21_4  (
            .in0(N__22532),
            .in1(N__21861),
            .in2(N__19977),
            .in3(N__21947),
            .lcout(\this_vga_signals.N_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_i_o3_1_LC_20_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_i_o3_1_LC_20_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_i_o3_1_LC_20_21_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_i_o3_1_LC_20_21_5  (
            .in0(N__21776),
            .in1(N__21813),
            .in2(_gnd_net_),
            .in3(N__22530),
            .lcout(\this_vga_signals.N_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_20_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_20_21_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_20_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_20_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23428),
            .lcout(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32601),
            .ce(N__23401),
            .sr(N__23314));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_x0_LC_20_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_x0_LC_20_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_x0_LC_20_21_7 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_x0_LC_20_21_7  (
            .in0(_gnd_net_),
            .in1(N__21768),
            .in2(N__20085),
            .in3(N__21812),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_602_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_20_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_20_22_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_20_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_20_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21389),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32610),
            .ce(N__23408),
            .sr(N__23316));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_20_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_20_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_20_22_1 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_20_22_1  (
            .in0(N__21770),
            .in1(N__20248),
            .in2(N__20147),
            .in3(N__20071),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_4_LC_20_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_4_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_4_LC_20_22_2 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_4_LC_20_22_2  (
            .in0(N__20026),
            .in1(N__20124),
            .in2(_gnd_net_),
            .in3(N__21691),
            .lcout(\this_vga_signals.r_N_4_mux ),
            .ltout(\this_vga_signals.r_N_4_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIEC471_LC_20_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIEC471_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIEC471_LC_20_22_3 .LUT_INIT=16'b1000101011100111;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIEC471_LC_20_22_3  (
            .in0(N__21811),
            .in1(N__21774),
            .in2(N__20154),
            .in3(N__22501),
            .lcout(\this_vga_signals.SUM_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_x1_LC_20_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_x1_LC_20_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_x1_LC_20_22_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_x1_LC_20_22_4  (
            .in0(N__20027),
            .in1(N__21810),
            .in2(N__22536),
            .in3(N__21692),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_ns_LC_20_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_ns_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_ns_LC_20_22_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_ns_LC_20_22_5  (
            .in0(N__20125),
            .in1(_gnd_net_),
            .in2(N__20103),
            .in3(N__20094),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a1_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_x0_LC_20_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_x0_LC_20_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_x0_LC_20_22_6 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_x0_LC_20_22_6  (
            .in0(_gnd_net_),
            .in1(N__21690),
            .in2(N__22535),
            .in3(N__21806),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_x1_LC_20_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_x1_LC_20_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_x1_LC_20_22_7 .LUT_INIT=16'b1111011111101111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_x1_LC_20_22_7  (
            .in0(N__21769),
            .in1(N__20070),
            .in2(N__21818),
            .in3(N__20025),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_602_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_3_x1_LC_20_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_3_x1_LC_20_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_3_x1_LC_20_23_0 .LUT_INIT=16'b1000100000001000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_3_x1_LC_20_23_0  (
            .in0(N__22537),
            .in1(N__21693),
            .in2(N__22044),
            .in3(N__23415),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_0_3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_1_LC_20_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_1_LC_20_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_1_LC_20_23_1 .LUT_INIT=16'b0101011010101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_1_LC_20_23_1  (
            .in0(N__22352),
            .in1(N__22997),
            .in2(N__23250),
            .in3(N__20687),
            .lcout(),
            .ltout(\this_vga_signals.g0_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_20_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_20_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_20_23_2 .LUT_INIT=16'b0111100011010010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_26_LC_20_23_2  (
            .in0(N__22998),
            .in1(N__23213),
            .in2(N__20670),
            .in3(N__20662),
            .lcout(\this_vga_signals.N_4_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_5_LC_20_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_5_LC_20_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_5_LC_20_23_3 .LUT_INIT=16'b1010010101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_5_LC_20_23_3  (
            .in0(N__22351),
            .in1(_gnd_net_),
            .in2(N__23249),
            .in3(N__22996),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_20_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_20_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_20_23_4 .LUT_INIT=16'b1000001111001011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_LC_20_23_4  (
            .in0(N__20601),
            .in1(N__20341),
            .in2(N__20592),
            .in3(N__20418),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_20_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_20_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_20_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_20_23_5  (
            .in0(_gnd_net_),
            .in1(N__20551),
            .in2(_gnd_net_),
            .in3(N__20508),
            .lcout(\this_vga_signals.vaddress_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_20_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_20_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_20_23_6 .LUT_INIT=16'b0000011011100111;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_1_LC_20_23_6  (
            .in0(N__22999),
            .in1(N__23214),
            .in2(N__22404),
            .in3(N__20419),
            .lcout(),
            .ltout(\this_vga_signals.g2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_LC_20_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_LC_20_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_LC_20_23_7 .LUT_INIT=16'b0100111010110001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_LC_20_23_7  (
            .in0(N__20342),
            .in1(N__20961),
            .in2(N__20301),
            .in3(N__20298),
            .lcout(\this_vga_signals.g0_i_x4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_1_LC_20_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_1_LC_20_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_1_LC_20_24_3 .LUT_INIT=16'b1010100101010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_0_a3_1_LC_20_24_3  (
            .in0(N__22841),
            .in1(N__23200),
            .in2(N__23093),
            .in3(N__22673),
            .lcout(\this_vga_signals.g0_3_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_5_LC_20_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_5_LC_20_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_5_LC_20_24_5 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_5_LC_20_24_5  (
            .in0(N__23073),
            .in1(N__23199),
            .in2(_gnd_net_),
            .in3(N__22356),
            .lcout(\this_vga_signals.vaddress_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIBR6R_1_LC_20_31_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIBR6R_1_LC_20_31_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIBR6R_1_LC_20_31_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \this_ppu.M_haddress_q_RNIBR6R_1_LC_20_31_4  (
            .in0(N__32102),
            .in1(N__20955),
            .in2(N__31934),
            .in3(N__20933),
            .lcout(M_this_ppu_sprites_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_21_11_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_21_11_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_21_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_21_11_6  (
            .in0(N__30106),
            .in1(N__20775),
            .in2(_gnd_net_),
            .in3(N__20760),
            .lcout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_4_LC_21_15_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_4_LC_21_15_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_4_LC_21_15_4.LUT_INIT=16'b0101110111010101;
    LogicCell40 M_this_sprites_address_q_4_LC_21_15_4 (
            .in0(N__21045),
            .in1(N__27517),
            .in2(N__24744),
            .in3(N__24708),
            .lcout(M_this_sprites_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32557),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIK6R81_LC_21_16_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIK6R81_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIK6R81_LC_21_16_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_start_data_delay.M_last_q_RNIK6R81_LC_21_16_2  (
            .in0(N__23472),
            .in1(N__23947),
            .in2(_gnd_net_),
            .in3(N__24164),
            .lcout(M_this_sprites_ram_write_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNICA9G3_LC_21_16_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNICA9G3_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNICA9G3_LC_21_16_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_start_data_delay.M_last_q_RNICA9G3_LC_21_16_4  (
            .in0(N__23731),
            .in1(N__20742),
            .in2(_gnd_net_),
            .in3(N__26876),
            .lcout(\this_start_data_delay.N_125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIOCPV6_0_LC_21_16_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIOCPV6_0_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIOCPV6_0_LC_21_16_6 .LUT_INIT=16'b0000111110111111;
    LogicCell40 \this_start_data_delay.M_last_q_RNIOCPV6_0_LC_21_16_6  (
            .in0(N__23799),
            .in1(N__23532),
            .in2(N__23577),
            .in3(N__24609),
            .lcout(),
            .ltout(\this_start_data_delay.un30_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNINS0N8_LC_21_16_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNINS0N8_LC_21_16_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNINS0N8_LC_21_16_7 .LUT_INIT=16'b0000000011110011;
    LogicCell40 \this_start_data_delay.M_last_q_RNINS0N8_LC_21_16_7  (
            .in0(_gnd_net_),
            .in1(N__27822),
            .in2(N__20700),
            .in3(N__26199),
            .lcout(\this_start_data_delay.N_990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIHV2L3_LC_21_17_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIHV2L3_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIHV2L3_LC_21_17_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \this_start_data_delay.M_last_q_RNIHV2L3_LC_21_17_0  (
            .in0(N__30573),
            .in1(N__28302),
            .in2(N__27658),
            .in3(N__27603),
            .lcout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_21_17_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_21_17_1 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_21_17_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_21_17_1  (
            .in0(N__20979),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21009),
            .lcout(\this_start_data_delay.M_last_qZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32576),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_0_LC_21_17_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_0_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_0_LC_21_17_2 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBJQQ_0_LC_21_17_2  (
            .in0(N__21010),
            .in1(N__21025),
            .in2(_gnd_net_),
            .in3(N__20978),
            .lcout(N_554_0),
            .ltout(N_554_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIIT6G1_LC_21_17_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIIT6G1_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIIT6G1_LC_21_17_3 .LUT_INIT=16'b0100010101000100;
    LogicCell40 \this_start_data_delay.M_last_q_RNIIT6G1_LC_21_17_3  (
            .in0(N__26185),
            .in1(N__21101),
            .in2(N__21108),
            .in3(N__21323),
            .lcout(\this_start_data_delay.N_992 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIIT6G1_0_LC_21_17_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIIT6G1_0_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIIT6G1_0_LC_21_17_4 .LUT_INIT=16'b0010001000110010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIIT6G1_0_LC_21_17_4  (
            .in0(N__21324),
            .in1(N__26186),
            .in2(N__21105),
            .in3(N__24161),
            .lcout(\this_start_data_delay.N_109 ),
            .ltout(\this_start_data_delay.N_109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI433C3_LC_21_17_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI433C3_LC_21_17_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI433C3_LC_21_17_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \this_start_data_delay.M_last_q_RNI433C3_LC_21_17_5  (
            .in0(N__28301),
            .in1(N__24745),
            .in2(N__21048),
            .in3(N__25330),
            .lcout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBOQ11_LC_21_18_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBOQ11_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBOQ11_LC_21_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBOQ11_LC_21_18_0  (
            .in0(_gnd_net_),
            .in1(N__21272),
            .in2(_gnd_net_),
            .in3(N__24128),
            .lcout(\this_start_data_delay.N_86_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_21_18_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_21_18_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBJQQ_LC_21_18_1  (
            .in0(N__21027),
            .in1(N__21011),
            .in2(_gnd_net_),
            .in3(N__20977),
            .lcout(\this_start_data_delay.N_555_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_21_18_2 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_21_18_2 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_21_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_21_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21036),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32587),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIDQQ11_LC_21_18_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIDQQ11_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIDQQ11_LC_21_18_3 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIDQQ11_LC_21_18_3  (
            .in0(N__21026),
            .in1(N__21012),
            .in2(N__23798),
            .in3(N__20976),
            .lcout(\this_start_data_delay.N_91_0 ),
            .ltout(\this_start_data_delay.N_91_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI12SC4_0_LC_21_18_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI12SC4_0_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI12SC4_0_LC_21_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI12SC4_0_LC_21_18_4  (
            .in0(N__28032),
            .in1(N__24474),
            .in2(N__21327),
            .in3(N__32874),
            .lcout(N_116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIKQ691_LC_21_18_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIKQ691_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIKQ691_LC_21_18_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIKQ691_LC_21_18_5  (
            .in0(N__24129),
            .in1(N__26184),
            .in2(_gnd_net_),
            .in3(N__21322),
            .lcout(\this_start_data_delay.N_110 ),
            .ltout(\this_start_data_delay.N_110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI653C3_0_LC_21_18_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI653C3_0_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI653C3_0_LC_21_18_6 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \this_start_data_delay.M_last_q_RNI653C3_0_LC_21_18_6  (
            .in0(N__26308),
            .in1(N__32875),
            .in2(N__21279),
            .in3(N__27645),
            .lcout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI6UUI2_LC_21_18_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI6UUI2_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI6UUI2_LC_21_18_7 .LUT_INIT=16'b0000000010100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNI6UUI2_LC_21_18_7  (
            .in0(N__24130),
            .in1(N__24680),
            .in2(N__21276),
            .in3(N__23791),
            .lcout(\this_start_data_delay.N_121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_21_19_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_21_19_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_21_19_0  (
            .in0(N__21249),
            .in1(N__21237),
            .in2(_gnd_net_),
            .in3(N__30036),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_19_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_19_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_19_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_19_1  (
            .in0(N__30035),
            .in1(N__21219),
            .in2(_gnd_net_),
            .in3(N__21204),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_21_19_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_21_19_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_21_19_2 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_21_19_2  (
            .in0(N__28727),
            .in1(N__28668),
            .in2(N__21186),
            .in3(N__21183),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_21_19_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_21_19_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_21_19_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_21_19_3  (
            .in0(N__28669),
            .in1(N__23583),
            .in2(N__21171),
            .in3(N__21168),
            .lcout(M_this_ppu_vram_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI12SC4_1_LC_21_19_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI12SC4_1_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI12SC4_1_LC_21_19_4 .LUT_INIT=16'b0011101100000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI12SC4_1_LC_21_19_4  (
            .in0(N__32892),
            .in1(N__28036),
            .in2(N__24473),
            .in3(N__23827),
            .lcout(\this_start_data_delay.M_this_state_q_ns_0_i_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_21_20_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_21_20_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_21_20_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_21_20_0  (
            .in0(N__21537),
            .in1(N__21568),
            .in2(N__21675),
            .in3(N__21674),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_21_20_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__32602),
            .ce(),
            .sr(N__23311));
    defparam \this_vga_signals.M_vcounter_q_1_LC_21_20_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_21_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_21_20_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_21_20_1  (
            .in0(N__21539),
            .in1(N__22898),
            .in2(_gnd_net_),
            .in3(N__21546),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__32602),
            .ce(),
            .sr(N__23311));
    defparam \this_vga_signals.M_vcounter_q_2_LC_21_20_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_21_20_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_21_20_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_21_20_2  (
            .in0(N__21538),
            .in1(N__22648),
            .in2(_gnd_net_),
            .in3(N__21543),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__32602),
            .ce(),
            .sr(N__23311));
    defparam \this_vga_signals.M_vcounter_q_3_LC_21_20_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_21_20_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_21_20_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_21_20_3  (
            .in0(N__21540),
            .in1(N__22771),
            .in2(_gnd_net_),
            .in3(N__21393),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__32602),
            .ce(),
            .sr(N__23311));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_21_20_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_21_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_21_20_4  (
            .in0(_gnd_net_),
            .in1(N__23285),
            .in2(_gnd_net_),
            .in3(N__21357),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_21_20_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_21_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_21_20_5  (
            .in0(_gnd_net_),
            .in1(N__23088),
            .in2(_gnd_net_),
            .in3(N__21336),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_21_20_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_21_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_21_20_6  (
            .in0(_gnd_net_),
            .in1(N__22320),
            .in2(_gnd_net_),
            .in3(N__21333),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_21_20_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_21_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_21_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_21_20_7  (
            .in0(_gnd_net_),
            .in1(N__21967),
            .in2(_gnd_net_),
            .in3(N__21330),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_21_21_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_21_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_21_21_0  (
            .in0(_gnd_net_),
            .in1(N__21882),
            .in2(_gnd_net_),
            .in3(N__22050),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_21_21_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_21_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_21_21_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_21_21_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_21_21_1  (
            .in0(_gnd_net_),
            .in1(N__22534),
            .in2(_gnd_net_),
            .in3(N__22047),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32611),
            .ce(N__23402),
            .sr(N__23312));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_21_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_21_21_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_21_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_21_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22031),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32611),
            .ce(N__23402),
            .sr(N__23312));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_21_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_21_21_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_21_21_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_21_21_3  (
            .in0(N__22032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32611),
            .ce(N__23402),
            .sr(N__23312));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_21_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_21_21_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_21_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_21_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22030),
            .lcout(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32611),
            .ce(N__23402),
            .sr(N__23312));
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_21_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_21_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_21_22_5 .LUT_INIT=16'b1011101111011101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_17_LC_21_22_5  (
            .in0(N__21872),
            .in1(N__21962),
            .in2(_gnd_net_),
            .in3(N__22503),
            .lcout(\this_vga_signals.N_4557_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_8_LC_21_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_8_LC_21_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_8_LC_21_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIROQM_8_LC_21_22_6  (
            .in0(N__21963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21873),
            .lcout(\this_vga_signals.m58_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_601_LC_21_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_601_LC_21_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_601_LC_21_22_7 .LUT_INIT=16'b1100111111110011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_601_LC_21_22_7  (
            .in0(_gnd_net_),
            .in1(N__21814),
            .in2(N__21777),
            .in3(N__22502),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_21_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_21_23_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_21_23_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_21_23_0  (
            .in0(_gnd_net_),
            .in1(N__21719),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32625),
            .ce(N__23406),
            .sr(N__23317));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_21_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_21_23_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_21_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_21_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23433),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32625),
            .ce(N__23406),
            .sr(N__23317));
    defparam \this_start_data_delay.M_last_q_RNI75F36_LC_21_24_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI75F36_LC_21_24_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI75F36_LC_21_24_0 .LUT_INIT=16'b1111111100011101;
    LogicCell40 \this_start_data_delay.M_last_q_RNI75F36_LC_21_24_0  (
            .in0(N__26755),
            .in1(N__26271),
            .in2(N__28275),
            .in3(N__26194),
            .lcout(M_this_external_address_q_3_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI97F36_LC_21_24_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI97F36_LC_21_24_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI97F36_LC_21_24_2 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNI97F36_LC_21_24_2  (
            .in0(N__23999),
            .in1(N__26272),
            .in2(N__28166),
            .in3(N__26195),
            .lcout(M_this_external_address_q_3_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_21_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_21_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_21_24_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_21_24_5  (
            .in0(N__23276),
            .in1(N__23089),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.m58_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNICVQL1_1_LC_21_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNICVQL1_1_LC_21_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNICVQL1_1_LC_21_24_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNICVQL1_1_LC_21_24_6  (
            .in0(N__22915),
            .in1(N__22842),
            .in2(N__22709),
            .in3(N__22569),
            .lcout(),
            .ltout(\this_vga_signals.m58_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_21_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_21_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_21_24_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_21_24_7  (
            .in0(N__22433),
            .in1(N__22413),
            .in2(N__22407),
            .in3(N__22360),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI12SC4_2_LC_21_25_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI12SC4_2_LC_21_25_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI12SC4_2_LC_21_25_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI12SC4_2_LC_21_25_4  (
            .in0(N__32800),
            .in1(N__24503),
            .in2(N__28044),
            .in3(N__23832),
            .lcout(N_911),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIJARF1_LC_22_15_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIJARF1_LC_22_15_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIJARF1_LC_22_15_6 .LUT_INIT=16'b0000000100110011;
    LogicCell40 \this_start_data_delay.M_last_q_RNIJARF1_LC_22_15_6  (
            .in0(N__22179),
            .in1(N__23954),
            .in2(N__23495),
            .in3(N__24204),
            .lcout(\this_start_data_delay.N_123 ),
            .ltout(\this_start_data_delay.N_123_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIUFEC3_LC_22_15_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIUFEC3_LC_22_15_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIUFEC3_LC_22_15_7 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIUFEC3_LC_22_15_7  (
            .in0(N__30935),
            .in1(N__24488),
            .in2(N__22137),
            .in3(N__27979),
            .lcout(N_812_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_7_LC_22_16_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_7_LC_22_16_0.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_7_LC_22_16_0.LUT_INIT=16'b0101110111010101;
    LogicCell40 M_this_sprites_address_q_7_LC_22_16_0 (
            .in0(N__23508),
            .in1(N__27518),
            .in2(N__25589),
            .in3(N__25554),
            .lcout(M_this_sprites_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32577),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI213C3_0_LC_22_16_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI213C3_0_LC_22_16_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI213C3_0_LC_22_16_7 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \this_start_data_delay.M_last_q_RNI213C3_0_LC_22_16_7  (
            .in0(N__27646),
            .in1(N__28471),
            .in2(N__25588),
            .in3(N__27611),
            .lcout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI12SC4_3_LC_22_17_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI12SC4_3_LC_22_17_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI12SC4_3_LC_22_17_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI12SC4_3_LC_22_17_0  (
            .in0(N__28014),
            .in1(N__32891),
            .in2(N__24487),
            .in3(N__23820),
            .lcout(\this_start_data_delay.N_938_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI0T8G3_LC_22_17_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI0T8G3_LC_22_17_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI0T8G3_LC_22_17_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI0T8G3_LC_22_17_1  (
            .in0(N__23901),
            .in1(N__23726),
            .in2(_gnd_net_),
            .in3(N__26871),
            .lcout(),
            .ltout(\this_start_data_delay.N_129_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_8_LC_22_17_2.C_ON=1'b0;
    defparam M_this_state_q_8_LC_22_17_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_8_LC_22_17_2.LUT_INIT=16'b0000000011110100;
    LogicCell40 M_this_state_q_8_LC_22_17_2 (
            .in0(N__24163),
            .in1(N__23474),
            .in2(N__23502),
            .in3(N__26223),
            .lcout(M_this_state_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32588),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIJ13L3_LC_22_17_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIJ13L3_LC_22_17_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIJ13L3_LC_22_17_3 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \this_start_data_delay.M_last_q_RNIJ13L3_LC_22_17_3  (
            .in0(N__27607),
            .in1(N__24458),
            .in2(N__30677),
            .in3(N__27657),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_12_LC_22_17_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_12_LC_22_17_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_12_LC_22_17_4.LUT_INIT=16'b0010111110001111;
    LogicCell40 M_this_sprites_address_q_12_LC_22_17_4 (
            .in0(N__27533),
            .in1(N__30657),
            .in2(N__23499),
            .in3(N__25395),
            .lcout(M_this_sprites_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32588),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIFSQ11_LC_22_17_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIFSQ11_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIFSQ11_LC_22_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIFSQ11_LC_22_17_5  (
            .in0(_gnd_net_),
            .in1(N__23473),
            .in2(_gnd_net_),
            .in3(N__24162),
            .lcout(\this_start_data_delay.N_821_0 ),
            .ltout(\this_start_data_delay.N_821_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_9_LC_22_17_6.C_ON=1'b0;
    defparam M_this_state_q_9_LC_22_17_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_9_LC_22_17_6.LUT_INIT=16'b0000000011110000;
    LogicCell40 M_this_state_q_9_LC_22_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23436),
            .in3(N__26224),
            .lcout(M_this_state_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32588),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_11_LC_22_17_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_11_LC_22_17_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_11_LC_22_17_7.LUT_INIT=16'b0101110111010101;
    LogicCell40 M_this_sprites_address_q_11_LC_22_17_7 (
            .in0(N__23625),
            .in1(N__27532),
            .in2(N__30592),
            .in3(N__25404),
            .lcout(M_this_sprites_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32588),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIFT2L3_LC_22_18_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIFT2L3_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIFT2L3_LC_22_18_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \this_start_data_delay.M_last_q_RNIFT2L3_LC_22_18_0  (
            .in0(N__27602),
            .in1(N__25435),
            .in2(N__31342),
            .in3(N__27653),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_10_LC_22_18_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_10_LC_22_18_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_10_LC_22_18_1.LUT_INIT=16'b0100111110001111;
    LogicCell40 M_this_sprites_address_q_10_LC_22_18_1 (
            .in0(N__25434),
            .in1(N__27557),
            .in2(N__23619),
            .in3(N__25413),
            .lcout(M_this_sprites_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32593),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_22_18_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_22_18_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_22_18_2  (
            .in0(N__23616),
            .in1(N__23598),
            .in2(_gnd_net_),
            .in3(N__30056),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIL33L3_LC_22_18_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIL33L3_LC_22_18_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIL33L3_LC_22_18_3 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \this_start_data_delay.M_last_q_RNIL33L3_LC_22_18_3  (
            .in0(N__30480),
            .in1(N__28127),
            .in2(N__27659),
            .in3(N__27601),
            .lcout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIOCPV6_LC_22_18_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIOCPV6_LC_22_18_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIOCPV6_LC_22_18_7 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIOCPV6_LC_22_18_7  (
            .in0(N__23796),
            .in1(N__24608),
            .in2(N__23572),
            .in3(N__23531),
            .lcout(un30_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI0V2C3_LC_22_19_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI0V2C3_LC_22_19_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI0V2C3_LC_22_19_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \this_start_data_delay.M_last_q_RNI0V2C3_LC_22_19_0  (
            .in0(N__25033),
            .in1(N__25300),
            .in2(N__32903),
            .in3(N__25352),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_2_LC_22_19_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_2_LC_22_19_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_2_LC_22_19_1.LUT_INIT=16'b0100111110001111;
    LogicCell40 M_this_sprites_address_q_2_LC_22_19_1 (
            .in0(N__25032),
            .in1(N__27558),
            .in2(N__23514),
            .in3(N__25008),
            .lcout(M_this_sprites_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32603),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI0T8G3_0_LC_22_19_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI0T8G3_0_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI0T8G3_0_LC_22_19_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI0T8G3_0_LC_22_19_2  (
            .in0(_gnd_net_),
            .in1(N__23889),
            .in2(_gnd_net_),
            .in3(N__23652),
            .lcout(),
            .ltout(\this_start_data_delay.N_913_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_22_19_3.C_ON=1'b0;
    defparam M_this_state_q_7_LC_22_19_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_22_19_3.LUT_INIT=16'b0101010101010100;
    LogicCell40 M_this_state_q_7_LC_22_19_3 (
            .in0(N__26222),
            .in1(N__24622),
            .in2(N__23511),
            .in3(N__23957),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32603),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI213C3_LC_22_19_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI213C3_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI213C3_LC_22_19_4 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \this_start_data_delay.M_last_q_RNI213C3_LC_22_19_4  (
            .in0(N__24889),
            .in1(N__25301),
            .in2(N__31355),
            .in3(N__25353),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_3_LC_22_19_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_3_LC_22_19_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_3_LC_22_19_5.LUT_INIT=16'b0100111110001111;
    LogicCell40 M_this_sprites_address_q_3_LC_22_19_5 (
            .in0(N__24888),
            .in1(N__27559),
            .in2(N__23868),
            .in3(N__24864),
            .lcout(M_this_sprites_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32603),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_13_LC_22_19_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_13_LC_22_19_6 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_13_LC_22_19_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \this_sprites_ram.mem_radreg_13_LC_22_19_6  (
            .in0(N__31919),
            .in1(N__32141),
            .in2(N__23865),
            .in3(N__23841),
            .lcout(\this_sprites_ram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32603),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI12SC4_LC_22_20_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI12SC4_LC_22_20_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI12SC4_LC_22_20_0 .LUT_INIT=16'b1101000000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI12SC4_LC_22_20_0  (
            .in0(N__32858),
            .in1(N__24445),
            .in2(N__28040),
            .in3(N__23828),
            .lcout(\this_start_data_delay.N_149 ),
            .ltout(\this_start_data_delay.N_149_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIF2NL5_LC_22_20_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIF2NL5_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIF2NL5_LC_22_20_1 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \this_start_data_delay.M_last_q_RNIF2NL5_LC_22_20_1  (
            .in0(N__24281),
            .in1(N__24178),
            .in2(N__23802),
            .in3(N__23797),
            .lcout(\this_start_data_delay.M_this_data_count_qlde_i_2_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNITK893_LC_22_20_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNITK893_LC_22_20_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNITK893_LC_22_20_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_start_data_delay.M_last_q_RNITK893_LC_22_20_3  (
            .in0(_gnd_net_),
            .in1(N__23732),
            .in2(_gnd_net_),
            .in3(N__26851),
            .lcout(\this_start_data_delay.N_820_0 ),
            .ltout(\this_start_data_delay.N_820_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI281SC_LC_22_20_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI281SC_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI281SC_LC_22_20_4 .LUT_INIT=16'b1100010011110101;
    LogicCell40 \this_start_data_delay.M_last_q_RNI281SC_LC_22_20_4  (
            .in0(N__23694),
            .in1(N__23685),
            .in2(N__23679),
            .in3(N__23676),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_data_count_qlde_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIC4IPK_LC_22_20_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIC4IPK_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIC4IPK_LC_22_20_5 .LUT_INIT=16'b1111111100101111;
    LogicCell40 \this_start_data_delay.M_last_q_RNIC4IPK_LC_22_20_5  (
            .in0(N__24647),
            .in1(N__23656),
            .in2(N__23628),
            .in3(N__26201),
            .lcout(N_35),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_5_LC_22_20_7.C_ON=1'b0;
    defparam M_this_state_q_5_LC_22_20_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_22_20_7.LUT_INIT=16'b0000000010111010;
    LogicCell40 M_this_state_q_5_LC_22_20_7 (
            .in0(N__24327),
            .in1(N__24179),
            .in2(N__24301),
            .in3(N__26202),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32612),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_d62_11_LC_22_21_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d62_11_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d62_11_LC_22_21_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.M_this_state_d62_11_LC_22_21_1  (
            .in0(N__28910),
            .in1(N__28939),
            .in2(N__28886),
            .in3(N__29136),
            .lcout(\this_start_data_delay.M_this_state_d62Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_5_LC_22_21_3.C_ON=1'b0;
    defparam M_this_data_count_q_5_LC_22_21_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_22_21_3.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_5_LC_22_21_3 (
            .in0(N__29195),
            .in1(N__28926),
            .in2(_gnd_net_),
            .in3(N__28940),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32618),
            .ce(N__29104),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_7_LC_22_21_4.C_ON=1'b0;
    defparam M_this_data_count_q_7_LC_22_21_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_22_21_4.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_7_LC_22_21_4 (
            .in0(N__28866),
            .in1(N__29196),
            .in2(_gnd_net_),
            .in3(N__28882),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32618),
            .ce(N__29104),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIOU691_0_LC_22_21_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIOU691_0_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIOU691_0_LC_22_21_5 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \this_start_data_delay.M_last_q_RNIOU691_0_LC_22_21_5  (
            .in0(N__24285),
            .in1(N__26198),
            .in2(_gnd_net_),
            .in3(N__24226),
            .lcout(),
            .ltout(this_start_data_delay_M_this_data_count_q_3_0_a3_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_6_LC_22_21_6.C_ON=1'b0;
    defparam M_this_data_count_q_6_LC_22_21_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_22_21_6.LUT_INIT=16'b1100000010101010;
    LogicCell40 M_this_data_count_q_6_LC_22_21_6 (
            .in0(N__28899),
            .in1(N__26765),
            .in2(N__24051),
            .in3(N__29194),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32618),
            .ce(N__29104),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNII9RA6_LC_22_21_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNII9RA6_LC_22_21_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNII9RA6_LC_22_21_7 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNII9RA6_LC_22_21_7  (
            .in0(N__24019),
            .in1(N__26971),
            .in2(N__32884),
            .in3(N__26197),
            .lcout(M_this_data_count_q_3_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_22_22_1.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_22_22_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_22_22_1.LUT_INIT=16'b0111001000100111;
    LogicCell40 M_this_data_count_q_13_LC_22_22_1 (
            .in0(N__29235),
            .in1(N__23970),
            .in2(N__29859),
            .in3(N__29879),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32626),
            .ce(N__29081),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_9_LC_22_22_2.C_ON=1'b0;
    defparam M_this_data_count_q_9_LC_22_22_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_22_22_2.LUT_INIT=16'b1100000010101010;
    LogicCell40 M_this_data_count_q_9_LC_22_22_2 (
            .in0(N__29979),
            .in1(N__26974),
            .in2(N__30914),
            .in3(N__29234),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32626),
            .ce(N__29081),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_8_LC_22_22_6.C_ON=1'b0;
    defparam M_this_data_count_q_8_LC_22_22_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_22_22_6.LUT_INIT=16'b1100000010101010;
    LogicCell40 M_this_data_count_q_8_LC_22_22_6 (
            .in0(N__28833),
            .in1(N__26973),
            .in2(N__28470),
            .in3(N__29233),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32626),
            .ce(N__29081),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_i_LC_22_23_1 .C_ON=1'b0;
    defparam \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_i_LC_22_23_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_i_LC_22_23_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_i_LC_22_23_1  (
            .in0(_gnd_net_),
            .in1(N__26192),
            .in2(_gnd_net_),
            .in3(N__24690),
            .lcout(N_39),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIEGBV8_LC_22_23_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIEGBV8_LC_22_23_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIEGBV8_LC_22_23_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \this_start_data_delay.M_last_q_RNIEGBV8_LC_22_23_7  (
            .in0(N__24669),
            .in1(N__26193),
            .in2(N__24654),
            .in3(N__24636),
            .lcout(N_37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNINT691_LC_22_24_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNINT691_LC_22_24_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNINT691_LC_22_24_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_start_data_delay.M_last_q_RNINT691_LC_22_24_4  (
            .in0(_gnd_net_),
            .in1(N__26270),
            .in2(_gnd_net_),
            .in3(N__26190),
            .lcout(M_this_external_address_d_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI86F36_LC_22_24_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI86F36_LC_22_24_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI86F36_LC_22_24_5 .LUT_INIT=16'b1010111010111111;
    LogicCell40 \this_start_data_delay.M_last_q_RNI86F36_LC_22_24_5  (
            .in0(N__26191),
            .in1(N__26273),
            .in2(N__24498),
            .in3(N__24623),
            .lcout(M_this_external_address_q_3_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNISDEC3_LC_23_15_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNISDEC3_LC_23_15_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNISDEC3_LC_23_15_0 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNISDEC3_LC_23_15_0  (
            .in0(N__28419),
            .in1(N__27980),
            .in2(N__28320),
            .in3(N__27823),
            .lcout(N_813_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI653C3_LC_23_16_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI653C3_LC_23_16_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI653C3_LC_23_16_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \this_start_data_delay.M_last_q_RNI653C3_LC_23_16_0  (
            .in0(N__27069),
            .in1(N__25302),
            .in2(N__24497),
            .in3(N__25343),
            .lcout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI873C3_LC_23_16_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI873C3_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI873C3_LC_23_16_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \this_start_data_delay.M_last_q_RNI873C3_LC_23_16_1  (
            .in0(N__25345),
            .in1(N__28109),
            .in2(N__25313),
            .in3(N__25720),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_6_LC_23_16_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_6_LC_23_16_2.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_6_LC_23_16_2.LUT_INIT=16'b0100111110001111;
    LogicCell40 M_this_sprites_address_q_6_LC_23_16_2 (
            .in0(N__25719),
            .in1(N__27543),
            .in2(N__24330),
            .in3(N__25698),
            .lcout(M_this_sprites_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32589),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIUS2C3_LC_23_16_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIUS2C3_LC_23_16_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIUS2C3_LC_23_16_5 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \this_start_data_delay.M_last_q_RNIUS2C3_LC_23_16_5  (
            .in0(N__25346),
            .in1(N__30930),
            .in2(N__25314),
            .in3(N__25168),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_1_LC_23_16_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_1_LC_23_16_6.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_1_LC_23_16_6.LUT_INIT=16'b0110111100001111;
    LogicCell40 M_this_sprites_address_q_1_LC_23_16_6 (
            .in0(N__25167),
            .in1(N__25146),
            .in2(N__25356),
            .in3(N__27542),
            .lcout(M_this_sprites_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32589),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNISQ2C3_LC_23_16_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNISQ2C3_LC_23_16_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNISQ2C3_LC_23_16_7 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \this_start_data_delay.M_last_q_RNISQ2C3_LC_23_16_7  (
            .in0(N__25344),
            .in1(N__28472),
            .in2(N__25312),
            .in3(N__26457),
            .lcout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_0_c_LC_23_17_0.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_0_c_LC_23_17_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_0_c_LC_23_17_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_0_c_LC_23_17_0 (
            .in0(_gnd_net_),
            .in1(N__25367),
            .in2(N__26459),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_23_17_0_),
            .carryout(un1_M_this_sprites_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_0_THRU_LUT4_0_LC_23_17_1.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_0_THRU_LUT4_0_LC_23_17_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_0_THRU_LUT4_0_LC_23_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_0_THRU_LUT4_0_LC_23_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25175),
            .in3(N__25140),
            .lcout(un1_M_this_sprites_address_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_0),
            .carryout(un1_M_this_sprites_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_1_THRU_LUT4_0_LC_23_17_2.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_1_THRU_LUT4_0_LC_23_17_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_1_THRU_LUT4_0_LC_23_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_1_THRU_LUT4_0_LC_23_17_2 (
            .in0(_gnd_net_),
            .in1(N__25040),
            .in2(_gnd_net_),
            .in3(N__24999),
            .lcout(un1_M_this_sprites_address_q_cry_1_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_1),
            .carryout(un1_M_this_sprites_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_2_THRU_LUT4_0_LC_23_17_3.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_2_THRU_LUT4_0_LC_23_17_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_2_THRU_LUT4_0_LC_23_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_2_THRU_LUT4_0_LC_23_17_3 (
            .in0(_gnd_net_),
            .in1(N__24902),
            .in2(_gnd_net_),
            .in3(N__24855),
            .lcout(un1_M_this_sprites_address_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_2),
            .carryout(un1_M_this_sprites_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_3_THRU_LUT4_0_LC_23_17_4.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_3_THRU_LUT4_0_LC_23_17_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_3_THRU_LUT4_0_LC_23_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_3_THRU_LUT4_0_LC_23_17_4 (
            .in0(_gnd_net_),
            .in1(N__24752),
            .in2(_gnd_net_),
            .in3(N__24696),
            .lcout(un1_M_this_sprites_address_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_3),
            .carryout(un1_M_this_sprites_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_4_THRU_LUT4_0_LC_23_17_5.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_4_THRU_LUT4_0_LC_23_17_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_4_THRU_LUT4_0_LC_23_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_4_THRU_LUT4_0_LC_23_17_5 (
            .in0(_gnd_net_),
            .in1(N__27070),
            .in2(_gnd_net_),
            .in3(N__24693),
            .lcout(un1_M_this_sprites_address_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_4),
            .carryout(un1_M_this_sprites_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_5_THRU_LUT4_0_LC_23_17_6.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_5_THRU_LUT4_0_LC_23_17_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_5_THRU_LUT4_0_LC_23_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_5_THRU_LUT4_0_LC_23_17_6 (
            .in0(_gnd_net_),
            .in1(N__25721),
            .in2(_gnd_net_),
            .in3(N__25692),
            .lcout(un1_M_this_sprites_address_q_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_5),
            .carryout(un1_M_this_sprites_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_6_THRU_LUT4_0_LC_23_17_7.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_6_THRU_LUT4_0_LC_23_17_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_6_THRU_LUT4_0_LC_23_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_6_THRU_LUT4_0_LC_23_17_7 (
            .in0(_gnd_net_),
            .in1(N__25578),
            .in2(_gnd_net_),
            .in3(N__25548),
            .lcout(un1_M_this_sprites_address_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_6),
            .carryout(un1_M_this_sprites_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_7_THRU_LUT4_0_LC_23_18_0.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_7_THRU_LUT4_0_LC_23_18_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_7_THRU_LUT4_0_LC_23_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_7_THRU_LUT4_0_LC_23_18_0 (
            .in0(_gnd_net_),
            .in1(N__27380),
            .in2(_gnd_net_),
            .in3(N__25545),
            .lcout(un1_M_this_sprites_address_q_cry_7_THRU_CO),
            .ltout(),
            .carryin(bfn_23_18_0_),
            .carryout(un1_M_this_sprites_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_8_THRU_LUT4_0_LC_23_18_1.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_8_THRU_LUT4_0_LC_23_18_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_8_THRU_LUT4_0_LC_23_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_8_THRU_LUT4_0_LC_23_18_1 (
            .in0(_gnd_net_),
            .in1(N__26301),
            .in2(_gnd_net_),
            .in3(N__25542),
            .lcout(un1_M_this_sprites_address_q_cry_8_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_8),
            .carryout(un1_M_this_sprites_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_9_THRU_LUT4_0_LC_23_18_2.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_9_THRU_LUT4_0_LC_23_18_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_9_THRU_LUT4_0_LC_23_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_9_THRU_LUT4_0_LC_23_18_2 (
            .in0(_gnd_net_),
            .in1(N__25436),
            .in2(_gnd_net_),
            .in3(N__25407),
            .lcout(un1_M_this_sprites_address_q_cry_9_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_9),
            .carryout(un1_M_this_sprites_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_10_THRU_LUT4_0_LC_23_18_3.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_10_THRU_LUT4_0_LC_23_18_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_10_THRU_LUT4_0_LC_23_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_10_THRU_LUT4_0_LC_23_18_3 (
            .in0(_gnd_net_),
            .in1(N__30572),
            .in2(_gnd_net_),
            .in3(N__25398),
            .lcout(un1_M_this_sprites_address_q_cry_10_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_10),
            .carryout(un1_M_this_sprites_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_11_THRU_LUT4_0_LC_23_18_4.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_11_THRU_LUT4_0_LC_23_18_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_11_THRU_LUT4_0_LC_23_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_sprites_address_q_cry_11_THRU_LUT4_0_LC_23_18_4 (
            .in0(_gnd_net_),
            .in1(N__30653),
            .in2(_gnd_net_),
            .in3(N__25389),
            .lcout(un1_M_this_sprites_address_q_cry_11_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_11),
            .carryout(un1_M_this_sprites_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_13_LC_23_18_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_13_LC_23_18_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_13_LC_23_18_5.LUT_INIT=16'b0011101110110011;
    LogicCell40 M_this_sprites_address_q_13_LC_23_18_5 (
            .in0(N__27562),
            .in1(N__25386),
            .in2(N__30513),
            .in3(N__25380),
            .lcout(M_this_sprites_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32604),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_0_LC_23_18_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_0_LC_23_18_6.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_0_LC_23_18_6.LUT_INIT=16'b0101110111010101;
    LogicCell40 M_this_sprites_address_q_0_LC_23_18_6 (
            .in0(N__25377),
            .in1(N__27561),
            .in2(N__26458),
            .in3(N__25368),
            .lcout(M_this_sprites_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32604),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_9_LC_23_18_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_9_LC_23_18_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_9_LC_23_18_7.LUT_INIT=16'b0011101110110011;
    LogicCell40 M_this_sprites_address_q_9_LC_23_18_7 (
            .in0(N__27563),
            .in1(N__26424),
            .in2(N__26309),
            .in3(N__26415),
            .lcout(M_this_sprites_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32604),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI96JM1_LC_23_19_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI96JM1_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI96JM1_LC_23_19_1 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \this_start_data_delay.M_last_q_RNI96JM1_LC_23_19_1  (
            .in0(N__27933),
            .in1(N__26274),
            .in2(_gnd_net_),
            .in3(N__26200),
            .lcout(this_start_data_delay_M_this_external_address_q_3_i_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_23_19_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_23_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_23_19_2  (
            .in0(N__25851),
            .in1(N__25839),
            .in2(_gnd_net_),
            .in3(N__30088),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_12_LC_23_20_2.C_ON=1'b0;
    defparam M_this_data_count_q_12_LC_23_20_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_23_20_2.LUT_INIT=16'b1110010001000100;
    LogicCell40 M_this_data_count_q_12_LC_23_20_2 (
            .in0(N__29226),
            .in1(N__29892),
            .in2(N__28294),
            .in3(N__26975),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32619),
            .ce(N__29109),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_0_LC_23_20_5.C_ON=1'b0;
    defparam M_this_data_count_q_0_LC_23_20_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_23_20_5.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_0_LC_23_20_5 (
            .in0(_gnd_net_),
            .in1(N__29225),
            .in2(_gnd_net_),
            .in3(N__28512),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32619),
            .ce(N__29109),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_d62_10_LC_23_21_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d62_10_LC_23_21_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d62_10_LC_23_21_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.M_this_state_d62_10_LC_23_21_1  (
            .in0(N__29020),
            .in1(N__28492),
            .in2(N__28995),
            .in3(N__28510),
            .lcout(\this_start_data_delay.M_this_state_d62Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_15_LC_23_21_3.C_ON=1'b0;
    defparam M_this_data_count_q_15_LC_23_21_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_15_LC_23_21_3.LUT_INIT=16'b1100000010101010;
    LogicCell40 M_this_data_count_q_15_LC_23_21_3 (
            .in0(N__29256),
            .in1(N__26972),
            .in2(N__27941),
            .in3(N__29227),
            .lcout(M_this_data_count_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32627),
            .ce(N__29101),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_1_LC_23_21_6.C_ON=1'b0;
    defparam M_this_data_count_q_1_LC_23_21_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_23_21_6.LUT_INIT=16'b0000101000000101;
    LogicCell40 M_this_data_count_q_1_LC_23_21_6 (
            .in0(N__28493),
            .in1(_gnd_net_),
            .in2(N__29238),
            .in3(N__28479),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32627),
            .ce(N__29101),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_2_LC_23_21_7.C_ON=1'b0;
    defparam M_this_data_count_q_2_LC_23_21_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_23_21_7.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_2_LC_23_21_7 (
            .in0(N__29021),
            .in1(N__29007),
            .in2(_gnd_net_),
            .in3(N__29231),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32627),
            .ce(N__29101),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_11_LC_23_22_0.C_ON=1'b0;
    defparam M_this_data_count_q_11_LC_23_22_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_23_22_0.LUT_INIT=16'b1110010001000100;
    LogicCell40 M_this_data_count_q_11_LC_23_22_0 (
            .in0(N__29236),
            .in1(N__29922),
            .in2(N__26979),
            .in3(N__31296),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32632),
            .ce(N__29085),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_d62_8_LC_23_22_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d62_8_LC_23_22_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d62_8_LC_23_22_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.M_this_state_d62_8_LC_23_22_1  (
            .in0(N__29959),
            .in1(N__28817),
            .in2(N__29937),
            .in3(N__28844),
            .lcout(\this_start_data_delay.M_this_state_d62Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_d62_9_LC_23_22_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d62_9_LC_23_22_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d62_9_LC_23_22_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.M_this_state_d62_9_LC_23_22_3  (
            .in0(N__29315),
            .in1(N__29875),
            .in2(N__29274),
            .in3(N__29909),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_state_d62Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_d62_LC_23_22_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d62_LC_23_22_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d62_LC_23_22_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_start_data_delay.M_this_state_d62_LC_23_22_4  (
            .in0(N__26898),
            .in1(N__26892),
            .in2(N__26886),
            .in3(N__26883),
            .lcout(\this_start_data_delay.M_this_state_dZ0Z62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_10_LC_23_22_5.C_ON=1'b0;
    defparam M_this_data_count_q_10_LC_23_22_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_23_22_5.LUT_INIT=16'b1111000010011001;
    LogicCell40 M_this_data_count_q_10_LC_23_22_5 (
            .in0(N__29960),
            .in1(N__29946),
            .in2(N__26811),
            .in3(N__29237),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32632),
            .ce(N__29085),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_8_LC_23_24_0.C_ON=1'b0;
    defparam M_this_external_address_q_8_LC_23_24_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_8_LC_23_24_0.LUT_INIT=16'b1100000010101010;
    LogicCell40 M_this_external_address_q_8_LC_23_24_0 (
            .in0(N__30969),
            .in1(N__32932),
            .in2(N__28455),
            .in3(N__32735),
            .lcout(M_this_external_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32641),
            .ce(N__32220),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_15_LC_23_24_6.C_ON=1'b0;
    defparam M_this_external_address_q_15_LC_23_24_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_15_LC_23_24_6.LUT_INIT=16'b0010001011110000;
    LogicCell40 M_this_external_address_q_15_LC_23_24_6 (
            .in0(N__26802),
            .in1(N__26787),
            .in2(N__31377),
            .in3(N__32734),
            .lcout(M_this_external_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32641),
            .ce(N__32220),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_13_LC_23_24_7.C_ON=1'b0;
    defparam M_this_external_address_q_13_LC_23_24_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_13_LC_23_24_7.LUT_INIT=16'b0001010010111110;
    LogicCell40 M_this_external_address_q_13_LC_23_24_7 (
            .in0(N__32733),
            .in1(N__31486),
            .in2(N__31467),
            .in3(N__26703),
            .lcout(M_this_external_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32641),
            .ce(N__32220),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI5F621_2_LC_23_31_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI5F621_2_LC_23_31_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI5F621_2_LC_23_31_1 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \this_ppu.M_state_q_RNI5F621_2_LC_23_31_1  (
            .in0(N__26697),
            .in1(N__26676),
            .in2(N__31964),
            .in3(N__32131),
            .lcout(M_this_ppu_sprites_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_13_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_13_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_13_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_13_1  (
            .in0(N__30519),
            .in1(N__30606),
            .in2(N__30697),
            .in3(N__30751),
            .lcout(\this_sprites_ram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_13_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_13_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_13_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_13_6  (
            .in0(N__30752),
            .in1(N__30520),
            .in2(N__30614),
            .in3(N__30681),
            .lcout(\this_sprites_ram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_14_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_14_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_14_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_14_1  (
            .in0(N__30754),
            .in1(N__30685),
            .in2(N__30526),
            .in3(N__30594),
            .lcout(\this_sprites_ram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_14_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_14_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_14_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_14_4  (
            .in0(N__30593),
            .in1(N__30515),
            .in2(N__30698),
            .in3(N__30753),
            .lcout(\this_sprites_ram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI0IEC3_LC_24_15_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI0IEC3_LC_24_15_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI0IEC3_LC_24_15_3 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNI0IEC3_LC_24_15_3  (
            .in0(N__32904),
            .in1(N__27984),
            .in2(N__28108),
            .in3(N__27830),
            .lcout(N_811_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_5_LC_24_16_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_5_LC_24_16_2.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_5_LC_24_16_2.LUT_INIT=16'b0101110111010101;
    LogicCell40 M_this_sprites_address_q_5_LC_24_16_2 (
            .in0(N__27186),
            .in1(N__27560),
            .in2(N__27074),
            .in3(N__27180),
            .lcout(M_this_sprites_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32594),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_17_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_17_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_17_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_17_0  (
            .in0(N__30481),
            .in1(N__30591),
            .in2(N__30699),
            .in3(N__30739),
            .lcout(\this_sprites_ram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_24_17_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_24_17_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_24_17_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_24_17_2  (
            .in0(N__27018),
            .in1(N__27006),
            .in2(_gnd_net_),
            .in3(N__30105),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3_0_LC_24_17_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3_0_LC_24_17_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3_0_LC_24_17_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3_0_LC_24_17_5  (
            .in0(N__28473),
            .in1(N__28285),
            .in2(N__30936),
            .in3(N__28096),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_0_LC_24_17_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_0_LC_24_17_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_0_LC_24_17_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_0_LC_24_17_6  (
            .in0(_gnd_net_),
            .in1(N__27916),
            .in2(N__28047),
            .in3(N__31323),
            .lcout(\this_start_data_delay.N_902_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI2KEC3_LC_24_17_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI2KEC3_LC_24_17_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI2KEC3_LC_24_17_7 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNI2KEC3_LC_24_17_7  (
            .in0(N__31322),
            .in1(N__27978),
            .in2(N__27929),
            .in3(N__27834),
            .lcout(N_41_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_24_18_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_24_18_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_24_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_24_18_0  (
            .in0(N__30089),
            .in1(N__27732),
            .in2(_gnd_net_),
            .in3(N__27726),
            .lcout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_24_18_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_24_18_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_24_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_24_18_1  (
            .in0(N__30090),
            .in1(N__27711),
            .in2(_gnd_net_),
            .in3(N__27705),
            .lcout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_24_18_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_24_18_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_24_18_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_24_18_3  (
            .in0(N__30091),
            .in1(N__27687),
            .in2(_gnd_net_),
            .in3(N__27675),
            .lcout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI433C3_0_LC_24_18_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI433C3_0_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI433C3_0_LC_24_18_4 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \this_start_data_delay.M_last_q_RNI433C3_0_LC_24_18_4  (
            .in0(N__27379),
            .in1(N__27663),
            .in2(N__30934),
            .in3(N__27612),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_sprites_address_q_0_0_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_8_LC_24_18_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_8_LC_24_18_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_8_LC_24_18_5.LUT_INIT=16'b0110111100001111;
    LogicCell40 M_this_sprites_address_q_8_LC_24_18_5 (
            .in0(N__27378),
            .in1(N__27573),
            .in2(N__27567),
            .in3(N__27564),
            .lcout(M_this_sprites_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32613),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_24_19_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_24_19_2 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_24_19_2  (
            .in0(N__28667),
            .in1(N__27354),
            .in2(N__28728),
            .in3(N__28806),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_24_19_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_24_19_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_24_19_3  (
            .in0(N__28676),
            .in1(N__29991),
            .in2(N__28800),
            .in3(N__28797),
            .lcout(M_this_ppu_vram_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_24_19_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_24_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_24_19_6  (
            .in0(N__30076),
            .in1(N__28755),
            .in2(_gnd_net_),
            .in3(N__28743),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_24_19_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_24_19_7 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_24_19_7  (
            .in0(N__28720),
            .in1(N__28686),
            .in2(N__28680),
            .in3(N__28666),
            .lcout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_24_20_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_24_20_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_24_20_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_24_20_0  (
            .in0(N__30095),
            .in1(N__28614),
            .in2(_gnd_net_),
            .in3(N__28602),
            .lcout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_20_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_20_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_20_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_20_3  (
            .in0(N__30755),
            .in1(N__30514),
            .in2(N__30704),
            .in3(N__30605),
            .lcout(\this_sprites_ram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_24_20_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_24_20_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_24_20_7  (
            .in0(N__28554),
            .in1(N__28539),
            .in2(_gnd_net_),
            .in3(N__30096),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_c_0_LC_24_21_0.C_ON=1'b1;
    defparam M_this_data_count_q_cry_c_0_LC_24_21_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_c_0_LC_24_21_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 M_this_data_count_q_cry_c_0_LC_24_21_0 (
            .in0(_gnd_net_),
            .in1(N__28511),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_24_21_0_),
            .carryout(M_this_data_count_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_24_21_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_24_21_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_24_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_0_THRU_LUT4_0_LC_24_21_1 (
            .in0(_gnd_net_),
            .in1(N__28494),
            .in2(N__29682),
            .in3(N__29025),
            .lcout(M_this_data_count_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_0),
            .carryout(M_this_data_count_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_24_21_2.C_ON=1'b1;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_24_21_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_24_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_1_THRU_LUT4_0_LC_24_21_2 (
            .in0(_gnd_net_),
            .in1(N__29022),
            .in2(N__29680),
            .in3(N__28998),
            .lcout(M_this_data_count_q_cry_1_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_1),
            .carryout(M_this_data_count_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_24_21_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_24_21_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_24_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_2_THRU_LUT4_0_LC_24_21_3 (
            .in0(_gnd_net_),
            .in1(N__28994),
            .in2(N__29683),
            .in3(N__28950),
            .lcout(M_this_data_count_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_2),
            .carryout(M_this_data_count_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_24_21_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_24_21_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_24_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_3_THRU_LUT4_0_LC_24_21_4 (
            .in0(_gnd_net_),
            .in1(N__29135),
            .in2(N__29681),
            .in3(N__28947),
            .lcout(M_this_data_count_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_3),
            .carryout(M_this_data_count_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_24_21_5.C_ON=1'b1;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_24_21_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_24_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_4_THRU_LUT4_0_LC_24_21_5 (
            .in0(_gnd_net_),
            .in1(N__28944),
            .in2(N__29684),
            .in3(N__28917),
            .lcout(M_this_data_count_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_4),
            .carryout(M_this_data_count_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_6_LC_24_21_6.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_6_LC_24_21_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_6_LC_24_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_6_LC_24_21_6 (
            .in0(_gnd_net_),
            .in1(N__28914),
            .in2(N__29679),
            .in3(N__28890),
            .lcout(M_this_data_count_q_s_6),
            .ltout(),
            .carryin(M_this_data_count_q_cry_5),
            .carryout(M_this_data_count_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_24_21_7.C_ON=1'b1;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_24_21_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_24_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_6_THRU_LUT4_0_LC_24_21_7 (
            .in0(_gnd_net_),
            .in1(N__28887),
            .in2(N__29685),
            .in3(N__28857),
            .lcout(M_this_data_count_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_6),
            .carryout(M_this_data_count_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_8_LC_24_22_0.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_8_LC_24_22_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_8_LC_24_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_8_LC_24_22_0 (
            .in0(_gnd_net_),
            .in1(N__29691),
            .in2(N__28854),
            .in3(N__28824),
            .lcout(M_this_data_count_q_s_8),
            .ltout(),
            .carryin(bfn_24_22_0_),
            .carryout(M_this_data_count_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_9_LC_24_22_1.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_9_LC_24_22_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_9_LC_24_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_9_LC_24_22_1 (
            .in0(_gnd_net_),
            .in1(N__28821),
            .in2(N__29752),
            .in3(N__29970),
            .lcout(M_this_data_count_q_s_9),
            .ltout(),
            .carryin(M_this_data_count_q_cry_8),
            .carryout(M_this_data_count_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_9_THRU_LUT4_0_LC_24_22_2.C_ON=1'b1;
    defparam M_this_data_count_q_cry_9_THRU_LUT4_0_LC_24_22_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_9_THRU_LUT4_0_LC_24_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_9_THRU_LUT4_0_LC_24_22_2 (
            .in0(_gnd_net_),
            .in1(N__29698),
            .in2(N__29967),
            .in3(N__29940),
            .lcout(M_this_data_count_q_cry_9_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_9),
            .carryout(M_this_data_count_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_11_LC_24_22_3.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_11_LC_24_22_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_11_LC_24_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_11_LC_24_22_3 (
            .in0(_gnd_net_),
            .in1(N__29936),
            .in2(N__29751),
            .in3(N__29916),
            .lcout(M_this_data_count_q_s_11),
            .ltout(),
            .carryin(M_this_data_count_q_cry_10),
            .carryout(M_this_data_count_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_12_LC_24_22_4.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_12_LC_24_22_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_12_LC_24_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_12_LC_24_22_4 (
            .in0(_gnd_net_),
            .in1(N__29689),
            .in2(N__29913),
            .in3(N__29883),
            .lcout(M_this_data_count_q_s_12),
            .ltout(),
            .carryin(M_this_data_count_q_cry_11),
            .carryout(M_this_data_count_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_12_THRU_LUT4_0_LC_24_22_5.C_ON=1'b1;
    defparam M_this_data_count_q_cry_12_THRU_LUT4_0_LC_24_22_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_12_THRU_LUT4_0_LC_24_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_12_THRU_LUT4_0_LC_24_22_5 (
            .in0(_gnd_net_),
            .in1(N__29880),
            .in2(N__29753),
            .in3(N__29847),
            .lcout(M_this_data_count_q_cry_12_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_12),
            .carryout(M_this_data_count_q_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_14_LC_24_22_6.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_14_LC_24_22_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_14_LC_24_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_14_LC_24_22_6 (
            .in0(_gnd_net_),
            .in1(N__29690),
            .in2(N__29319),
            .in3(N__29277),
            .lcout(M_this_data_count_q_s_14),
            .ltout(),
            .carryin(M_this_data_count_q_cry_13),
            .carryout(M_this_data_count_q_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_15_LC_24_22_7.C_ON=1'b0;
    defparam M_this_data_count_q_RNO_0_15_LC_24_22_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_15_LC_24_22_7.LUT_INIT=16'b1100110000110011;
    LogicCell40 M_this_data_count_q_RNO_0_15_LC_24_22_7 (
            .in0(_gnd_net_),
            .in1(N__29273),
            .in2(_gnd_net_),
            .in3(N__29259),
            .lcout(M_this_data_count_q_s_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_4_LC_24_23_0.C_ON=1'b0;
    defparam M_this_data_count_q_4_LC_24_23_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_24_23_0.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_4_LC_24_23_0 (
            .in0(N__29247),
            .in1(N__29232),
            .in2(_gnd_net_),
            .in3(N__29131),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32642),
            .ce(N__29102),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_12_LC_24_24_0.C_ON=1'b0;
    defparam M_this_external_address_q_12_LC_24_24_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_12_LC_24_24_0.LUT_INIT=16'b0011001101011010;
    LogicCell40 M_this_external_address_q_12_LC_24_24_0 (
            .in0(N__31512),
            .in1(N__30954),
            .in2(N__31538),
            .in3(N__32760),
            .lcout(M_this_external_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32644),
            .ce(N__32235),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_14_LC_24_24_1.C_ON=1'b0;
    defparam M_this_external_address_q_14_LC_24_24_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_14_LC_24_24_1.LUT_INIT=16'b1011111000010100;
    LogicCell40 M_this_external_address_q_14_LC_24_24_1 (
            .in0(N__32758),
            .in1(N__31416),
            .in2(N__31442),
            .in3(N__30945),
            .lcout(M_this_external_address_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32644),
            .ce(N__32235),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_9_LC_24_24_6.C_ON=1'b0;
    defparam M_this_external_address_q_9_LC_24_24_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_9_LC_24_24_6.LUT_INIT=16'b1100000010101010;
    LogicCell40 M_this_external_address_q_9_LC_24_24_6 (
            .in0(N__31560),
            .in1(N__32941),
            .in2(N__30915),
            .in3(N__32759),
            .lcout(M_this_external_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32644),
            .ce(N__32235),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_25_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_25_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_25_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_25_1  (
            .in0(N__30527),
            .in1(N__30610),
            .in2(N__30705),
            .in3(N__30761),
            .lcout(\this_sprites_ram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_25_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_25_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_25_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_25_2  (
            .in0(N__30762),
            .in1(N__30700),
            .in2(N__30615),
            .in3(N__30528),
            .lcout(\this_sprites_ram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIP0T41_2_LC_24_31_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIP0T41_2_LC_24_31_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIP0T41_2_LC_24_31_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \this_ppu.M_state_q_RNIP0T41_2_LC_24_31_4  (
            .in0(N__32129),
            .in1(N__31960),
            .in2(N__30429),
            .in3(N__30405),
            .lcout(M_this_ppu_sprites_addr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNI2HC01_2_LC_24_31_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNI2HC01_2_LC_24_31_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNI2HC01_2_LC_24_31_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \this_ppu.M_vaddress_q_RNI2HC01_2_LC_24_31_7  (
            .in0(N__30291),
            .in1(N__32128),
            .in2(N__31969),
            .in3(N__30249),
            .lcout(M_this_ppu_sprites_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_26_17_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_26_17_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_26_17_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_26_17_0  (
            .in0(N__30135),
            .in1(N__30117),
            .in2(_gnd_net_),
            .in3(N__30107),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_0_LC_26_23_0.C_ON=1'b1;
    defparam M_this_external_address_q_0_LC_26_23_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_0_LC_26_23_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_0_LC_26_23_0 (
            .in0(N__32752),
            .in1(N__31178),
            .in2(_gnd_net_),
            .in3(N__31167),
            .lcout(M_this_external_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_26_23_0_),
            .carryout(M_this_external_address_q_cry_0),
            .clk(N__32648),
            .ce(N__32233),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_1_LC_26_23_1.C_ON=1'b1;
    defparam M_this_external_address_q_1_LC_26_23_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_1_LC_26_23_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_1_LC_26_23_1 (
            .in0(N__32748),
            .in1(N__31157),
            .in2(_gnd_net_),
            .in3(N__31146),
            .lcout(M_this_external_address_qZ0Z_1),
            .ltout(),
            .carryin(M_this_external_address_q_cry_0),
            .carryout(M_this_external_address_q_cry_1),
            .clk(N__32648),
            .ce(N__32233),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_2_LC_26_23_2.C_ON=1'b1;
    defparam M_this_external_address_q_2_LC_26_23_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_2_LC_26_23_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_2_LC_26_23_2 (
            .in0(N__32753),
            .in1(N__31130),
            .in2(_gnd_net_),
            .in3(N__31119),
            .lcout(M_this_external_address_qZ0Z_2),
            .ltout(),
            .carryin(M_this_external_address_q_cry_1),
            .carryout(M_this_external_address_q_cry_2),
            .clk(N__32648),
            .ce(N__32233),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_3_LC_26_23_3.C_ON=1'b1;
    defparam M_this_external_address_q_3_LC_26_23_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_3_LC_26_23_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_3_LC_26_23_3 (
            .in0(N__32749),
            .in1(N__31103),
            .in2(_gnd_net_),
            .in3(N__31092),
            .lcout(M_this_external_address_qZ0Z_3),
            .ltout(),
            .carryin(M_this_external_address_q_cry_2),
            .carryout(M_this_external_address_q_cry_3),
            .clk(N__32648),
            .ce(N__32233),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_4_LC_26_23_4.C_ON=1'b1;
    defparam M_this_external_address_q_4_LC_26_23_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_4_LC_26_23_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_4_LC_26_23_4 (
            .in0(N__32754),
            .in1(N__31085),
            .in2(_gnd_net_),
            .in3(N__31074),
            .lcout(M_this_external_address_qZ0Z_4),
            .ltout(),
            .carryin(M_this_external_address_q_cry_3),
            .carryout(M_this_external_address_q_cry_4),
            .clk(N__32648),
            .ce(N__32233),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_5_LC_26_23_5.C_ON=1'b1;
    defparam M_this_external_address_q_5_LC_26_23_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_5_LC_26_23_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_5_LC_26_23_5 (
            .in0(N__32750),
            .in1(N__31061),
            .in2(_gnd_net_),
            .in3(N__31050),
            .lcout(M_this_external_address_qZ0Z_5),
            .ltout(),
            .carryin(M_this_external_address_q_cry_4),
            .carryout(M_this_external_address_q_cry_5),
            .clk(N__32648),
            .ce(N__32233),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_6_LC_26_23_6.C_ON=1'b1;
    defparam M_this_external_address_q_6_LC_26_23_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_6_LC_26_23_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_6_LC_26_23_6 (
            .in0(N__32755),
            .in1(N__31040),
            .in2(_gnd_net_),
            .in3(N__31029),
            .lcout(M_this_external_address_qZ0Z_6),
            .ltout(),
            .carryin(M_this_external_address_q_cry_5),
            .carryout(M_this_external_address_q_cry_6),
            .clk(N__32648),
            .ce(N__32233),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_7_LC_26_23_7.C_ON=1'b1;
    defparam M_this_external_address_q_7_LC_26_23_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_7_LC_26_23_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_7_LC_26_23_7 (
            .in0(N__32751),
            .in1(N__31010),
            .in2(_gnd_net_),
            .in3(N__30999),
            .lcout(M_this_external_address_qZ0Z_7),
            .ltout(),
            .carryin(M_this_external_address_q_cry_6),
            .carryout(M_this_external_address_q_cry_7),
            .clk(N__32648),
            .ce(N__32233),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNO_0_8_LC_26_24_0.C_ON=1'b1;
    defparam M_this_external_address_q_RNO_0_8_LC_26_24_0.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNO_0_8_LC_26_24_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_external_address_q_RNO_0_8_LC_26_24_0 (
            .in0(_gnd_net_),
            .in1(N__30986),
            .in2(_gnd_net_),
            .in3(N__30957),
            .lcout(M_this_external_address_q_s_8),
            .ltout(),
            .carryin(bfn_26_24_0_),
            .carryout(M_this_external_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNO_0_9_LC_26_24_1.C_ON=1'b1;
    defparam M_this_external_address_q_RNO_0_9_LC_26_24_1.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNO_0_9_LC_26_24_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_external_address_q_RNO_0_9_LC_26_24_1 (
            .in0(_gnd_net_),
            .in1(N__31577),
            .in2(_gnd_net_),
            .in3(N__31551),
            .lcout(M_this_external_address_q_s_9),
            .ltout(),
            .carryin(M_this_external_address_q_cry_8),
            .carryout(M_this_external_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNO_0_10_LC_26_24_2.C_ON=1'b1;
    defparam M_this_external_address_q_RNO_0_10_LC_26_24_2.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNO_0_10_LC_26_24_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_external_address_q_RNO_0_10_LC_26_24_2 (
            .in0(_gnd_net_),
            .in1(N__32675),
            .in2(_gnd_net_),
            .in3(N__31548),
            .lcout(M_this_external_address_q_s_10),
            .ltout(),
            .carryin(M_this_external_address_q_cry_9),
            .carryout(M_this_external_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNO_0_11_LC_26_24_3.C_ON=1'b1;
    defparam M_this_external_address_q_RNO_0_11_LC_26_24_3.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNO_0_11_LC_26_24_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_external_address_q_RNO_0_11_LC_26_24_3 (
            .in0(_gnd_net_),
            .in1(N__31202),
            .in2(_gnd_net_),
            .in3(N__31545),
            .lcout(M_this_external_address_q_s_11),
            .ltout(),
            .carryin(M_this_external_address_q_cry_10),
            .carryout(M_this_external_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_cry_11_THRU_LUT4_0_LC_26_24_4.C_ON=1'b1;
    defparam M_this_external_address_q_cry_11_THRU_LUT4_0_LC_26_24_4.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_cry_11_THRU_LUT4_0_LC_26_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_external_address_q_cry_11_THRU_LUT4_0_LC_26_24_4 (
            .in0(_gnd_net_),
            .in1(N__31537),
            .in2(_gnd_net_),
            .in3(N__31503),
            .lcout(M_this_external_address_q_cry_11_THRU_CO),
            .ltout(),
            .carryin(M_this_external_address_q_cry_11),
            .carryout(M_this_external_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_cry_12_THRU_LUT4_0_LC_26_24_5.C_ON=1'b1;
    defparam M_this_external_address_q_cry_12_THRU_LUT4_0_LC_26_24_5.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_cry_12_THRU_LUT4_0_LC_26_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_external_address_q_cry_12_THRU_LUT4_0_LC_26_24_5 (
            .in0(_gnd_net_),
            .in1(N__31490),
            .in2(_gnd_net_),
            .in3(N__31455),
            .lcout(M_this_external_address_q_cry_12_THRU_CO),
            .ltout(),
            .carryin(M_this_external_address_q_cry_12),
            .carryout(M_this_external_address_q_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_cry_13_THRU_LUT4_0_LC_26_24_6.C_ON=1'b1;
    defparam M_this_external_address_q_cry_13_THRU_LUT4_0_LC_26_24_6.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_cry_13_THRU_LUT4_0_LC_26_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_external_address_q_cry_13_THRU_LUT4_0_LC_26_24_6 (
            .in0(_gnd_net_),
            .in1(N__31441),
            .in2(_gnd_net_),
            .in3(N__31407),
            .lcout(M_this_external_address_q_cry_13_THRU_CO),
            .ltout(),
            .carryin(M_this_external_address_q_cry_13),
            .carryout(M_this_external_address_q_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNO_0_15_LC_26_24_7.C_ON=1'b0;
    defparam M_this_external_address_q_RNO_0_15_LC_26_24_7.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNO_0_15_LC_26_24_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 M_this_external_address_q_RNO_0_15_LC_26_24_7 (
            .in0(_gnd_net_),
            .in1(N__31397),
            .in2(_gnd_net_),
            .in3(N__31380),
            .lcout(M_this_external_address_q_s_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_11_LC_26_25_1.C_ON=1'b0;
    defparam M_this_external_address_q_11_LC_26_25_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_11_LC_26_25_1.LUT_INIT=16'b1110010001000100;
    LogicCell40 M_this_external_address_q_11_LC_26_25_1 (
            .in0(N__32756),
            .in1(N__31365),
            .in2(N__31295),
            .in3(N__32949),
            .lcout(M_this_external_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32654),
            .ce(N__32234),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_10_LC_26_25_2.C_ON=1'b0;
    defparam M_this_external_address_q_10_LC_26_25_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_10_LC_26_25_2.LUT_INIT=16'b1100000010101010;
    LogicCell40 M_this_external_address_q_10_LC_26_25_2 (
            .in0(N__32955),
            .in1(N__32948),
            .in2(N__32819),
            .in3(N__32757),
            .lcout(M_this_external_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32654),
            .ce(N__32234),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIVCB01_1_LC_26_31_2 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIVCB01_1_LC_26_31_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIVCB01_1_LC_26_31_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \this_ppu.M_vaddress_q_RNIVCB01_1_LC_26_31_2  (
            .in0(N__32187),
            .in1(N__32130),
            .in2(N__31970),
            .in3(N__31806),
            .lcout(M_this_ppu_sprites_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un1_M_this_state_q_17_i_o2_1_4_LC_32_19_7 .C_ON=1'b0;
    defparam \this_start_data_delay.un1_M_this_state_q_17_i_o2_1_4_LC_32_19_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un1_M_this_state_q_17_i_o2_1_4_LC_32_19_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.un1_M_this_state_q_17_i_o2_1_4_LC_32_19_7  (
            .in0(N__31689),
            .in1(N__31668),
            .in2(N__31656),
            .in3(N__31608),
            .lcout(\this_start_data_delay.un1_M_this_state_q_17_i_o2_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
