// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     Jun 1 2022 09:54:43

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    led,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    inout [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output [7:0] led;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__44416;
    wire N__44415;
    wire N__44414;
    wire N__44405;
    wire N__44404;
    wire N__44403;
    wire N__44396;
    wire N__44395;
    wire N__44394;
    wire N__44387;
    wire N__44386;
    wire N__44385;
    wire N__44378;
    wire N__44377;
    wire N__44376;
    wire N__44369;
    wire N__44368;
    wire N__44367;
    wire N__44360;
    wire N__44359;
    wire N__44358;
    wire N__44351;
    wire N__44350;
    wire N__44349;
    wire N__44342;
    wire N__44341;
    wire N__44340;
    wire N__44333;
    wire N__44332;
    wire N__44331;
    wire N__44324;
    wire N__44323;
    wire N__44322;
    wire N__44315;
    wire N__44314;
    wire N__44313;
    wire N__44306;
    wire N__44305;
    wire N__44304;
    wire N__44297;
    wire N__44296;
    wire N__44295;
    wire N__44288;
    wire N__44287;
    wire N__44286;
    wire N__44279;
    wire N__44278;
    wire N__44277;
    wire N__44270;
    wire N__44269;
    wire N__44268;
    wire N__44261;
    wire N__44260;
    wire N__44259;
    wire N__44252;
    wire N__44251;
    wire N__44250;
    wire N__44243;
    wire N__44242;
    wire N__44241;
    wire N__44234;
    wire N__44233;
    wire N__44232;
    wire N__44225;
    wire N__44224;
    wire N__44223;
    wire N__44216;
    wire N__44215;
    wire N__44214;
    wire N__44207;
    wire N__44206;
    wire N__44205;
    wire N__44198;
    wire N__44197;
    wire N__44196;
    wire N__44189;
    wire N__44188;
    wire N__44187;
    wire N__44180;
    wire N__44179;
    wire N__44178;
    wire N__44171;
    wire N__44170;
    wire N__44169;
    wire N__44162;
    wire N__44161;
    wire N__44160;
    wire N__44153;
    wire N__44152;
    wire N__44151;
    wire N__44144;
    wire N__44143;
    wire N__44142;
    wire N__44135;
    wire N__44134;
    wire N__44133;
    wire N__44126;
    wire N__44125;
    wire N__44124;
    wire N__44117;
    wire N__44116;
    wire N__44115;
    wire N__44108;
    wire N__44107;
    wire N__44106;
    wire N__44099;
    wire N__44098;
    wire N__44097;
    wire N__44090;
    wire N__44089;
    wire N__44088;
    wire N__44081;
    wire N__44080;
    wire N__44079;
    wire N__44072;
    wire N__44071;
    wire N__44070;
    wire N__44063;
    wire N__44062;
    wire N__44061;
    wire N__44054;
    wire N__44053;
    wire N__44052;
    wire N__44045;
    wire N__44044;
    wire N__44043;
    wire N__44036;
    wire N__44035;
    wire N__44034;
    wire N__44027;
    wire N__44026;
    wire N__44025;
    wire N__44018;
    wire N__44017;
    wire N__44016;
    wire N__44009;
    wire N__44008;
    wire N__44007;
    wire N__44000;
    wire N__43999;
    wire N__43998;
    wire N__43991;
    wire N__43990;
    wire N__43989;
    wire N__43982;
    wire N__43981;
    wire N__43980;
    wire N__43973;
    wire N__43972;
    wire N__43971;
    wire N__43964;
    wire N__43963;
    wire N__43962;
    wire N__43955;
    wire N__43954;
    wire N__43953;
    wire N__43936;
    wire N__43935;
    wire N__43932;
    wire N__43929;
    wire N__43926;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43912;
    wire N__43909;
    wire N__43906;
    wire N__43903;
    wire N__43900;
    wire N__43897;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43874;
    wire N__43869;
    wire N__43866;
    wire N__43861;
    wire N__43858;
    wire N__43855;
    wire N__43854;
    wire N__43851;
    wire N__43848;
    wire N__43847;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43835;
    wire N__43832;
    wire N__43829;
    wire N__43826;
    wire N__43823;
    wire N__43820;
    wire N__43813;
    wire N__43810;
    wire N__43807;
    wire N__43806;
    wire N__43803;
    wire N__43800;
    wire N__43799;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43781;
    wire N__43778;
    wire N__43775;
    wire N__43772;
    wire N__43767;
    wire N__43764;
    wire N__43761;
    wire N__43756;
    wire N__43753;
    wire N__43750;
    wire N__43747;
    wire N__43746;
    wire N__43743;
    wire N__43740;
    wire N__43737;
    wire N__43734;
    wire N__43731;
    wire N__43728;
    wire N__43725;
    wire N__43722;
    wire N__43719;
    wire N__43714;
    wire N__43711;
    wire N__43708;
    wire N__43705;
    wire N__43704;
    wire N__43703;
    wire N__43700;
    wire N__43697;
    wire N__43696;
    wire N__43695;
    wire N__43692;
    wire N__43687;
    wire N__43682;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43665;
    wire N__43664;
    wire N__43659;
    wire N__43656;
    wire N__43653;
    wire N__43650;
    wire N__43647;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43612;
    wire N__43609;
    wire N__43608;
    wire N__43605;
    wire N__43602;
    wire N__43599;
    wire N__43596;
    wire N__43593;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43576;
    wire N__43575;
    wire N__43574;
    wire N__43573;
    wire N__43572;
    wire N__43569;
    wire N__43568;
    wire N__43567;
    wire N__43566;
    wire N__43565;
    wire N__43564;
    wire N__43563;
    wire N__43562;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43548;
    wire N__43547;
    wire N__43546;
    wire N__43545;
    wire N__43544;
    wire N__43543;
    wire N__43530;
    wire N__43529;
    wire N__43528;
    wire N__43517;
    wire N__43504;
    wire N__43503;
    wire N__43502;
    wire N__43501;
    wire N__43500;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43490;
    wire N__43489;
    wire N__43488;
    wire N__43487;
    wire N__43486;
    wire N__43485;
    wire N__43484;
    wire N__43481;
    wire N__43478;
    wire N__43475;
    wire N__43472;
    wire N__43471;
    wire N__43470;
    wire N__43467;
    wire N__43464;
    wire N__43461;
    wire N__43460;
    wire N__43457;
    wire N__43454;
    wire N__43447;
    wire N__43440;
    wire N__43433;
    wire N__43432;
    wire N__43431;
    wire N__43428;
    wire N__43425;
    wire N__43420;
    wire N__43417;
    wire N__43416;
    wire N__43415;
    wire N__43412;
    wire N__43405;
    wire N__43402;
    wire N__43401;
    wire N__43398;
    wire N__43389;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43373;
    wire N__43372;
    wire N__43371;
    wire N__43366;
    wire N__43365;
    wire N__43362;
    wire N__43357;
    wire N__43356;
    wire N__43355;
    wire N__43354;
    wire N__43351;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43335;
    wire N__43332;
    wire N__43329;
    wire N__43326;
    wire N__43323;
    wire N__43318;
    wire N__43311;
    wire N__43306;
    wire N__43285;
    wire N__43282;
    wire N__43279;
    wire N__43276;
    wire N__43275;
    wire N__43272;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43259;
    wire N__43252;
    wire N__43251;
    wire N__43250;
    wire N__43249;
    wire N__43248;
    wire N__43245;
    wire N__43244;
    wire N__43243;
    wire N__43242;
    wire N__43241;
    wire N__43240;
    wire N__43239;
    wire N__43238;
    wire N__43237;
    wire N__43236;
    wire N__43235;
    wire N__43234;
    wire N__43233;
    wire N__43232;
    wire N__43229;
    wire N__43228;
    wire N__43227;
    wire N__43226;
    wire N__43225;
    wire N__43224;
    wire N__43223;
    wire N__43222;
    wire N__43221;
    wire N__43220;
    wire N__43219;
    wire N__43218;
    wire N__43217;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43197;
    wire N__43194;
    wire N__43191;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43166;
    wire N__43163;
    wire N__43158;
    wire N__43153;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43138;
    wire N__43135;
    wire N__43132;
    wire N__43131;
    wire N__43130;
    wire N__43129;
    wire N__43128;
    wire N__43127;
    wire N__43126;
    wire N__43125;
    wire N__43124;
    wire N__43123;
    wire N__43122;
    wire N__43121;
    wire N__43120;
    wire N__43119;
    wire N__43118;
    wire N__43117;
    wire N__43116;
    wire N__43115;
    wire N__43114;
    wire N__43113;
    wire N__43112;
    wire N__43111;
    wire N__43110;
    wire N__43109;
    wire N__43108;
    wire N__43107;
    wire N__43106;
    wire N__43105;
    wire N__43104;
    wire N__43103;
    wire N__43102;
    wire N__43101;
    wire N__43100;
    wire N__43099;
    wire N__43098;
    wire N__43097;
    wire N__43094;
    wire N__43091;
    wire N__43088;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43067;
    wire N__43064;
    wire N__43061;
    wire N__43058;
    wire N__43055;
    wire N__43052;
    wire N__43049;
    wire N__43046;
    wire N__43043;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43028;
    wire N__43025;
    wire N__43022;
    wire N__42901;
    wire N__42898;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42880;
    wire N__42877;
    wire N__42874;
    wire N__42871;
    wire N__42870;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42847;
    wire N__42844;
    wire N__42835;
    wire N__42834;
    wire N__42831;
    wire N__42830;
    wire N__42829;
    wire N__42828;
    wire N__42825;
    wire N__42822;
    wire N__42817;
    wire N__42814;
    wire N__42807;
    wire N__42804;
    wire N__42801;
    wire N__42796;
    wire N__42793;
    wire N__42792;
    wire N__42791;
    wire N__42788;
    wire N__42785;
    wire N__42782;
    wire N__42775;
    wire N__42774;
    wire N__42773;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42765;
    wire N__42764;
    wire N__42761;
    wire N__42758;
    wire N__42757;
    wire N__42754;
    wire N__42751;
    wire N__42750;
    wire N__42747;
    wire N__42744;
    wire N__42741;
    wire N__42738;
    wire N__42735;
    wire N__42732;
    wire N__42729;
    wire N__42726;
    wire N__42723;
    wire N__42720;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42710;
    wire N__42703;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42689;
    wire N__42686;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42670;
    wire N__42667;
    wire N__42658;
    wire N__42655;
    wire N__42652;
    wire N__42649;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42637;
    wire N__42636;
    wire N__42633;
    wire N__42630;
    wire N__42625;
    wire N__42622;
    wire N__42619;
    wire N__42616;
    wire N__42615;
    wire N__42614;
    wire N__42611;
    wire N__42608;
    wire N__42605;
    wire N__42598;
    wire N__42595;
    wire N__42594;
    wire N__42593;
    wire N__42592;
    wire N__42589;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42568;
    wire N__42565;
    wire N__42562;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42544;
    wire N__42543;
    wire N__42542;
    wire N__42541;
    wire N__42540;
    wire N__42539;
    wire N__42536;
    wire N__42533;
    wire N__42530;
    wire N__42529;
    wire N__42526;
    wire N__42523;
    wire N__42520;
    wire N__42517;
    wire N__42514;
    wire N__42509;
    wire N__42508;
    wire N__42507;
    wire N__42500;
    wire N__42499;
    wire N__42496;
    wire N__42493;
    wire N__42490;
    wire N__42487;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42463;
    wire N__42460;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42449;
    wire N__42446;
    wire N__42445;
    wire N__42444;
    wire N__42443;
    wire N__42440;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42430;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42416;
    wire N__42415;
    wire N__42412;
    wire N__42407;
    wire N__42404;
    wire N__42401;
    wire N__42398;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42368;
    wire N__42363;
    wire N__42358;
    wire N__42355;
    wire N__42352;
    wire N__42347;
    wire N__42342;
    wire N__42339;
    wire N__42334;
    wire N__42329;
    wire N__42324;
    wire N__42319;
    wire N__42316;
    wire N__42313;
    wire N__42310;
    wire N__42307;
    wire N__42304;
    wire N__42301;
    wire N__42298;
    wire N__42295;
    wire N__42294;
    wire N__42293;
    wire N__42290;
    wire N__42289;
    wire N__42288;
    wire N__42285;
    wire N__42284;
    wire N__42283;
    wire N__42280;
    wire N__42277;
    wire N__42274;
    wire N__42271;
    wire N__42268;
    wire N__42263;
    wire N__42262;
    wire N__42261;
    wire N__42260;
    wire N__42259;
    wire N__42258;
    wire N__42255;
    wire N__42250;
    wire N__42247;
    wire N__42244;
    wire N__42241;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42227;
    wire N__42220;
    wire N__42217;
    wire N__42214;
    wire N__42211;
    wire N__42208;
    wire N__42205;
    wire N__42190;
    wire N__42187;
    wire N__42184;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42174;
    wire N__42171;
    wire N__42168;
    wire N__42167;
    wire N__42164;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42152;
    wire N__42145;
    wire N__42144;
    wire N__42143;
    wire N__42142;
    wire N__42141;
    wire N__42140;
    wire N__42139;
    wire N__42138;
    wire N__42137;
    wire N__42136;
    wire N__42135;
    wire N__42134;
    wire N__42133;
    wire N__42132;
    wire N__42131;
    wire N__42130;
    wire N__42129;
    wire N__42128;
    wire N__42127;
    wire N__42126;
    wire N__42125;
    wire N__42124;
    wire N__42123;
    wire N__42122;
    wire N__42121;
    wire N__42120;
    wire N__42119;
    wire N__42118;
    wire N__42117;
    wire N__42116;
    wire N__42115;
    wire N__42114;
    wire N__42113;
    wire N__42112;
    wire N__42111;
    wire N__42110;
    wire N__42109;
    wire N__42108;
    wire N__42107;
    wire N__42106;
    wire N__42105;
    wire N__42104;
    wire N__42103;
    wire N__42102;
    wire N__42101;
    wire N__42100;
    wire N__42099;
    wire N__42098;
    wire N__42097;
    wire N__42096;
    wire N__42095;
    wire N__42094;
    wire N__42093;
    wire N__42092;
    wire N__42091;
    wire N__42090;
    wire N__42089;
    wire N__42088;
    wire N__42087;
    wire N__42086;
    wire N__42085;
    wire N__42084;
    wire N__42083;
    wire N__42082;
    wire N__42081;
    wire N__42080;
    wire N__42079;
    wire N__42078;
    wire N__42077;
    wire N__42076;
    wire N__42075;
    wire N__42074;
    wire N__42073;
    wire N__42072;
    wire N__42071;
    wire N__42070;
    wire N__42069;
    wire N__42068;
    wire N__42067;
    wire N__42066;
    wire N__42065;
    wire N__42064;
    wire N__42063;
    wire N__42062;
    wire N__42061;
    wire N__42060;
    wire N__42059;
    wire N__42058;
    wire N__42057;
    wire N__42056;
    wire N__42055;
    wire N__42054;
    wire N__42053;
    wire N__42052;
    wire N__42051;
    wire N__42050;
    wire N__42049;
    wire N__42048;
    wire N__42047;
    wire N__42046;
    wire N__42045;
    wire N__42044;
    wire N__42043;
    wire N__42042;
    wire N__42041;
    wire N__42040;
    wire N__42039;
    wire N__42038;
    wire N__42037;
    wire N__42036;
    wire N__42035;
    wire N__42034;
    wire N__42033;
    wire N__42032;
    wire N__42031;
    wire N__42030;
    wire N__42029;
    wire N__42028;
    wire N__42027;
    wire N__42026;
    wire N__42025;
    wire N__42024;
    wire N__42023;
    wire N__42022;
    wire N__42021;
    wire N__42020;
    wire N__42019;
    wire N__42018;
    wire N__42017;
    wire N__42016;
    wire N__42015;
    wire N__42014;
    wire N__42013;
    wire N__42012;
    wire N__42011;
    wire N__42010;
    wire N__42009;
    wire N__42008;
    wire N__42007;
    wire N__42006;
    wire N__42005;
    wire N__42004;
    wire N__42003;
    wire N__42002;
    wire N__42001;
    wire N__42000;
    wire N__41999;
    wire N__41998;
    wire N__41997;
    wire N__41996;
    wire N__41995;
    wire N__41994;
    wire N__41993;
    wire N__41992;
    wire N__41991;
    wire N__41990;
    wire N__41989;
    wire N__41988;
    wire N__41987;
    wire N__41986;
    wire N__41985;
    wire N__41984;
    wire N__41659;
    wire N__41656;
    wire N__41653;
    wire N__41652;
    wire N__41651;
    wire N__41650;
    wire N__41649;
    wire N__41648;
    wire N__41647;
    wire N__41646;
    wire N__41645;
    wire N__41644;
    wire N__41643;
    wire N__41642;
    wire N__41641;
    wire N__41640;
    wire N__41639;
    wire N__41608;
    wire N__41605;
    wire N__41602;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41589;
    wire N__41586;
    wire N__41581;
    wire N__41578;
    wire N__41575;
    wire N__41572;
    wire N__41569;
    wire N__41566;
    wire N__41563;
    wire N__41560;
    wire N__41557;
    wire N__41554;
    wire N__41551;
    wire N__41550;
    wire N__41549;
    wire N__41546;
    wire N__41543;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41533;
    wire N__41530;
    wire N__41527;
    wire N__41524;
    wire N__41515;
    wire N__41514;
    wire N__41513;
    wire N__41512;
    wire N__41511;
    wire N__41510;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41494;
    wire N__41491;
    wire N__41488;
    wire N__41485;
    wire N__41482;
    wire N__41475;
    wire N__41474;
    wire N__41471;
    wire N__41470;
    wire N__41467;
    wire N__41466;
    wire N__41461;
    wire N__41458;
    wire N__41455;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41437;
    wire N__41434;
    wire N__41431;
    wire N__41426;
    wire N__41421;
    wire N__41418;
    wire N__41413;
    wire N__41410;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41398;
    wire N__41395;
    wire N__41386;
    wire N__41383;
    wire N__41380;
    wire N__41377;
    wire N__41374;
    wire N__41371;
    wire N__41368;
    wire N__41365;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41355;
    wire N__41350;
    wire N__41347;
    wire N__41344;
    wire N__41341;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41323;
    wire N__41322;
    wire N__41319;
    wire N__41316;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41296;
    wire N__41295;
    wire N__41292;
    wire N__41289;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41257;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41249;
    wire N__41246;
    wire N__41243;
    wire N__41240;
    wire N__41233;
    wire N__41230;
    wire N__41227;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41214;
    wire N__41213;
    wire N__41210;
    wire N__41207;
    wire N__41204;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41185;
    wire N__41184;
    wire N__41181;
    wire N__41178;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41161;
    wire N__41160;
    wire N__41157;
    wire N__41154;
    wire N__41153;
    wire N__41152;
    wire N__41151;
    wire N__41146;
    wire N__41145;
    wire N__41142;
    wire N__41137;
    wire N__41136;
    wire N__41135;
    wire N__41134;
    wire N__41133;
    wire N__41132;
    wire N__41131;
    wire N__41130;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41097;
    wire N__41096;
    wire N__41095;
    wire N__41092;
    wire N__41085;
    wire N__41082;
    wire N__41079;
    wire N__41076;
    wire N__41069;
    wire N__41062;
    wire N__41061;
    wire N__41060;
    wire N__41053;
    wire N__41050;
    wire N__41045;
    wire N__41038;
    wire N__41035;
    wire N__41032;
    wire N__41029;
    wire N__41026;
    wire N__41023;
    wire N__41020;
    wire N__41017;
    wire N__41014;
    wire N__41011;
    wire N__41008;
    wire N__41005;
    wire N__41004;
    wire N__41001;
    wire N__40998;
    wire N__40993;
    wire N__40990;
    wire N__40987;
    wire N__40984;
    wire N__40981;
    wire N__40978;
    wire N__40975;
    wire N__40972;
    wire N__40971;
    wire N__40968;
    wire N__40967;
    wire N__40964;
    wire N__40961;
    wire N__40958;
    wire N__40955;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40929;
    wire N__40926;
    wire N__40923;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40909;
    wire N__40906;
    wire N__40903;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40891;
    wire N__40890;
    wire N__40885;
    wire N__40882;
    wire N__40881;
    wire N__40880;
    wire N__40877;
    wire N__40874;
    wire N__40871;
    wire N__40866;
    wire N__40863;
    wire N__40862;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40852;
    wire N__40849;
    wire N__40840;
    wire N__40839;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40825;
    wire N__40822;
    wire N__40819;
    wire N__40816;
    wire N__40813;
    wire N__40812;
    wire N__40809;
    wire N__40808;
    wire N__40805;
    wire N__40802;
    wire N__40799;
    wire N__40796;
    wire N__40793;
    wire N__40786;
    wire N__40785;
    wire N__40784;
    wire N__40783;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40764;
    wire N__40763;
    wire N__40760;
    wire N__40757;
    wire N__40752;
    wire N__40751;
    wire N__40748;
    wire N__40747;
    wire N__40744;
    wire N__40739;
    wire N__40736;
    wire N__40733;
    wire N__40730;
    wire N__40727;
    wire N__40726;
    wire N__40723;
    wire N__40718;
    wire N__40715;
    wire N__40710;
    wire N__40709;
    wire N__40706;
    wire N__40705;
    wire N__40702;
    wire N__40697;
    wire N__40694;
    wire N__40689;
    wire N__40686;
    wire N__40685;
    wire N__40680;
    wire N__40677;
    wire N__40672;
    wire N__40669;
    wire N__40662;
    wire N__40659;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40617;
    wire N__40614;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40572;
    wire N__40569;
    wire N__40566;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40536;
    wire N__40533;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40519;
    wire N__40516;
    wire N__40513;
    wire N__40510;
    wire N__40507;
    wire N__40504;
    wire N__40503;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40491;
    wire N__40488;
    wire N__40485;
    wire N__40480;
    wire N__40479;
    wire N__40476;
    wire N__40473;
    wire N__40470;
    wire N__40467;
    wire N__40464;
    wire N__40459;
    wire N__40458;
    wire N__40455;
    wire N__40452;
    wire N__40449;
    wire N__40444;
    wire N__40443;
    wire N__40440;
    wire N__40437;
    wire N__40436;
    wire N__40435;
    wire N__40430;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40420;
    wire N__40419;
    wire N__40416;
    wire N__40415;
    wire N__40412;
    wire N__40411;
    wire N__40408;
    wire N__40405;
    wire N__40404;
    wire N__40401;
    wire N__40398;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40388;
    wire N__40383;
    wire N__40378;
    wire N__40375;
    wire N__40372;
    wire N__40369;
    wire N__40364;
    wire N__40361;
    wire N__40358;
    wire N__40355;
    wire N__40352;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40336;
    wire N__40331;
    wire N__40328;
    wire N__40325;
    wire N__40322;
    wire N__40319;
    wire N__40312;
    wire N__40311;
    wire N__40308;
    wire N__40305;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40281;
    wire N__40280;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40254;
    wire N__40249;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40237;
    wire N__40236;
    wire N__40233;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40220;
    wire N__40215;
    wire N__40210;
    wire N__40207;
    wire N__40204;
    wire N__40201;
    wire N__40198;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40180;
    wire N__40177;
    wire N__40174;
    wire N__40171;
    wire N__40168;
    wire N__40165;
    wire N__40162;
    wire N__40159;
    wire N__40156;
    wire N__40155;
    wire N__40154;
    wire N__40153;
    wire N__40152;
    wire N__40151;
    wire N__40150;
    wire N__40149;
    wire N__40146;
    wire N__40141;
    wire N__40136;
    wire N__40133;
    wire N__40130;
    wire N__40129;
    wire N__40126;
    wire N__40123;
    wire N__40122;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40096;
    wire N__40093;
    wire N__40088;
    wire N__40085;
    wire N__40080;
    wire N__40075;
    wire N__40072;
    wire N__40069;
    wire N__40068;
    wire N__40065;
    wire N__40062;
    wire N__40061;
    wire N__40060;
    wire N__40059;
    wire N__40058;
    wire N__40053;
    wire N__40052;
    wire N__40049;
    wire N__40046;
    wire N__40043;
    wire N__40040;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40032;
    wire N__40029;
    wire N__40022;
    wire N__40019;
    wire N__40016;
    wire N__40013;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__40000;
    wire N__39995;
    wire N__39990;
    wire N__39987;
    wire N__39982;
    wire N__39979;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39965;
    wire N__39960;
    wire N__39957;
    wire N__39952;
    wire N__39949;
    wire N__39946;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39936;
    wire N__39931;
    wire N__39928;
    wire N__39927;
    wire N__39926;
    wire N__39923;
    wire N__39920;
    wire N__39917;
    wire N__39910;
    wire N__39907;
    wire N__39906;
    wire N__39905;
    wire N__39902;
    wire N__39899;
    wire N__39898;
    wire N__39897;
    wire N__39894;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39877;
    wire N__39874;
    wire N__39871;
    wire N__39870;
    wire N__39867;
    wire N__39860;
    wire N__39857;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39847;
    wire N__39844;
    wire N__39839;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39823;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39805;
    wire N__39802;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39784;
    wire N__39783;
    wire N__39782;
    wire N__39781;
    wire N__39778;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39761;
    wire N__39760;
    wire N__39757;
    wire N__39754;
    wire N__39753;
    wire N__39750;
    wire N__39745;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39729;
    wire N__39728;
    wire N__39725;
    wire N__39720;
    wire N__39717;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39698;
    wire N__39695;
    wire N__39690;
    wire N__39687;
    wire N__39686;
    wire N__39681;
    wire N__39678;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39664;
    wire N__39661;
    wire N__39658;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39634;
    wire N__39633;
    wire N__39632;
    wire N__39629;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39586;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39565;
    wire N__39564;
    wire N__39563;
    wire N__39562;
    wire N__39559;
    wire N__39556;
    wire N__39551;
    wire N__39548;
    wire N__39547;
    wire N__39544;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39527;
    wire N__39520;
    wire N__39517;
    wire N__39514;
    wire N__39511;
    wire N__39508;
    wire N__39507;
    wire N__39506;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39467;
    wire N__39462;
    wire N__39461;
    wire N__39460;
    wire N__39459;
    wire N__39456;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39431;
    wire N__39422;
    wire N__39415;
    wire N__39412;
    wire N__39409;
    wire N__39406;
    wire N__39403;
    wire N__39400;
    wire N__39397;
    wire N__39394;
    wire N__39391;
    wire N__39388;
    wire N__39385;
    wire N__39382;
    wire N__39381;
    wire N__39378;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39365;
    wire N__39364;
    wire N__39361;
    wire N__39358;
    wire N__39355;
    wire N__39352;
    wire N__39349;
    wire N__39340;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39318;
    wire N__39317;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39305;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39289;
    wire N__39286;
    wire N__39283;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39273;
    wire N__39272;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39260;
    wire N__39253;
    wire N__39250;
    wire N__39247;
    wire N__39244;
    wire N__39241;
    wire N__39238;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39228;
    wire N__39227;
    wire N__39224;
    wire N__39221;
    wire N__39218;
    wire N__39215;
    wire N__39208;
    wire N__39205;
    wire N__39202;
    wire N__39199;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39187;
    wire N__39184;
    wire N__39181;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39117;
    wire N__39114;
    wire N__39113;
    wire N__39112;
    wire N__39111;
    wire N__39110;
    wire N__39109;
    wire N__39108;
    wire N__39107;
    wire N__39106;
    wire N__39105;
    wire N__39104;
    wire N__39101;
    wire N__39100;
    wire N__39099;
    wire N__39098;
    wire N__39097;
    wire N__39094;
    wire N__39081;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39062;
    wire N__39059;
    wire N__39056;
    wire N__39051;
    wire N__39034;
    wire N__39031;
    wire N__39028;
    wire N__39025;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38995;
    wire N__38992;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38925;
    wire N__38924;
    wire N__38923;
    wire N__38922;
    wire N__38921;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38904;
    wire N__38903;
    wire N__38902;
    wire N__38895;
    wire N__38892;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38866;
    wire N__38865;
    wire N__38862;
    wire N__38861;
    wire N__38860;
    wire N__38859;
    wire N__38858;
    wire N__38855;
    wire N__38848;
    wire N__38847;
    wire N__38846;
    wire N__38843;
    wire N__38840;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38830;
    wire N__38827;
    wire N__38824;
    wire N__38819;
    wire N__38814;
    wire N__38811;
    wire N__38802;
    wire N__38797;
    wire N__38796;
    wire N__38795;
    wire N__38794;
    wire N__38793;
    wire N__38790;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38776;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38759;
    wire N__38756;
    wire N__38755;
    wire N__38748;
    wire N__38745;
    wire N__38740;
    wire N__38737;
    wire N__38734;
    wire N__38731;
    wire N__38728;
    wire N__38719;
    wire N__38718;
    wire N__38717;
    wire N__38716;
    wire N__38713;
    wire N__38710;
    wire N__38709;
    wire N__38704;
    wire N__38703;
    wire N__38702;
    wire N__38701;
    wire N__38698;
    wire N__38695;
    wire N__38692;
    wire N__38689;
    wire N__38682;
    wire N__38679;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38657;
    wire N__38650;
    wire N__38647;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38622;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38608;
    wire N__38607;
    wire N__38606;
    wire N__38605;
    wire N__38602;
    wire N__38599;
    wire N__38598;
    wire N__38597;
    wire N__38596;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38588;
    wire N__38587;
    wire N__38586;
    wire N__38581;
    wire N__38578;
    wire N__38571;
    wire N__38566;
    wire N__38563;
    wire N__38560;
    wire N__38557;
    wire N__38550;
    wire N__38545;
    wire N__38536;
    wire N__38535;
    wire N__38534;
    wire N__38533;
    wire N__38532;
    wire N__38527;
    wire N__38524;
    wire N__38519;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38491;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38479;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38461;
    wire N__38458;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38446;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38438;
    wire N__38437;
    wire N__38432;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38414;
    wire N__38413;
    wire N__38408;
    wire N__38405;
    wire N__38402;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38368;
    wire N__38365;
    wire N__38364;
    wire N__38361;
    wire N__38358;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38346;
    wire N__38343;
    wire N__38340;
    wire N__38337;
    wire N__38334;
    wire N__38331;
    wire N__38328;
    wire N__38323;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38287;
    wire N__38286;
    wire N__38285;
    wire N__38282;
    wire N__38277;
    wire N__38276;
    wire N__38275;
    wire N__38270;
    wire N__38265;
    wire N__38260;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38226;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38209;
    wire N__38206;
    wire N__38205;
    wire N__38204;
    wire N__38199;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38189;
    wire N__38188;
    wire N__38187;
    wire N__38184;
    wire N__38179;
    wire N__38178;
    wire N__38177;
    wire N__38176;
    wire N__38175;
    wire N__38174;
    wire N__38169;
    wire N__38164;
    wire N__38163;
    wire N__38152;
    wire N__38151;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38132;
    wire N__38129;
    wire N__38126;
    wire N__38121;
    wire N__38114;
    wire N__38107;
    wire N__38106;
    wire N__38105;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38097;
    wire N__38094;
    wire N__38091;
    wire N__38090;
    wire N__38087;
    wire N__38084;
    wire N__38081;
    wire N__38080;
    wire N__38079;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38069;
    wire N__38068;
    wire N__38063;
    wire N__38060;
    wire N__38057;
    wire N__38054;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38040;
    wire N__38039;
    wire N__38038;
    wire N__38037;
    wire N__38034;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37997;
    wire N__37994;
    wire N__37991;
    wire N__37986;
    wire N__37983;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37946;
    wire N__37943;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37929;
    wire N__37924;
    wire N__37921;
    wire N__37912;
    wire N__37909;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37879;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37831;
    wire N__37828;
    wire N__37825;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37804;
    wire N__37801;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37789;
    wire N__37786;
    wire N__37785;
    wire N__37782;
    wire N__37781;
    wire N__37778;
    wire N__37775;
    wire N__37772;
    wire N__37769;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37755;
    wire N__37752;
    wire N__37749;
    wire N__37748;
    wire N__37747;
    wire N__37744;
    wire N__37741;
    wire N__37740;
    wire N__37737;
    wire N__37736;
    wire N__37735;
    wire N__37734;
    wire N__37731;
    wire N__37730;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37706;
    wire N__37703;
    wire N__37700;
    wire N__37697;
    wire N__37696;
    wire N__37693;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37677;
    wire N__37674;
    wire N__37671;
    wire N__37668;
    wire N__37665;
    wire N__37662;
    wire N__37657;
    wire N__37654;
    wire N__37639;
    wire N__37636;
    wire N__37635;
    wire N__37632;
    wire N__37629;
    wire N__37624;
    wire N__37623;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37612;
    wire N__37611;
    wire N__37610;
    wire N__37609;
    wire N__37608;
    wire N__37607;
    wire N__37606;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37585;
    wire N__37584;
    wire N__37581;
    wire N__37578;
    wire N__37577;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37563;
    wire N__37562;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37549;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37530;
    wire N__37527;
    wire N__37524;
    wire N__37521;
    wire N__37514;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37496;
    wire N__37493;
    wire N__37488;
    wire N__37481;
    wire N__37478;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37464;
    wire N__37459;
    wire N__37456;
    wire N__37455;
    wire N__37452;
    wire N__37449;
    wire N__37446;
    wire N__37441;
    wire N__37438;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37427;
    wire N__37426;
    wire N__37423;
    wire N__37420;
    wire N__37417;
    wire N__37414;
    wire N__37405;
    wire N__37402;
    wire N__37399;
    wire N__37396;
    wire N__37395;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37387;
    wire N__37386;
    wire N__37383;
    wire N__37378;
    wire N__37375;
    wire N__37372;
    wire N__37369;
    wire N__37360;
    wire N__37357;
    wire N__37354;
    wire N__37351;
    wire N__37348;
    wire N__37345;
    wire N__37344;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37330;
    wire N__37329;
    wire N__37322;
    wire N__37319;
    wire N__37318;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37298;
    wire N__37291;
    wire N__37290;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37264;
    wire N__37261;
    wire N__37260;
    wire N__37259;
    wire N__37256;
    wire N__37255;
    wire N__37254;
    wire N__37253;
    wire N__37252;
    wire N__37251;
    wire N__37250;
    wire N__37245;
    wire N__37242;
    wire N__37239;
    wire N__37238;
    wire N__37237;
    wire N__37236;
    wire N__37235;
    wire N__37234;
    wire N__37233;
    wire N__37222;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37210;
    wire N__37207;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37177;
    wire N__37176;
    wire N__37173;
    wire N__37170;
    wire N__37169;
    wire N__37166;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37147;
    wire N__37142;
    wire N__37135;
    wire N__37134;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37123;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37111;
    wire N__37108;
    wire N__37105;
    wire N__37100;
    wire N__37093;
    wire N__37090;
    wire N__37087;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37063;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37038;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37027;
    wire N__37020;
    wire N__37017;
    wire N__37014;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__37002;
    wire N__37001;
    wire N__37000;
    wire N__36999;
    wire N__36996;
    wire N__36995;
    wire N__36992;
    wire N__36987;
    wire N__36980;
    wire N__36979;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36964;
    wire N__36961;
    wire N__36952;
    wire N__36949;
    wire N__36946;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36793;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36757;
    wire N__36754;
    wire N__36751;
    wire N__36748;
    wire N__36745;
    wire N__36742;
    wire N__36739;
    wire N__36736;
    wire N__36733;
    wire N__36730;
    wire N__36727;
    wire N__36724;
    wire N__36721;
    wire N__36718;
    wire N__36715;
    wire N__36712;
    wire N__36709;
    wire N__36706;
    wire N__36703;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36691;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36676;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36655;
    wire N__36652;
    wire N__36649;
    wire N__36646;
    wire N__36643;
    wire N__36640;
    wire N__36637;
    wire N__36634;
    wire N__36631;
    wire N__36628;
    wire N__36625;
    wire N__36622;
    wire N__36619;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36607;
    wire N__36604;
    wire N__36601;
    wire N__36598;
    wire N__36595;
    wire N__36594;
    wire N__36591;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36571;
    wire N__36568;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36543;
    wire N__36538;
    wire N__36535;
    wire N__36534;
    wire N__36533;
    wire N__36532;
    wire N__36531;
    wire N__36528;
    wire N__36525;
    wire N__36522;
    wire N__36519;
    wire N__36518;
    wire N__36515;
    wire N__36514;
    wire N__36513;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36492;
    wire N__36485;
    wire N__36484;
    wire N__36479;
    wire N__36478;
    wire N__36477;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36462;
    wire N__36459;
    wire N__36456;
    wire N__36445;
    wire N__36444;
    wire N__36443;
    wire N__36442;
    wire N__36439;
    wire N__36438;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36430;
    wire N__36427;
    wire N__36424;
    wire N__36421;
    wire N__36418;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36398;
    wire N__36395;
    wire N__36392;
    wire N__36379;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36369;
    wire N__36364;
    wire N__36361;
    wire N__36358;
    wire N__36355;
    wire N__36354;
    wire N__36351;
    wire N__36350;
    wire N__36347;
    wire N__36344;
    wire N__36343;
    wire N__36340;
    wire N__36337;
    wire N__36336;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36318;
    wire N__36307;
    wire N__36306;
    wire N__36301;
    wire N__36300;
    wire N__36299;
    wire N__36298;
    wire N__36295;
    wire N__36288;
    wire N__36287;
    wire N__36282;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36272;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36260;
    wire N__36255;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36243;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36235;
    wire N__36232;
    wire N__36227;
    wire N__36226;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36214;
    wire N__36211;
    wire N__36210;
    wire N__36207;
    wire N__36200;
    wire N__36197;
    wire N__36196;
    wire N__36195;
    wire N__36192;
    wire N__36189;
    wire N__36186;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36170;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36156;
    wire N__36155;
    wire N__36154;
    wire N__36153;
    wire N__36152;
    wire N__36149;
    wire N__36146;
    wire N__36141;
    wire N__36138;
    wire N__36135;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36114;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36101;
    wire N__36100;
    wire N__36099;
    wire N__36096;
    wire N__36091;
    wire N__36088;
    wire N__36085;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36064;
    wire N__36061;
    wire N__36058;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__36000;
    wire N__35995;
    wire N__35992;
    wire N__35989;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35977;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35965;
    wire N__35964;
    wire N__35961;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35950;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35937;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35918;
    wire N__35915;
    wire N__35914;
    wire N__35911;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35886;
    wire N__35883;
    wire N__35878;
    wire N__35875;
    wire N__35868;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35851;
    wire N__35848;
    wire N__35847;
    wire N__35846;
    wire N__35845;
    wire N__35842;
    wire N__35841;
    wire N__35840;
    wire N__35839;
    wire N__35834;
    wire N__35831;
    wire N__35830;
    wire N__35827;
    wire N__35822;
    wire N__35819;
    wire N__35814;
    wire N__35811;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35793;
    wire N__35788;
    wire N__35785;
    wire N__35784;
    wire N__35783;
    wire N__35782;
    wire N__35781;
    wire N__35778;
    wire N__35777;
    wire N__35774;
    wire N__35773;
    wire N__35770;
    wire N__35767;
    wire N__35764;
    wire N__35763;
    wire N__35760;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35748;
    wire N__35743;
    wire N__35740;
    wire N__35733;
    wire N__35726;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35712;
    wire N__35711;
    wire N__35710;
    wire N__35709;
    wire N__35706;
    wire N__35705;
    wire N__35698;
    wire N__35693;
    wire N__35690;
    wire N__35685;
    wire N__35684;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35665;
    wire N__35664;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35656;
    wire N__35653;
    wire N__35648;
    wire N__35645;
    wire N__35642;
    wire N__35637;
    wire N__35634;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35617;
    wire N__35616;
    wire N__35615;
    wire N__35612;
    wire N__35611;
    wire N__35610;
    wire N__35609;
    wire N__35608;
    wire N__35605;
    wire N__35604;
    wire N__35603;
    wire N__35602;
    wire N__35595;
    wire N__35592;
    wire N__35587;
    wire N__35582;
    wire N__35577;
    wire N__35566;
    wire N__35563;
    wire N__35560;
    wire N__35557;
    wire N__35554;
    wire N__35553;
    wire N__35552;
    wire N__35549;
    wire N__35548;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35520;
    wire N__35519;
    wire N__35518;
    wire N__35517;
    wire N__35516;
    wire N__35515;
    wire N__35514;
    wire N__35511;
    wire N__35508;
    wire N__35505;
    wire N__35498;
    wire N__35495;
    wire N__35492;
    wire N__35491;
    wire N__35490;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35472;
    wire N__35469;
    wire N__35466;
    wire N__35465;
    wire N__35464;
    wire N__35461;
    wire N__35460;
    wire N__35453;
    wire N__35448;
    wire N__35443;
    wire N__35440;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35426;
    wire N__35423;
    wire N__35410;
    wire N__35409;
    wire N__35408;
    wire N__35407;
    wire N__35406;
    wire N__35405;
    wire N__35402;
    wire N__35401;
    wire N__35400;
    wire N__35399;
    wire N__35398;
    wire N__35393;
    wire N__35392;
    wire N__35387;
    wire N__35386;
    wire N__35385;
    wire N__35384;
    wire N__35381;
    wire N__35380;
    wire N__35377;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35361;
    wire N__35358;
    wire N__35353;
    wire N__35346;
    wire N__35329;
    wire N__35326;
    wire N__35323;
    wire N__35322;
    wire N__35321;
    wire N__35320;
    wire N__35319;
    wire N__35318;
    wire N__35317;
    wire N__35316;
    wire N__35315;
    wire N__35314;
    wire N__35311;
    wire N__35308;
    wire N__35307;
    wire N__35306;
    wire N__35305;
    wire N__35304;
    wire N__35303;
    wire N__35302;
    wire N__35301;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35286;
    wire N__35279;
    wire N__35276;
    wire N__35271;
    wire N__35266;
    wire N__35263;
    wire N__35260;
    wire N__35257;
    wire N__35252;
    wire N__35249;
    wire N__35248;
    wire N__35245;
    wire N__35242;
    wire N__35241;
    wire N__35240;
    wire N__35237;
    wire N__35232;
    wire N__35229;
    wire N__35220;
    wire N__35219;
    wire N__35216;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35197;
    wire N__35190;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35170;
    wire N__35155;
    wire N__35154;
    wire N__35153;
    wire N__35152;
    wire N__35151;
    wire N__35150;
    wire N__35147;
    wire N__35146;
    wire N__35143;
    wire N__35142;
    wire N__35141;
    wire N__35138;
    wire N__35137;
    wire N__35136;
    wire N__35135;
    wire N__35134;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35115;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35100;
    wire N__35099;
    wire N__35096;
    wire N__35093;
    wire N__35090;
    wire N__35089;
    wire N__35086;
    wire N__35079;
    wire N__35076;
    wire N__35075;
    wire N__35072;
    wire N__35065;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35046;
    wire N__35039;
    wire N__35036;
    wire N__35029;
    wire N__35014;
    wire N__35013;
    wire N__35012;
    wire N__35009;
    wire N__35006;
    wire N__35005;
    wire N__35004;
    wire N__35001;
    wire N__35000;
    wire N__34999;
    wire N__34996;
    wire N__34995;
    wire N__34994;
    wire N__34993;
    wire N__34992;
    wire N__34991;
    wire N__34990;
    wire N__34987;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34973;
    wire N__34972;
    wire N__34971;
    wire N__34968;
    wire N__34967;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34955;
    wire N__34948;
    wire N__34947;
    wire N__34946;
    wire N__34945;
    wire N__34944;
    wire N__34943;
    wire N__34942;
    wire N__34939;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34924;
    wire N__34921;
    wire N__34916;
    wire N__34913;
    wire N__34908;
    wire N__34901;
    wire N__34898;
    wire N__34897;
    wire N__34894;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34881;
    wire N__34880;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34865;
    wire N__34858;
    wire N__34855;
    wire N__34846;
    wire N__34843;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34831;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34804;
    wire N__34801;
    wire N__34796;
    wire N__34787;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34751;
    wire N__34750;
    wire N__34749;
    wire N__34748;
    wire N__34747;
    wire N__34746;
    wire N__34745;
    wire N__34744;
    wire N__34739;
    wire N__34736;
    wire N__34735;
    wire N__34732;
    wire N__34729;
    wire N__34726;
    wire N__34723;
    wire N__34720;
    wire N__34717;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34706;
    wire N__34705;
    wire N__34704;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34692;
    wire N__34685;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34662;
    wire N__34651;
    wire N__34648;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34597;
    wire N__34594;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34579;
    wire N__34578;
    wire N__34577;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34566;
    wire N__34565;
    wire N__34562;
    wire N__34557;
    wire N__34554;
    wire N__34553;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34498;
    wire N__34493;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34469;
    wire N__34464;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34454;
    wire N__34451;
    wire N__34448;
    wire N__34445;
    wire N__34438;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34430;
    wire N__34427;
    wire N__34424;
    wire N__34421;
    wire N__34418;
    wire N__34413;
    wire N__34408;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34374;
    wire N__34371;
    wire N__34370;
    wire N__34369;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34357;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34341;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34321;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34285;
    wire N__34284;
    wire N__34281;
    wire N__34278;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34252;
    wire N__34251;
    wire N__34250;
    wire N__34249;
    wire N__34248;
    wire N__34247;
    wire N__34246;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34221;
    wire N__34220;
    wire N__34219;
    wire N__34218;
    wire N__34217;
    wire N__34216;
    wire N__34215;
    wire N__34214;
    wire N__34211;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34141;
    wire N__34138;
    wire N__34137;
    wire N__34136;
    wire N__34133;
    wire N__34132;
    wire N__34131;
    wire N__34130;
    wire N__34127;
    wire N__34126;
    wire N__34125;
    wire N__34124;
    wire N__34123;
    wire N__34120;
    wire N__34119;
    wire N__34118;
    wire N__34115;
    wire N__34110;
    wire N__34101;
    wire N__34098;
    wire N__34095;
    wire N__34088;
    wire N__34075;
    wire N__34074;
    wire N__34073;
    wire N__34072;
    wire N__34071;
    wire N__34070;
    wire N__34069;
    wire N__34068;
    wire N__34061;
    wire N__34058;
    wire N__34053;
    wire N__34048;
    wire N__34039;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34012;
    wire N__34009;
    wire N__34006;
    wire N__34003;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33943;
    wire N__33940;
    wire N__33937;
    wire N__33934;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33891;
    wire N__33890;
    wire N__33887;
    wire N__33886;
    wire N__33885;
    wire N__33882;
    wire N__33881;
    wire N__33880;
    wire N__33877;
    wire N__33876;
    wire N__33873;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33860;
    wire N__33857;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33814;
    wire N__33813;
    wire N__33806;
    wire N__33801;
    wire N__33798;
    wire N__33795;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33773;
    wire N__33770;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33754;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33740;
    wire N__33737;
    wire N__33732;
    wire N__33729;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33708;
    wire N__33701;
    wire N__33700;
    wire N__33697;
    wire N__33692;
    wire N__33689;
    wire N__33682;
    wire N__33679;
    wire N__33678;
    wire N__33675;
    wire N__33674;
    wire N__33673;
    wire N__33670;
    wire N__33669;
    wire N__33666;
    wire N__33663;
    wire N__33662;
    wire N__33659;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33651;
    wire N__33650;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33620;
    wire N__33617;
    wire N__33616;
    wire N__33611;
    wire N__33608;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33597;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33549;
    wire N__33546;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33500;
    wire N__33497;
    wire N__33492;
    wire N__33483;
    wire N__33482;
    wire N__33479;
    wire N__33474;
    wire N__33469;
    wire N__33466;
    wire N__33457;
    wire N__33454;
    wire N__33453;
    wire N__33452;
    wire N__33449;
    wire N__33448;
    wire N__33445;
    wire N__33444;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33434;
    wire N__33433;
    wire N__33432;
    wire N__33431;
    wire N__33430;
    wire N__33427;
    wire N__33424;
    wire N__33423;
    wire N__33420;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33403;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33386;
    wire N__33383;
    wire N__33380;
    wire N__33373;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33299;
    wire N__33296;
    wire N__33293;
    wire N__33286;
    wire N__33281;
    wire N__33276;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33264;
    wire N__33261;
    wire N__33254;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33236;
    wire N__33233;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33217;
    wire N__33216;
    wire N__33215;
    wire N__33214;
    wire N__33213;
    wire N__33212;
    wire N__33211;
    wire N__33210;
    wire N__33209;
    wire N__33208;
    wire N__33207;
    wire N__33206;
    wire N__33205;
    wire N__33204;
    wire N__33195;
    wire N__33186;
    wire N__33181;
    wire N__33172;
    wire N__33171;
    wire N__33170;
    wire N__33165;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33128;
    wire N__33125;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33090;
    wire N__33089;
    wire N__33088;
    wire N__33087;
    wire N__33084;
    wire N__33081;
    wire N__33076;
    wire N__33075;
    wire N__33074;
    wire N__33073;
    wire N__33070;
    wire N__33063;
    wire N__33056;
    wire N__33053;
    wire N__33052;
    wire N__33051;
    wire N__33048;
    wire N__33043;
    wire N__33038;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33021;
    wire N__33020;
    wire N__33019;
    wire N__33016;
    wire N__33015;
    wire N__33014;
    wire N__33013;
    wire N__33008;
    wire N__33005;
    wire N__33000;
    wire N__32995;
    wire N__32990;
    wire N__32989;
    wire N__32988;
    wire N__32987;
    wire N__32982;
    wire N__32981;
    wire N__32980;
    wire N__32977;
    wire N__32970;
    wire N__32967;
    wire N__32962;
    wire N__32953;
    wire N__32950;
    wire N__32947;
    wire N__32944;
    wire N__32943;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32935;
    wire N__32934;
    wire N__32933;
    wire N__32932;
    wire N__32929;
    wire N__32928;
    wire N__32927;
    wire N__32924;
    wire N__32921;
    wire N__32916;
    wire N__32913;
    wire N__32908;
    wire N__32903;
    wire N__32890;
    wire N__32887;
    wire N__32884;
    wire N__32881;
    wire N__32878;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32856;
    wire N__32853;
    wire N__32850;
    wire N__32845;
    wire N__32844;
    wire N__32843;
    wire N__32840;
    wire N__32839;
    wire N__32838;
    wire N__32837;
    wire N__32834;
    wire N__32831;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32816;
    wire N__32815;
    wire N__32812;
    wire N__32809;
    wire N__32806;
    wire N__32803;
    wire N__32800;
    wire N__32797;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32783;
    wire N__32782;
    wire N__32779;
    wire N__32776;
    wire N__32773;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32761;
    wire N__32758;
    wire N__32755;
    wire N__32752;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32742;
    wire N__32735;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32702;
    wire N__32697;
    wire N__32694;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32673;
    wire N__32668;
    wire N__32665;
    wire N__32662;
    wire N__32661;
    wire N__32656;
    wire N__32651;
    wire N__32648;
    wire N__32641;
    wire N__32638;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32634;
    wire N__32633;
    wire N__32632;
    wire N__32631;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32623;
    wire N__32620;
    wire N__32617;
    wire N__32614;
    wire N__32613;
    wire N__32610;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32602;
    wire N__32601;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32550;
    wire N__32547;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32511;
    wire N__32508;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32487;
    wire N__32482;
    wire N__32477;
    wire N__32474;
    wire N__32471;
    wire N__32466;
    wire N__32459;
    wire N__32456;
    wire N__32453;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32441;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32425;
    wire N__32422;
    wire N__32419;
    wire N__32416;
    wire N__32411;
    wire N__32398;
    wire N__32395;
    wire N__32392;
    wire N__32391;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32381;
    wire N__32380;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32372;
    wire N__32369;
    wire N__32366;
    wire N__32365;
    wire N__32362;
    wire N__32361;
    wire N__32360;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32333;
    wire N__32332;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32313;
    wire N__32310;
    wire N__32307;
    wire N__32304;
    wire N__32301;
    wire N__32298;
    wire N__32297;
    wire N__32296;
    wire N__32293;
    wire N__32290;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32259;
    wire N__32254;
    wire N__32249;
    wire N__32246;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32227;
    wire N__32222;
    wire N__32215;
    wire N__32212;
    wire N__32211;
    wire N__32208;
    wire N__32201;
    wire N__32198;
    wire N__32191;
    wire N__32188;
    wire N__32187;
    wire N__32184;
    wire N__32183;
    wire N__32182;
    wire N__32179;
    wire N__32176;
    wire N__32173;
    wire N__32172;
    wire N__32171;
    wire N__32170;
    wire N__32167;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32150;
    wire N__32149;
    wire N__32146;
    wire N__32143;
    wire N__32140;
    wire N__32139;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32107;
    wire N__32104;
    wire N__32101;
    wire N__32100;
    wire N__32099;
    wire N__32096;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32068;
    wire N__32065;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32055;
    wire N__32050;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32028;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32009;
    wire N__32002;
    wire N__31999;
    wire N__31998;
    wire N__31995;
    wire N__31990;
    wire N__31987;
    wire N__31984;
    wire N__31975;
    wire N__31972;
    wire N__31971;
    wire N__31970;
    wire N__31967;
    wire N__31966;
    wire N__31963;
    wire N__31962;
    wire N__31961;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31945;
    wire N__31942;
    wire N__31941;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31925;
    wire N__31922;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31911;
    wire N__31910;
    wire N__31909;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31888;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31869;
    wire N__31866;
    wire N__31861;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31830;
    wire N__31825;
    wire N__31820;
    wire N__31817;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31792;
    wire N__31783;
    wire N__31780;
    wire N__31779;
    wire N__31776;
    wire N__31769;
    wire N__31766;
    wire N__31759;
    wire N__31756;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31748;
    wire N__31747;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31736;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31728;
    wire N__31727;
    wire N__31724;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31714;
    wire N__31713;
    wire N__31712;
    wire N__31709;
    wire N__31708;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31694;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31678;
    wire N__31675;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31606;
    wire N__31601;
    wire N__31596;
    wire N__31593;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31581;
    wire N__31576;
    wire N__31573;
    wire N__31568;
    wire N__31563;
    wire N__31560;
    wire N__31549;
    wire N__31546;
    wire N__31545;
    wire N__31544;
    wire N__31543;
    wire N__31540;
    wire N__31539;
    wire N__31538;
    wire N__31535;
    wire N__31534;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31526;
    wire N__31525;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31515;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31493;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31476;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31460;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31444;
    wire N__31441;
    wire N__31438;
    wire N__31435;
    wire N__31432;
    wire N__31425;
    wire N__31424;
    wire N__31417;
    wire N__31414;
    wire N__31411;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31385;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31371;
    wire N__31366;
    wire N__31361;
    wire N__31358;
    wire N__31351;
    wire N__31348;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31340;
    wire N__31339;
    wire N__31338;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31324;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31316;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31296;
    wire N__31295;
    wire N__31292;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31282;
    wire N__31277;
    wire N__31274;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31242;
    wire N__31241;
    wire N__31236;
    wire N__31229;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31213;
    wire N__31210;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31191;
    wire N__31188;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31163;
    wire N__31160;
    wire N__31159;
    wire N__31156;
    wire N__31151;
    wire N__31148;
    wire N__31141;
    wire N__31138;
    wire N__31137;
    wire N__31132;
    wire N__31129;
    wire N__31126;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31089;
    wire N__31088;
    wire N__31085;
    wire N__31080;
    wire N__31079;
    wire N__31076;
    wire N__31075;
    wire N__31072;
    wire N__31069;
    wire N__31068;
    wire N__31067;
    wire N__31066;
    wire N__31065;
    wire N__31064;
    wire N__31063;
    wire N__31060;
    wire N__31059;
    wire N__31056;
    wire N__31055;
    wire N__31054;
    wire N__31049;
    wire N__31040;
    wire N__31035;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31020;
    wire N__31017;
    wire N__31012;
    wire N__31009;
    wire N__30994;
    wire N__30991;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30973;
    wire N__30970;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30955;
    wire N__30952;
    wire N__30949;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30929;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30918;
    wire N__30915;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30888;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30837;
    wire N__30836;
    wire N__30835;
    wire N__30834;
    wire N__30833;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30792;
    wire N__30791;
    wire N__30790;
    wire N__30785;
    wire N__30780;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30730;
    wire N__30727;
    wire N__30726;
    wire N__30725;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30700;
    wire N__30699;
    wire N__30694;
    wire N__30693;
    wire N__30692;
    wire N__30689;
    wire N__30688;
    wire N__30687;
    wire N__30686;
    wire N__30685;
    wire N__30684;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30670;
    wire N__30669;
    wire N__30664;
    wire N__30661;
    wire N__30656;
    wire N__30653;
    wire N__30652;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30638;
    wire N__30637;
    wire N__30634;
    wire N__30627;
    wire N__30624;
    wire N__30619;
    wire N__30610;
    wire N__30605;
    wire N__30600;
    wire N__30589;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30571;
    wire N__30568;
    wire N__30567;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30548;
    wire N__30541;
    wire N__30540;
    wire N__30539;
    wire N__30536;
    wire N__30535;
    wire N__30534;
    wire N__30533;
    wire N__30532;
    wire N__30527;
    wire N__30524;
    wire N__30521;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30503;
    wire N__30502;
    wire N__30501;
    wire N__30498;
    wire N__30487;
    wire N__30482;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30468;
    wire N__30467;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30459;
    wire N__30458;
    wire N__30457;
    wire N__30456;
    wire N__30455;
    wire N__30454;
    wire N__30453;
    wire N__30452;
    wire N__30451;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30429;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30421;
    wire N__30420;
    wire N__30415;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30398;
    wire N__30393;
    wire N__30390;
    wire N__30385;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30356;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30315;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30297;
    wire N__30296;
    wire N__30293;
    wire N__30288;
    wire N__30283;
    wire N__30280;
    wire N__30277;
    wire N__30274;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30240;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30173;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30157;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30108;
    wire N__30107;
    wire N__30104;
    wire N__30103;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30043;
    wire N__30040;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30030;
    wire N__30029;
    wire N__30028;
    wire N__30025;
    wire N__30020;
    wire N__30019;
    wire N__30018;
    wire N__30017;
    wire N__30016;
    wire N__30013;
    wire N__30008;
    wire N__30003;
    wire N__29998;
    wire N__29989;
    wire N__29988;
    wire N__29987;
    wire N__29984;
    wire N__29983;
    wire N__29982;
    wire N__29981;
    wire N__29980;
    wire N__29979;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29964;
    wire N__29959;
    wire N__29954;
    wire N__29951;
    wire N__29938;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29930;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29912;
    wire N__29909;
    wire N__29902;
    wire N__29899;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29886;
    wire N__29881;
    wire N__29880;
    wire N__29877;
    wire N__29876;
    wire N__29873;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29851;
    wire N__29850;
    wire N__29849;
    wire N__29844;
    wire N__29843;
    wire N__29842;
    wire N__29839;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29831;
    wire N__29828;
    wire N__29823;
    wire N__29818;
    wire N__29815;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29788;
    wire N__29785;
    wire N__29782;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29766;
    wire N__29765;
    wire N__29764;
    wire N__29761;
    wire N__29760;
    wire N__29757;
    wire N__29756;
    wire N__29755;
    wire N__29754;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29737;
    wire N__29730;
    wire N__29719;
    wire N__29718;
    wire N__29717;
    wire N__29716;
    wire N__29715;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29707;
    wire N__29706;
    wire N__29705;
    wire N__29704;
    wire N__29703;
    wire N__29698;
    wire N__29693;
    wire N__29690;
    wire N__29683;
    wire N__29676;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29647;
    wire N__29644;
    wire N__29643;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29635;
    wire N__29632;
    wire N__29627;
    wire N__29626;
    wire N__29623;
    wire N__29622;
    wire N__29621;
    wire N__29620;
    wire N__29619;
    wire N__29618;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29602;
    wire N__29599;
    wire N__29594;
    wire N__29591;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29571;
    wire N__29570;
    wire N__29569;
    wire N__29566;
    wire N__29559;
    wire N__29558;
    wire N__29557;
    wire N__29554;
    wire N__29551;
    wire N__29546;
    wire N__29539;
    wire N__29536;
    wire N__29533;
    wire N__29532;
    wire N__29531;
    wire N__29528;
    wire N__29527;
    wire N__29524;
    wire N__29523;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29509;
    wire N__29506;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29490;
    wire N__29489;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29481;
    wire N__29480;
    wire N__29477;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29463;
    wire N__29458;
    wire N__29449;
    wire N__29446;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29428;
    wire N__29427;
    wire N__29424;
    wire N__29423;
    wire N__29422;
    wire N__29419;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29411;
    wire N__29408;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29376;
    wire N__29375;
    wire N__29370;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29348;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29314;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29289;
    wire N__29286;
    wire N__29285;
    wire N__29282;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29271;
    wire N__29268;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29248;
    wire N__29245;
    wire N__29244;
    wire N__29241;
    wire N__29240;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29223;
    wire N__29222;
    wire N__29221;
    wire N__29216;
    wire N__29211;
    wire N__29206;
    wire N__29205;
    wire N__29202;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29194;
    wire N__29191;
    wire N__29190;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29171;
    wire N__29168;
    wire N__29161;
    wire N__29158;
    wire N__29155;
    wire N__29152;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29144;
    wire N__29143;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29128;
    wire N__29121;
    wire N__29116;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29082;
    wire N__29081;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29069;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29053;
    wire N__29052;
    wire N__29047;
    wire N__29046;
    wire N__29043;
    wire N__29042;
    wire N__29041;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29007;
    wire N__29004;
    wire N__29003;
    wire N__29002;
    wire N__28999;
    wire N__28992;
    wire N__28987;
    wire N__28986;
    wire N__28983;
    wire N__28982;
    wire N__28981;
    wire N__28978;
    wire N__28977;
    wire N__28972;
    wire N__28969;
    wire N__28964;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28937;
    wire N__28936;
    wire N__28935;
    wire N__28932;
    wire N__28931;
    wire N__28930;
    wire N__28929;
    wire N__28928;
    wire N__28925;
    wire N__28918;
    wire N__28915;
    wire N__28910;
    wire N__28909;
    wire N__28906;
    wire N__28905;
    wire N__28904;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28880;
    wire N__28875;
    wire N__28858;
    wire N__28857;
    wire N__28856;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28844;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28785;
    wire N__28784;
    wire N__28781;
    wire N__28776;
    wire N__28771;
    wire N__28770;
    wire N__28769;
    wire N__28768;
    wire N__28767;
    wire N__28766;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28750;
    wire N__28749;
    wire N__28748;
    wire N__28745;
    wire N__28742;
    wire N__28737;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28717;
    wire N__28714;
    wire N__28713;
    wire N__28712;
    wire N__28711;
    wire N__28706;
    wire N__28705;
    wire N__28704;
    wire N__28703;
    wire N__28702;
    wire N__28697;
    wire N__28694;
    wire N__28693;
    wire N__28690;
    wire N__28683;
    wire N__28678;
    wire N__28675;
    wire N__28666;
    wire N__28665;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28651;
    wire N__28650;
    wire N__28649;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire N__28634;
    wire N__28629;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28540;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28528;
    wire N__28525;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28517;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28453;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28438;
    wire N__28435;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28425;
    wire N__28424;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28392;
    wire N__28387;
    wire N__28384;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28336;
    wire N__28333;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28293;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28275;
    wire N__28270;
    wire N__28269;
    wire N__28264;
    wire N__28261;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28253;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28230;
    wire N__28229;
    wire N__28224;
    wire N__28221;
    wire N__28216;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28201;
    wire N__28200;
    wire N__28197;
    wire N__28196;
    wire N__28195;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28180;
    wire N__28171;
    wire N__28168;
    wire N__28167;
    wire N__28166;
    wire N__28165;
    wire N__28164;
    wire N__28163;
    wire N__28162;
    wire N__28157;
    wire N__28150;
    wire N__28145;
    wire N__28138;
    wire N__28135;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28115;
    wire N__28114;
    wire N__28109;
    wire N__28106;
    wire N__28105;
    wire N__28102;
    wire N__28097;
    wire N__28094;
    wire N__28093;
    wire N__28090;
    wire N__28085;
    wire N__28082;
    wire N__28081;
    wire N__28080;
    wire N__28077;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28047;
    wire N__28042;
    wire N__28039;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28031;
    wire N__28030;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__27994;
    wire N__27991;
    wire N__27990;
    wire N__27989;
    wire N__27986;
    wire N__27983;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27971;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27957;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27949;
    wire N__27946;
    wire N__27945;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27915;
    wire N__27914;
    wire N__27911;
    wire N__27910;
    wire N__27909;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27873;
    wire N__27872;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27860;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27817;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27709;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27681;
    wire N__27680;
    wire N__27679;
    wire N__27676;
    wire N__27675;
    wire N__27672;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27647;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27627;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27615;
    wire N__27614;
    wire N__27613;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27592;
    wire N__27589;
    wire N__27588;
    wire N__27587;
    wire N__27586;
    wire N__27585;
    wire N__27582;
    wire N__27577;
    wire N__27572;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27550;
    wire N__27549;
    wire N__27548;
    wire N__27547;
    wire N__27546;
    wire N__27545;
    wire N__27544;
    wire N__27543;
    wire N__27542;
    wire N__27541;
    wire N__27540;
    wire N__27539;
    wire N__27538;
    wire N__27537;
    wire N__27532;
    wire N__27521;
    wire N__27506;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27490;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27482;
    wire N__27481;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27467;
    wire N__27466;
    wire N__27465;
    wire N__27464;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27445;
    wire N__27436;
    wire N__27433;
    wire N__27432;
    wire N__27431;
    wire N__27428;
    wire N__27427;
    wire N__27426;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27411;
    wire N__27408;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27384;
    wire N__27383;
    wire N__27382;
    wire N__27379;
    wire N__27376;
    wire N__27371;
    wire N__27364;
    wire N__27361;
    wire N__27360;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27345;
    wire N__27344;
    wire N__27343;
    wire N__27336;
    wire N__27335;
    wire N__27334;
    wire N__27333;
    wire N__27330;
    wire N__27329;
    wire N__27328;
    wire N__27327;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27313;
    wire N__27312;
    wire N__27309;
    wire N__27304;
    wire N__27299;
    wire N__27298;
    wire N__27297;
    wire N__27296;
    wire N__27295;
    wire N__27294;
    wire N__27293;
    wire N__27292;
    wire N__27291;
    wire N__27286;
    wire N__27281;
    wire N__27280;
    wire N__27279;
    wire N__27274;
    wire N__27271;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27255;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27235;
    wire N__27230;
    wire N__27225;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27117;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27103;
    wire N__27102;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27083;
    wire N__27082;
    wire N__27075;
    wire N__27074;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27062;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27047;
    wire N__27042;
    wire N__27037;
    wire N__27028;
    wire N__27027;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27017;
    wire N__27010;
    wire N__27007;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26988;
    wire N__26985;
    wire N__26982;
    wire N__26981;
    wire N__26978;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26956;
    wire N__26953;
    wire N__26944;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26925;
    wire N__26924;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26897;
    wire N__26890;
    wire N__26889;
    wire N__26888;
    wire N__26887;
    wire N__26884;
    wire N__26881;
    wire N__26880;
    wire N__26877;
    wire N__26876;
    wire N__26875;
    wire N__26870;
    wire N__26867;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26845;
    wire N__26844;
    wire N__26843;
    wire N__26842;
    wire N__26841;
    wire N__26840;
    wire N__26839;
    wire N__26838;
    wire N__26835;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26810;
    wire N__26797;
    wire N__26796;
    wire N__26793;
    wire N__26792;
    wire N__26791;
    wire N__26790;
    wire N__26789;
    wire N__26786;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26766;
    wire N__26761;
    wire N__26760;
    wire N__26759;
    wire N__26758;
    wire N__26757;
    wire N__26754;
    wire N__26749;
    wire N__26748;
    wire N__26747;
    wire N__26744;
    wire N__26741;
    wire N__26740;
    wire N__26739;
    wire N__26738;
    wire N__26737;
    wire N__26736;
    wire N__26735;
    wire N__26734;
    wire N__26733;
    wire N__26732;
    wire N__26731;
    wire N__26730;
    wire N__26729;
    wire N__26728;
    wire N__26727;
    wire N__26726;
    wire N__26725;
    wire N__26724;
    wire N__26723;
    wire N__26722;
    wire N__26721;
    wire N__26720;
    wire N__26719;
    wire N__26718;
    wire N__26713;
    wire N__26708;
    wire N__26703;
    wire N__26698;
    wire N__26689;
    wire N__26680;
    wire N__26675;
    wire N__26674;
    wire N__26667;
    wire N__26658;
    wire N__26649;
    wire N__26644;
    wire N__26643;
    wire N__26642;
    wire N__26641;
    wire N__26638;
    wire N__26633;
    wire N__26628;
    wire N__26625;
    wire N__26618;
    wire N__26615;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26599;
    wire N__26594;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26559;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26544;
    wire N__26541;
    wire N__26538;
    wire N__26535;
    wire N__26532;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26498;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26448;
    wire N__26447;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26431;
    wire N__26428;
    wire N__26427;
    wire N__26426;
    wire N__26423;
    wire N__26418;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26403;
    wire N__26400;
    wire N__26399;
    wire N__26398;
    wire N__26397;
    wire N__26394;
    wire N__26391;
    wire N__26388;
    wire N__26383;
    wire N__26380;
    wire N__26377;
    wire N__26368;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26341;
    wire N__26338;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26287;
    wire N__26284;
    wire N__26283;
    wire N__26280;
    wire N__26277;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26265;
    wire N__26262;
    wire N__26259;
    wire N__26254;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26236;
    wire N__26235;
    wire N__26232;
    wire N__26229;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26203;
    wire N__26200;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26173;
    wire N__26170;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26143;
    wire N__26142;
    wire N__26141;
    wire N__26138;
    wire N__26137;
    wire N__26136;
    wire N__26135;
    wire N__26132;
    wire N__26131;
    wire N__26130;
    wire N__26129;
    wire N__26128;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26118;
    wire N__26117;
    wire N__26116;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26106;
    wire N__26103;
    wire N__26098;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26086;
    wire N__26081;
    wire N__26078;
    wire N__26077;
    wire N__26076;
    wire N__26075;
    wire N__26074;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26028;
    wire N__26025;
    wire N__26018;
    wire N__26013;
    wire N__26010;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25942;
    wire N__25939;
    wire N__25938;
    wire N__25933;
    wire N__25932;
    wire N__25931;
    wire N__25928;
    wire N__25923;
    wire N__25918;
    wire N__25917;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25906;
    wire N__25899;
    wire N__25896;
    wire N__25891;
    wire N__25888;
    wire N__25887;
    wire N__25886;
    wire N__25885;
    wire N__25880;
    wire N__25879;
    wire N__25876;
    wire N__25873;
    wire N__25870;
    wire N__25863;
    wire N__25860;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25798;
    wire N__25795;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25737;
    wire N__25734;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25717;
    wire N__25716;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25686;
    wire N__25685;
    wire N__25682;
    wire N__25681;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25644;
    wire N__25641;
    wire N__25638;
    wire N__25633;
    wire N__25632;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25605;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25588;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25551;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25533;
    wire N__25528;
    wire N__25527;
    wire N__25526;
    wire N__25525;
    wire N__25524;
    wire N__25523;
    wire N__25520;
    wire N__25509;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25482;
    wire N__25481;
    wire N__25480;
    wire N__25479;
    wire N__25478;
    wire N__25475;
    wire N__25464;
    wire N__25463;
    wire N__25462;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25450;
    wire N__25441;
    wire N__25440;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25390;
    wire N__25389;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25366;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25358;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25327;
    wire N__25324;
    wire N__25321;
    wire N__25318;
    wire N__25315;
    wire N__25312;
    wire N__25311;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25263;
    wire N__25262;
    wire N__25261;
    wire N__25260;
    wire N__25259;
    wire N__25256;
    wire N__25255;
    wire N__25252;
    wire N__25251;
    wire N__25248;
    wire N__25247;
    wire N__25244;
    wire N__25243;
    wire N__25240;
    wire N__25237;
    wire N__25236;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25228;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25220;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25206;
    wire N__25205;
    wire N__25204;
    wire N__25203;
    wire N__25200;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25177;
    wire N__25176;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25164;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25142;
    wire N__25139;
    wire N__25138;
    wire N__25135;
    wire N__25134;
    wire N__25133;
    wire N__25126;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25110;
    wire N__25103;
    wire N__25100;
    wire N__25093;
    wire N__25088;
    wire N__25085;
    wire N__25084;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25076;
    wire N__25075;
    wire N__25074;
    wire N__25073;
    wire N__25072;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25061;
    wire N__25060;
    wire N__25059;
    wire N__25050;
    wire N__25047;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25025;
    wire N__25022;
    wire N__25021;
    wire N__25020;
    wire N__25019;
    wire N__25018;
    wire N__25017;
    wire N__25014;
    wire N__25013;
    wire N__25010;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24999;
    wire N__24992;
    wire N__24991;
    wire N__24988;
    wire N__24987;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24958;
    wire N__24955;
    wire N__24954;
    wire N__24951;
    wire N__24950;
    wire N__24947;
    wire N__24934;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24907;
    wire N__24906;
    wire N__24899;
    wire N__24896;
    wire N__24891;
    wire N__24890;
    wire N__24889;
    wire N__24888;
    wire N__24887;
    wire N__24886;
    wire N__24871;
    wire N__24870;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24856;
    wire N__24853;
    wire N__24852;
    wire N__24847;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24833;
    wire N__24830;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24796;
    wire N__24791;
    wire N__24788;
    wire N__24779;
    wire N__24776;
    wire N__24771;
    wire N__24766;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24743;
    wire N__24738;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24707;
    wire N__24704;
    wire N__24697;
    wire N__24694;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24682;
    wire N__24681;
    wire N__24680;
    wire N__24679;
    wire N__24678;
    wire N__24677;
    wire N__24676;
    wire N__24675;
    wire N__24674;
    wire N__24671;
    wire N__24670;
    wire N__24669;
    wire N__24668;
    wire N__24667;
    wire N__24666;
    wire N__24665;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24644;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24615;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24600;
    wire N__24597;
    wire N__24588;
    wire N__24583;
    wire N__24582;
    wire N__24581;
    wire N__24580;
    wire N__24577;
    wire N__24570;
    wire N__24569;
    wire N__24562;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24504;
    wire N__24501;
    wire N__24500;
    wire N__24497;
    wire N__24492;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24474;
    wire N__24473;
    wire N__24470;
    wire N__24465;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24451;
    wire N__24450;
    wire N__24449;
    wire N__24446;
    wire N__24441;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24429;
    wire N__24428;
    wire N__24425;
    wire N__24424;
    wire N__24423;
    wire N__24422;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24401;
    wire N__24398;
    wire N__24393;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24377;
    wire N__24374;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24342;
    wire N__24341;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24319;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24301;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24278;
    wire N__24271;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24222;
    wire N__24221;
    wire N__24220;
    wire N__24219;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24201;
    wire N__24198;
    wire N__24193;
    wire N__24184;
    wire N__24183;
    wire N__24182;
    wire N__24181;
    wire N__24180;
    wire N__24179;
    wire N__24178;
    wire N__24177;
    wire N__24176;
    wire N__24175;
    wire N__24174;
    wire N__24173;
    wire N__24172;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24164;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24142;
    wire N__24141;
    wire N__24140;
    wire N__24139;
    wire N__24138;
    wire N__24137;
    wire N__24136;
    wire N__24135;
    wire N__24134;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24115;
    wire N__24114;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24102;
    wire N__24097;
    wire N__24096;
    wire N__24095;
    wire N__24094;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24082;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24056;
    wire N__24051;
    wire N__24044;
    wire N__24041;
    wire N__24034;
    wire N__24031;
    wire N__24026;
    wire N__24023;
    wire N__24018;
    wire N__24017;
    wire N__24016;
    wire N__24013;
    wire N__24012;
    wire N__24011;
    wire N__24010;
    wire N__24009;
    wire N__24008;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23994;
    wire N__23993;
    wire N__23986;
    wire N__23977;
    wire N__23968;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23946;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23886;
    wire N__23885;
    wire N__23882;
    wire N__23877;
    wire N__23872;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23835;
    wire N__23832;
    wire N__23829;
    wire N__23826;
    wire N__23823;
    wire N__23822;
    wire N__23819;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23797;
    wire N__23794;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23786;
    wire N__23781;
    wire N__23778;
    wire N__23773;
    wire N__23772;
    wire N__23771;
    wire N__23770;
    wire N__23769;
    wire N__23766;
    wire N__23757;
    wire N__23752;
    wire N__23751;
    wire N__23750;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23698;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23667;
    wire N__23666;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23658;
    wire N__23657;
    wire N__23654;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23628;
    wire N__23625;
    wire N__23614;
    wire N__23613;
    wire N__23612;
    wire N__23611;
    wire N__23610;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23602;
    wire N__23597;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23567;
    wire N__23554;
    wire N__23553;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23528;
    wire N__23525;
    wire N__23520;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23499;
    wire N__23498;
    wire N__23497;
    wire N__23494;
    wire N__23487;
    wire N__23482;
    wire N__23481;
    wire N__23480;
    wire N__23479;
    wire N__23470;
    wire N__23467;
    wire N__23466;
    wire N__23465;
    wire N__23462;
    wire N__23461;
    wire N__23456;
    wire N__23455;
    wire N__23454;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23437;
    wire N__23434;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23407;
    wire N__23404;
    wire N__23401;
    wire N__23400;
    wire N__23399;
    wire N__23398;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23390;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23353;
    wire N__23350;
    wire N__23347;
    wire N__23346;
    wire N__23345;
    wire N__23344;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23330;
    wire N__23327;
    wire N__23320;
    wire N__23317;
    wire N__23316;
    wire N__23313;
    wire N__23312;
    wire N__23311;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23285;
    wire N__23282;
    wire N__23275;
    wire N__23272;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23254;
    wire N__23251;
    wire N__23250;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23242;
    wire N__23239;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23223;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23203;
    wire N__23202;
    wire N__23201;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23172;
    wire N__23171;
    wire N__23170;
    wire N__23167;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23140;
    wire N__23133;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23112;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23088;
    wire N__23083;
    wire N__23082;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23074;
    wire N__23073;
    wire N__23068;
    wire N__23065;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22987;
    wire N__22986;
    wire N__22983;
    wire N__22980;
    wire N__22977;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22939;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22888;
    wire N__22887;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22867;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22842;
    wire N__22839;
    wire N__22838;
    wire N__22835;
    wire N__22830;
    wire N__22825;
    wire N__22824;
    wire N__22823;
    wire N__22820;
    wire N__22815;
    wire N__22810;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22795;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22765;
    wire N__22764;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22747;
    wire N__22746;
    wire N__22743;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22669;
    wire N__22666;
    wire N__22663;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22587;
    wire N__22586;
    wire N__22583;
    wire N__22578;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22563;
    wire N__22562;
    wire N__22559;
    wire N__22554;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22542;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22527;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22425;
    wire N__22424;
    wire N__22421;
    wire N__22416;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22404;
    wire N__22403;
    wire N__22402;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22354;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22313;
    wire N__22312;
    wire N__22309;
    wire N__22302;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22281;
    wire N__22280;
    wire N__22277;
    wire N__22272;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22233;
    wire N__22230;
    wire N__22229;
    wire N__22226;
    wire N__22225;
    wire N__22224;
    wire N__22221;
    wire N__22212;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22198;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22185;
    wire N__22182;
    wire N__22181;
    wire N__22180;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22165;
    wire N__22164;
    wire N__22161;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22136;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22102;
    wire N__22099;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22081;
    wire N__22080;
    wire N__22079;
    wire N__22078;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22029;
    wire N__22026;
    wire N__22025;
    wire N__22022;
    wire N__22017;
    wire N__22014;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21991;
    wire N__21988;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21952;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21918;
    wire N__21917;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21905;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21889;
    wire N__21886;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21540;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21489;
    wire N__21486;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21243;
    wire N__21242;
    wire N__21239;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21171;
    wire N__21168;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21153;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21135;
    wire N__21134;
    wire N__21133;
    wire N__21132;
    wire N__21129;
    wire N__21128;
    wire N__21127;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21116;
    wire N__21113;
    wire N__21112;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21104;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21084;
    wire N__21083;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20974;
    wire N__20971;
    wire N__20966;
    wire N__20961;
    wire N__20956;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20926;
    wire N__20923;
    wire N__20920;
    wire N__20915;
    wire N__20912;
    wire N__20905;
    wire N__20902;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20881;
    wire N__20878;
    wire N__20875;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20857;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20845;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20833;
    wire N__20832;
    wire N__20831;
    wire N__20830;
    wire N__20829;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20803;
    wire N__20802;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20757;
    wire N__20752;
    wire N__20749;
    wire N__20744;
    wire N__20741;
    wire N__20738;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20722;
    wire N__20715;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20654;
    wire N__20653;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20642;
    wire N__20641;
    wire N__20640;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20632;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20610;
    wire N__20609;
    wire N__20606;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20513;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20493;
    wire N__20490;
    wire N__20485;
    wire N__20482;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20461;
    wire N__20454;
    wire N__20451;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20421;
    wire N__20420;
    wire N__20413;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20370;
    wire N__20367;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20355;
    wire N__20350;
    wire N__20347;
    wire N__20346;
    wire N__20343;
    wire N__20342;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20311;
    wire N__20308;
    wire N__20307;
    wire N__20306;
    wire N__20305;
    wire N__20304;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20286;
    wire N__20281;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20140;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20132;
    wire N__20131;
    wire N__20130;
    wire N__20129;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20118;
    wire N__20117;
    wire N__20116;
    wire N__20115;
    wire N__20114;
    wire N__20113;
    wire N__20112;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20008;
    wire N__19997;
    wire N__19988;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19938;
    wire N__19937;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19929;
    wire N__19928;
    wire N__19925;
    wire N__19924;
    wire N__19923;
    wire N__19922;
    wire N__19919;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19887;
    wire N__19886;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19844;
    wire N__19843;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19757;
    wire N__19750;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19716;
    wire N__19715;
    wire N__19714;
    wire N__19713;
    wire N__19710;
    wire N__19709;
    wire N__19706;
    wire N__19705;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19694;
    wire N__19693;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19685;
    wire N__19684;
    wire N__19683;
    wire N__19682;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19581;
    wire N__19578;
    wire N__19571;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19547;
    wire N__19544;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19518;
    wire N__19517;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19509;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19501;
    wire N__19500;
    wire N__19499;
    wire N__19498;
    wire N__19497;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19486;
    wire N__19485;
    wire N__19482;
    wire N__19481;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19384;
    wire N__19377;
    wire N__19374;
    wire N__19363;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19345;
    wire N__19340;
    wire N__19335;
    wire N__19332;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19256;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19240;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19225;
    wire N__19224;
    wire N__19223;
    wire N__19222;
    wire N__19221;
    wire N__19220;
    wire N__19217;
    wire N__19216;
    wire N__19215;
    wire N__19212;
    wire N__19211;
    wire N__19210;
    wire N__19209;
    wire N__19206;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19178;
    wire N__19171;
    wire N__19164;
    wire N__19153;
    wire N__19152;
    wire N__19151;
    wire N__19150;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19138;
    wire N__19135;
    wire N__19126;
    wire N__19125;
    wire N__19124;
    wire N__19123;
    wire N__19122;
    wire N__19121;
    wire N__19120;
    wire N__19119;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19108;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19073;
    wire N__19072;
    wire N__19067;
    wire N__19064;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19042;
    wire N__19041;
    wire N__19038;
    wire N__19035;
    wire N__19034;
    wire N__19031;
    wire N__19030;
    wire N__19029;
    wire N__19028;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19008;
    wire N__18997;
    wire N__18996;
    wire N__18993;
    wire N__18990;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18943;
    wire N__18940;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18921;
    wire N__18918;
    wire N__18917;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18906;
    wire N__18905;
    wire N__18904;
    wire N__18903;
    wire N__18900;
    wire N__18899;
    wire N__18898;
    wire N__18897;
    wire N__18896;
    wire N__18895;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18854;
    wire N__18851;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18795;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18750;
    wire N__18743;
    wire N__18738;
    wire N__18735;
    wire N__18730;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18718;
    wire N__18715;
    wire N__18714;
    wire N__18713;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18621;
    wire N__18620;
    wire N__18619;
    wire N__18618;
    wire N__18615;
    wire N__18614;
    wire N__18611;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18603;
    wire N__18600;
    wire N__18595;
    wire N__18594;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18571;
    wire N__18568;
    wire N__18553;
    wire N__18550;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18538;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18508;
    wire N__18505;
    wire N__18502;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18447;
    wire N__18446;
    wire N__18439;
    wire N__18438;
    wire N__18437;
    wire N__18434;
    wire N__18429;
    wire N__18428;
    wire N__18423;
    wire N__18420;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18408;
    wire N__18405;
    wire N__18404;
    wire N__18399;
    wire N__18398;
    wire N__18395;
    wire N__18394;
    wire N__18391;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18355;
    wire N__18354;
    wire N__18353;
    wire N__18350;
    wire N__18349;
    wire N__18348;
    wire N__18343;
    wire N__18342;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18318;
    wire N__18315;
    wire N__18312;
    wire N__18307;
    wire N__18304;
    wire N__18303;
    wire N__18302;
    wire N__18301;
    wire N__18300;
    wire N__18295;
    wire N__18294;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18256;
    wire N__18253;
    wire N__18250;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18238;
    wire N__18235;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18187;
    wire N__18184;
    wire N__18181;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18109;
    wire N__18106;
    wire N__18105;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18097;
    wire N__18096;
    wire N__18093;
    wire N__18092;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18080;
    wire N__18075;
    wire N__18072;
    wire N__18061;
    wire N__18058;
    wire N__18057;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18019;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18007;
    wire N__18004;
    wire N__18001;
    wire N__17998;
    wire N__17995;
    wire N__17992;
    wire N__17989;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17953;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17941;
    wire N__17938;
    wire N__17937;
    wire N__17934;
    wire N__17931;
    wire N__17930;
    wire N__17929;
    wire N__17924;
    wire N__17921;
    wire N__17920;
    wire N__17917;
    wire N__17916;
    wire N__17915;
    wire N__17914;
    wire N__17909;
    wire N__17906;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17894;
    wire N__17889;
    wire N__17886;
    wire N__17875;
    wire N__17874;
    wire N__17871;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17860;
    wire N__17857;
    wire N__17856;
    wire N__17855;
    wire N__17854;
    wire N__17853;
    wire N__17848;
    wire N__17845;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17824;
    wire N__17821;
    wire N__17806;
    wire N__17805;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17788;
    wire N__17787;
    wire N__17786;
    wire N__17785;
    wire N__17784;
    wire N__17781;
    wire N__17778;
    wire N__17775;
    wire N__17774;
    wire N__17773;
    wire N__17770;
    wire N__17769;
    wire N__17766;
    wire N__17761;
    wire N__17758;
    wire N__17755;
    wire N__17752;
    wire N__17749;
    wire N__17744;
    wire N__17739;
    wire N__17728;
    wire N__17727;
    wire N__17724;
    wire N__17721;
    wire N__17716;
    wire N__17713;
    wire N__17712;
    wire N__17711;
    wire N__17710;
    wire N__17709;
    wire N__17708;
    wire N__17707;
    wire N__17706;
    wire N__17703;
    wire N__17702;
    wire N__17701;
    wire N__17694;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17675;
    wire N__17670;
    wire N__17659;
    wire N__17656;
    wire N__17655;
    wire N__17650;
    wire N__17649;
    wire N__17646;
    wire N__17643;
    wire N__17638;
    wire N__17635;
    wire N__17634;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17605;
    wire N__17604;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17530;
    wire N__17527;
    wire N__17524;
    wire N__17521;
    wire N__17518;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17508;
    wire N__17505;
    wire N__17502;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17442;
    wire N__17439;
    wire N__17436;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17419;
    wire N__17418;
    wire N__17417;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17409;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17392;
    wire N__17383;
    wire N__17380;
    wire N__17379;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17358;
    wire N__17355;
    wire N__17348;
    wire N__17347;
    wire N__17346;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17336;
    wire N__17329;
    wire N__17320;
    wire N__17319;
    wire N__17318;
    wire N__17317;
    wire N__17314;
    wire N__17307;
    wire N__17306;
    wire N__17305;
    wire N__17304;
    wire N__17299;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17284;
    wire N__17277;
    wire N__17274;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17217;
    wire N__17216;
    wire N__17213;
    wire N__17208;
    wire N__17207;
    wire N__17206;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17194;
    wire N__17193;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17178;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17010;
    wire N__17007;
    wire N__17004;
    wire N__17001;
    wire N__16998;
    wire N__16995;
    wire N__16992;
    wire N__16987;
    wire N__16984;
    wire N__16981;
    wire N__16978;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16959;
    wire N__16958;
    wire N__16957;
    wire N__16956;
    wire N__16955;
    wire N__16952;
    wire N__16947;
    wire N__16942;
    wire N__16939;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16879;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16840;
    wire N__16837;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16825;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16809;
    wire N__16806;
    wire N__16803;
    wire N__16798;
    wire N__16795;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16785;
    wire N__16782;
    wire N__16777;
    wire N__16774;
    wire N__16771;
    wire N__16768;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16752;
    wire N__16749;
    wire N__16746;
    wire N__16741;
    wire N__16738;
    wire N__16735;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16708;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16696;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16678;
    wire N__16675;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16662;
    wire N__16661;
    wire N__16660;
    wire N__16657;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16632;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16624;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16610;
    wire N__16609;
    wire N__16608;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16593;
    wire N__16590;
    wire N__16585;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16567;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16549;
    wire N__16546;
    wire N__16543;
    wire N__16540;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16366;
    wire N__16363;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16342;
    wire N__16339;
    wire N__16338;
    wire N__16333;
    wire N__16330;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16233;
    wire N__16230;
    wire N__16227;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16183;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16111;
    wire N__16108;
    wire N__16105;
    wire N__16102;
    wire N__16099;
    wire N__16098;
    wire N__16093;
    wire N__16090;
    wire N__16089;
    wire N__16086;
    wire N__16083;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16053;
    wire N__16050;
    wire N__16049;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16022;
    wire N__16019;
    wire N__16012;
    wire N__16009;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15999;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15987;
    wire N__15984;
    wire N__15981;
    wire N__15978;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15928;
    wire N__15925;
    wire N__15924;
    wire N__15921;
    wire N__15918;
    wire N__15915;
    wire N__15912;
    wire N__15909;
    wire N__15906;
    wire N__15903;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15883;
    wire N__15880;
    wire N__15877;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15867;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15853;
    wire N__15852;
    wire N__15851;
    wire N__15848;
    wire N__15847;
    wire N__15846;
    wire N__15845;
    wire N__15836;
    wire N__15835;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15817;
    wire N__15814;
    wire N__15811;
    wire N__15808;
    wire N__15805;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15795;
    wire N__15794;
    wire N__15791;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15781;
    wire N__15778;
    wire N__15775;
    wire N__15770;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15747;
    wire N__15746;
    wire N__15743;
    wire N__15738;
    wire N__15737;
    wire N__15734;
    wire N__15733;
    wire N__15732;
    wire N__15729;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15705;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15685;
    wire N__15682;
    wire N__15679;
    wire N__15678;
    wire N__15677;
    wire N__15676;
    wire N__15675;
    wire N__15674;
    wire N__15673;
    wire N__15672;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15657;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15621;
    wire N__15620;
    wire N__15619;
    wire N__15616;
    wire N__15615;
    wire N__15612;
    wire N__15609;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15599;
    wire N__15596;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15574;
    wire N__15573;
    wire N__15572;
    wire N__15571;
    wire N__15570;
    wire N__15565;
    wire N__15562;
    wire N__15557;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15528;
    wire N__15527;
    wire N__15524;
    wire N__15523;
    wire N__15520;
    wire N__15517;
    wire N__15514;
    wire N__15511;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15495;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15441;
    wire N__15440;
    wire N__15439;
    wire N__15436;
    wire N__15435;
    wire N__15432;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15414;
    wire N__15411;
    wire N__15408;
    wire N__15405;
    wire N__15394;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15376;
    wire N__15373;
    wire N__15370;
    wire N__15367;
    wire N__15364;
    wire N__15361;
    wire N__15358;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15343;
    wire N__15340;
    wire N__15337;
    wire N__15334;
    wire N__15331;
    wire N__15328;
    wire N__15325;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15277;
    wire N__15274;
    wire N__15271;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15244;
    wire N__15241;
    wire N__15238;
    wire N__15235;
    wire N__15232;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15213;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15181;
    wire N__15178;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15145;
    wire N__15142;
    wire N__15139;
    wire N__15136;
    wire N__15133;
    wire N__15130;
    wire N__15127;
    wire N__15124;
    wire N__15121;
    wire N__15118;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15055;
    wire N__15052;
    wire N__15049;
    wire N__15046;
    wire N__15043;
    wire N__15040;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15021;
    wire N__15018;
    wire N__15015;
    wire N__15010;
    wire N__15007;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14962;
    wire N__14961;
    wire N__14958;
    wire N__14955;
    wire N__14952;
    wire N__14947;
    wire N__14946;
    wire N__14945;
    wire N__14942;
    wire N__14937;
    wire N__14934;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14895;
    wire N__14894;
    wire N__14891;
    wire N__14886;
    wire N__14883;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14856;
    wire N__14855;
    wire N__14854;
    wire N__14851;
    wire N__14844;
    wire N__14839;
    wire N__14836;
    wire N__14833;
    wire N__14830;
    wire N__14827;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14812;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14752;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14737;
    wire N__14734;
    wire N__14731;
    wire N__14728;
    wire N__14725;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14602;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14490;
    wire N__14487;
    wire N__14484;
    wire N__14483;
    wire N__14482;
    wire N__14481;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14470;
    wire N__14467;
    wire N__14466;
    wire N__14463;
    wire N__14460;
    wire N__14459;
    wire N__14458;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14416;
    wire N__14413;
    wire N__14410;
    wire N__14409;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14386;
    wire N__14385;
    wire N__14380;
    wire N__14377;
    wire N__14370;
    wire N__14365;
    wire N__14364;
    wire N__14361;
    wire N__14358;
    wire N__14355;
    wire N__14352;
    wire N__14349;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14327;
    wire N__14324;
    wire N__14321;
    wire N__14314;
    wire N__14311;
    wire N__14306;
    wire N__14303;
    wire N__14298;
    wire N__14295;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14283;
    wire N__14282;
    wire N__14281;
    wire N__14280;
    wire N__14277;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14269;
    wire N__14268;
    wire N__14267;
    wire N__14266;
    wire N__14265;
    wire N__14264;
    wire N__14263;
    wire N__14262;
    wire N__14259;
    wire N__14258;
    wire N__14257;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14242;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14147;
    wire N__14140;
    wire N__14131;
    wire N__14128;
    wire N__14121;
    wire N__14118;
    wire N__14115;
    wire N__14112;
    wire N__14109;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14091;
    wire N__14086;
    wire N__14083;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire VCCG0;
    wire \this_vga_signals.N_1307_0 ;
    wire N_428;
    wire N_842;
    wire rgb_c_4;
    wire M_vcounter_q_esr_RNIQ82H7_9;
    wire M_this_oam_ram_read_data_13;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_13 ;
    wire rgb_c_2;
    wire rgb_c_5;
    wire \this_ppu.oam_cache.N_561_0 ;
    wire \this_ppu.oam_cache.mem_17 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_17 ;
    wire \this_ppu.M_oam_cache_read_data_i_16 ;
    wire bfn_7_19_0_;
    wire \this_ppu.M_oam_cache_read_data_i_17 ;
    wire M_this_ppu_spr_addr_4;
    wire \this_ppu.offset_y_cry_0 ;
    wire \this_ppu.offset_y_cry_1 ;
    wire M_this_ppu_spr_addr_5;
    wire \this_ppu.oam_cache.mem_16 ;
    wire \this_ppu.oam_cache.mem_18 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_18 ;
    wire port_clk_c;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire M_this_oam_ram_read_data_12;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_12 ;
    wire \this_ppu.oam_cache.N_579_0 ;
    wire M_this_oam_ram_read_data_26;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_26 ;
    wire N_84;
    wire rgb_c_0;
    wire M_this_oam_ram_read_data_15;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_15 ;
    wire \this_ppu.oam_cache.N_577_0 ;
    wire \this_ppu.oam_cache.N_567_0 ;
    wire M_this_oam_ram_read_data_8;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_8 ;
    wire M_this_oam_ram_read_data_9;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_9 ;
    wire M_this_oam_ram_read_data_10;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_10 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_16 ;
    wire \this_ppu.oam_cache.mem_4 ;
    wire \this_ppu.N_985_0 ;
    wire \this_ppu.N_671_0 ;
    wire \this_ppu.N_426_0_cascade_ ;
    wire \this_ppu.un1_M_oam_curr_q_1_c2_cascade_ ;
    wire \this_ppu.N_986_0 ;
    wire \this_ppu.un1_M_oam_curr_q_1_c4_cascade_ ;
    wire \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_cascade_ ;
    wire \this_ppu.N_841_0 ;
    wire \this_ppu.N_841_0_cascade_ ;
    wire \this_ppu.N_669_0 ;
    wire \this_ppu.m18_i_o2_1_cascade_ ;
    wire \this_ppu.N_426_0 ;
    wire M_this_vga_signals_address_2;
    wire \this_ppu.oam_cache.mem_2 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_21 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_22 ;
    wire M_this_oam_ram_read_data_3;
    wire M_this_oam_ram_read_data_6;
    wire M_this_oam_ram_read_data_25;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_25 ;
    wire M_this_warmup_qZ0Z_1;
    wire M_this_warmup_qZ0Z_0;
    wire bfn_9_22_0_;
    wire M_this_warmup_qZ0Z_2;
    wire un1_M_this_warmup_d_cry_1;
    wire M_this_warmup_qZ0Z_3;
    wire un1_M_this_warmup_d_cry_2;
    wire M_this_warmup_qZ0Z_4;
    wire un1_M_this_warmup_d_cry_3;
    wire M_this_warmup_qZ0Z_5;
    wire un1_M_this_warmup_d_cry_4;
    wire M_this_warmup_qZ0Z_6;
    wire un1_M_this_warmup_d_cry_5;
    wire M_this_warmup_qZ0Z_7;
    wire un1_M_this_warmup_d_cry_6;
    wire M_this_warmup_qZ0Z_8;
    wire un1_M_this_warmup_d_cry_7;
    wire un1_M_this_warmup_d_cry_8;
    wire M_this_warmup_qZ0Z_9;
    wire bfn_9_23_0_;
    wire M_this_warmup_qZ0Z_10;
    wire un1_M_this_warmup_d_cry_9;
    wire M_this_warmup_qZ0Z_11;
    wire un1_M_this_warmup_d_cry_10;
    wire M_this_warmup_qZ0Z_12;
    wire un1_M_this_warmup_d_cry_11;
    wire M_this_warmup_qZ0Z_13;
    wire un1_M_this_warmup_d_cry_12;
    wire M_this_warmup_qZ0Z_14;
    wire un1_M_this_warmup_d_cry_13;
    wire M_this_warmup_qZ0Z_15;
    wire un1_M_this_warmup_d_cry_14;
    wire M_this_warmup_qZ0Z_16;
    wire un1_M_this_warmup_d_cry_15;
    wire un1_M_this_warmup_d_cry_16;
    wire M_this_warmup_qZ0Z_17;
    wire bfn_9_24_0_;
    wire M_this_warmup_qZ0Z_18;
    wire un1_M_this_warmup_d_cry_17;
    wire M_this_warmup_qZ0Z_19;
    wire un1_M_this_warmup_d_cry_18;
    wire M_this_warmup_qZ0Z_20;
    wire un1_M_this_warmup_d_cry_19;
    wire M_this_warmup_qZ0Z_21;
    wire un1_M_this_warmup_d_cry_20;
    wire M_this_warmup_qZ0Z_22;
    wire un1_M_this_warmup_d_cry_21;
    wire M_this_warmup_qZ0Z_23;
    wire un1_M_this_warmup_d_cry_22;
    wire M_this_warmup_qZ0Z_24;
    wire un1_M_this_warmup_d_cry_23;
    wire un1_M_this_warmup_d_cry_24;
    wire M_this_warmup_qZ0Z_25;
    wire bfn_9_25_0_;
    wire M_this_warmup_qZ0Z_26;
    wire un1_M_this_warmup_d_cry_25;
    wire un1_M_this_warmup_d_cry_26;
    wire M_this_warmup_qZ0Z_27;
    wire M_this_oam_ram_write_data_18;
    wire M_this_oam_ram_write_data_23;
    wire M_this_oam_ram_write_data_20;
    wire M_this_oam_ram_write_data_19;
    wire M_this_oam_ram_write_data_17;
    wire rgb_c_1;
    wire M_this_oam_ram_read_data_0;
    wire \this_ppu.oam_cache.N_586_0 ;
    wire \this_ppu.oam_cache.mem_10 ;
    wire \this_ppu.N_844_0 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_10 ;
    wire bfn_10_17_0_;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_0 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_1 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_2 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_3 ;
    wire \this_ppu.oam_cache.mem_7 ;
    wire N_41_0;
    wire M_this_ppu_oam_addr_1;
    wire \this_ppu.M_oam_cache_cnt_qZ0Z_4 ;
    wire \this_ppu.m62_0_a2_0_o2_0_cascade_ ;
    wire \this_ppu.un1_M_oam_curr_q_1_c4 ;
    wire \this_ppu.M_oam_curr_qc_0_1 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO ;
    wire \this_ppu.M_oam_cache_cnt_qZ0Z_1 ;
    wire \this_ppu.m62_0_a2_0_o2_1 ;
    wire M_this_ppu_oam_addr_3;
    wire M_this_ppu_oam_addr_2;
    wire M_this_ppu_oam_addr_4;
    wire \this_ppu.un1_M_oam_curr_q_1_c2 ;
    wire \this_ppu.un1_M_oam_curr_q_1_c5 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO ;
    wire \this_ppu.M_oam_cache_cnt_qZ0Z_3 ;
    wire M_this_oam_ram_read_data_24;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_24 ;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire M_this_oam_ram_read_data_7;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axb1_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_c3_cascade_ ;
    wire \this_vga_signals.haddress_1_0 ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_0_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_cascade_ ;
    wire \this_vga_signals.if_m2 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3 ;
    wire M_this_vga_signals_address_1;
    wire \this_vga_signals.mult1_un75_sum_axb1 ;
    wire \this_ppu.M_oam_cache_cnt_qZ1Z_0 ;
    wire M_this_vga_signals_address_3;
    wire M_this_oam_ram_read_data_16;
    wire \this_ppu.M_this_oam_ram_read_data_i_16 ;
    wire bfn_10_22_0_;
    wire \this_ppu.M_this_oam_ram_read_data_i_17 ;
    wire \this_ppu.un1_oam_data_1_cry_0 ;
    wire \this_ppu.M_this_oam_ram_read_data_i_18 ;
    wire \this_ppu.un1_oam_data_1_cry_1 ;
    wire \this_ppu.un1_oam_data_1_cry_2 ;
    wire \this_ppu.un1_oam_data_1_cry_3 ;
    wire \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0 ;
    wire \this_ppu.un1_oam_data_1_cry_4 ;
    wire \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0 ;
    wire \this_ppu.un1_oam_data_1_cry_5 ;
    wire \this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0 ;
    wire \this_ppu.un1_oam_data_1_cry_2_c_RNIR4HDZ0 ;
    wire \this_ppu.un1_oam_data_1_cry_6 ;
    wire \this_ppu.m28_e_i_o3_2 ;
    wire M_this_oam_ram_read_data_18;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_18 ;
    wire M_this_oam_ram_write_data_5;
    wire M_this_oam_ram_read_data_22;
    wire M_this_oam_ram_read_data_i_22;
    wire M_this_oam_ram_read_data_29;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_29 ;
    wire M_this_oam_ram_read_data_21;
    wire M_this_oam_ram_read_data_i_21;
    wire M_this_oam_ram_read_data_31;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_31 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_19 ;
    wire M_this_oam_ram_read_data_19;
    wire M_this_oam_ram_read_data_i_19;
    wire M_this_oam_ram_write_data_10;
    wire N_260;
    wire M_this_oam_ram_read_data_28;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_28 ;
    wire M_this_oam_ram_write_data_9;
    wire M_this_oam_ram_read_data_i_20;
    wire M_this_oam_ram_write_data_28;
    wire M_this_oam_ram_write_data_8;
    wire M_this_oam_ram_write_data_31;
    wire M_this_oam_ram_write_data_16;
    wire M_this_oam_ram_write_data_24;
    wire \this_vga_signals.hsync_1_i_0_0_1 ;
    wire M_this_oam_ram_read_data_14;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_14 ;
    wire \this_vga_signals.hsync_1_i_0_0_a3_0_0 ;
    wire \this_vga_signals.N_811_0 ;
    wire rgb_c_3;
    wire M_this_ppu_oam_addr_5;
    wire M_this_ppu_oam_addr_0;
    wire \this_ppu.m35_i_0_a3_1_3 ;
    wire \this_ppu.N_1394 ;
    wire M_this_oam_ram_read_data_2;
    wire \this_ppu.m28_e_i_a3_4 ;
    wire \this_ppu.m28_e_i_a3_3 ;
    wire \this_ppu.N_1184_7_cascade_ ;
    wire \this_ppu.m18_i_1 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0_2 ;
    wire \this_ppu.oam_cache.mem_12 ;
    wire M_this_oam_ram_read_data_5;
    wire \this_ppu.oam_cache.N_569_0 ;
    wire M_this_oam_ram_read_data_4;
    wire \this_ppu.oam_cache.N_575_0 ;
    wire \this_ppu.N_1182 ;
    wire \this_vga_signals.if_N_9_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_c3 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_2_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_1 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0 ;
    wire \this_vga_signals.mult1_un75_sum_c2_0 ;
    wire \this_vga_signals.mult1_un75_sum_c2_0_cascade_ ;
    wire \this_vga_signals.if_N_8_i ;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire M_this_oam_ram_read_data_27;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_27 ;
    wire \this_ppu.oam_cache.mem_0 ;
    wire \this_ppu.un1_oam_data_1_axb_7 ;
    wire M_this_oam_ram_write_data_6;
    wire M_this_data_tmp_qZ0Z_6;
    wire M_this_oam_ram_write_data_7;
    wire M_this_data_tmp_qZ0Z_7;
    wire M_this_oam_ram_read_data_17;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_17 ;
    wire M_this_data_tmp_qZ0Z_10;
    wire M_this_data_tmp_qZ0Z_8;
    wire M_this_data_tmp_qZ0Z_9;
    wire M_this_oam_ram_write_data_26;
    wire M_this_oam_ram_write_data_27;
    wire M_this_oam_ram_write_data_30;
    wire M_this_data_tmp_qZ0Z_15;
    wire M_this_oam_ram_write_data_15;
    wire M_this_data_tmp_qZ0Z_16;
    wire M_this_data_tmp_qZ0Z_17;
    wire M_this_data_tmp_qZ0Z_19;
    wire M_this_data_tmp_qZ0Z_20;
    wire M_this_data_tmp_qZ0Z_18;
    wire M_this_oam_ram_write_data_0;
    wire \this_vga_ramdac.N_852_i_reto ;
    wire \this_vga_signals.N_298_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_d7_0_i_0_o3_0_o3_4_a2_0 ;
    wire \this_vga_signals.N_1044_0_cascade_ ;
    wire \this_vga_signals.N_298_0 ;
    wire \this_vga_signals.hsync_1_i_0_0_a3_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire bfn_12_17_0_;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_12_18_0_;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz ;
    wire \this_ppu.N_1184_7 ;
    wire \this_ppu.un1_M_state_q_7_i_0 ;
    wire M_this_oam_ram_read_data_11;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_11 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_12 ;
    wire \this_ppu.oam_cache.mem_15 ;
    wire \this_vga_signals.mult1_un54_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.N_968 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.N_968_cascade_ ;
    wire \this_vga_signals.N_291_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb1 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_2 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb2 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_0 ;
    wire M_this_oam_ram_read_data_20;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_20 ;
    wire \this_ppu.oam_cache.mem_13 ;
    wire M_this_vga_signals_address_4;
    wire N_852_0;
    wire \this_vga_signals.mult1_un54_sum_c3 ;
    wire M_this_vga_signals_address_5;
    wire M_this_oam_ram_write_data_3;
    wire M_this_data_tmp_qZ0Z_3;
    wire M_this_oam_ram_write_data_4;
    wire M_this_data_tmp_qZ0Z_4;
    wire M_this_data_tmp_qZ0Z_5;
    wire M_this_oam_ram_write_data_29;
    wire M_this_oam_ram_write_data_21;
    wire M_this_oam_ram_write_data_1;
    wire M_this_oam_ram_write_data_25;
    wire M_this_data_tmp_qZ0Z_21;
    wire M_this_data_tmp_qZ0Z_23;
    wire M_this_data_tmp_qZ0Z_0;
    wire \this_vga_ramdac.N_3856_reto ;
    wire \this_vga_ramdac.i2_mux_cascade_ ;
    wire \this_vga_ramdac.N_3858_reto ;
    wire \this_vga_ramdac.N_24_mux ;
    wire M_this_vram_read_data_0;
    wire M_this_vram_read_data_2;
    wire M_this_vram_read_data_3;
    wire M_this_vram_read_data_1;
    wire \this_vga_ramdac.m6_cascade_ ;
    wire \this_vga_ramdac.N_3857_reto ;
    wire \this_ppu.oam_cache.mem_9 ;
    wire \this_vga_signals.M_pcounter_q_ret_RNIB85CZ0Z3_cascade_ ;
    wire \this_vga_signals.N_3_0_cascade_ ;
    wire \this_vga_ramdac.m16 ;
    wire M_pcounter_q_ret_1_RNIOILK7_cascade_;
    wire \this_vga_ramdac.N_3859_reto ;
    wire \this_vga_signals.N_2_0 ;
    wire \this_vga_signals.N_2_0_cascade_ ;
    wire \this_vga_ramdac.m19 ;
    wire \this_vga_ramdac.N_3860_reto ;
    wire \this_ppu.oam_cache.mem_14 ;
    wire \this_ppu.m35_i_0_a3_0_cascade_ ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_9 ;
    wire \this_ppu.oam_cache.mem_11 ;
    wire \this_ppu.oam_cache.mem_1 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_14 ;
    wire \this_ppu.N_1196_1 ;
    wire \this_ppu.M_oam_curr_qZ0Z_6 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_13 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9_cascade_ ;
    wire \this_vga_signals.N_1307_1 ;
    wire \this_ppu.oam_cache.mem_8 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_11 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc1_0 ;
    wire this_pixel_clk_M_counter_q_0;
    wire this_pixel_clk_M_counter_q_i_1;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_2 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_3 ;
    wire \this_vga_signals.M_hcounter_q_RNII1437Z0Z_3 ;
    wire M_this_oam_ram_read_data_30;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_30 ;
    wire \this_ppu.oam_cache.mem_3 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_1 ;
    wire read_data_RNI5QFJ1_1;
    wire \this_ppu.M_oam_cache_read_data_16 ;
    wire M_this_ppu_spr_addr_3;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_2 ;
    wire read_data_RNI6RFJ1_2;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_3 ;
    wire read_data_RNI7SFJ1_3;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_4 ;
    wire read_data_RNI9TFJ1_4;
    wire \this_vga_signals.M_pcounter_q_0Z0Z_1 ;
    wire M_this_data_tmp_qZ0Z_11;
    wire M_this_oam_ram_write_data_11;
    wire M_this_oam_ram_write_data_12;
    wire M_this_oam_ram_write_data_13;
    wire M_this_oam_ram_write_data_14;
    wire M_this_data_tmp_qZ0Z_12;
    wire M_this_data_tmp_qZ0Z_14;
    wire M_this_data_tmp_qZ0Z_1;
    wire M_this_oam_ram_write_data_22;
    wire M_this_data_tmp_qZ0Z_22;
    wire M_this_map_ram_read_data_1;
    wire N_724_0;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire \this_vga_signals.N_1417 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_0 ;
    wire \this_vga_ramdac.i2_mux_0 ;
    wire M_pcounter_q_ret_1_RNIOILK7;
    wire \this_vga_ramdac.N_3861_reto ;
    wire \this_ppu.un1_M_surface_x_q_ac0_11 ;
    wire M_this_ppu_spr_addr_0;
    wire \this_ppu.M_oam_cache_read_data_8 ;
    wire \this_ppu.M_oam_cache_read_data_i_8 ;
    wire bfn_14_19_0_;
    wire \this_ppu.M_oam_cache_read_data_i_9 ;
    wire M_this_ppu_spr_addr_1;
    wire \this_ppu.offset_x_cry_0 ;
    wire \this_ppu.M_oam_cache_read_data_i_10 ;
    wire M_this_ppu_spr_addr_2;
    wire \this_ppu.offset_x_cry_1 ;
    wire \this_ppu.M_oam_cache_read_data_i_11 ;
    wire \this_ppu.m68_0_o2_0 ;
    wire \this_ppu.offset_x_cry_2 ;
    wire \this_ppu.M_oam_cache_read_data_i_12 ;
    wire \this_ppu.offset_x_4 ;
    wire \this_ppu.offset_x_cry_3 ;
    wire \this_ppu.M_oam_cache_read_data_i_13 ;
    wire \this_ppu.offset_x_5 ;
    wire \this_ppu.offset_x_cry_4 ;
    wire \this_ppu.M_oam_cache_read_data_i_14 ;
    wire M_this_ppu_map_addr_3;
    wire \this_ppu.offset_x_6 ;
    wire \this_ppu.offset_x_cry_5 ;
    wire GNDG0;
    wire \this_ppu.offset_x_cry_6 ;
    wire \this_ppu.offset_x_cry_6_THRU_CRY_0_THRU_CO ;
    wire \this_ppu.M_oam_cache_read_data_15 ;
    wire M_this_ppu_map_addr_4;
    wire bfn_14_20_0_;
    wire \this_ppu.offset_x_7 ;
    wire \this_ppu.m13_0_i_1 ;
    wire bfn_14_21_0_;
    wire \this_ppu.offset_y ;
    wire \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO ;
    wire \this_ppu.M_screen_y_q_esr_RNI453Q6Z0Z_1 ;
    wire \this_ppu.M_surface_y_qZ0Z_1 ;
    wire \this_ppu.un1_M_surface_y_d_cry_0 ;
    wire \this_ppu.M_surface_y_qZ0Z_2 ;
    wire \this_ppu.un1_M_surface_y_d_cry_1 ;
    wire M_this_ppu_map_addr_5;
    wire \this_ppu.un1_M_surface_y_d_cry_2 ;
    wire \this_ppu.M_screen_y_q_RNI8FJF7Z0Z_4 ;
    wire M_this_ppu_map_addr_6;
    wire \this_ppu.un1_M_surface_y_d_cry_3 ;
    wire M_this_ppu_map_addr_7;
    wire \this_ppu.un1_M_surface_y_d_cry_4 ;
    wire M_this_ppu_map_addr_8;
    wire \this_ppu.un1_M_surface_y_d_cry_5 ;
    wire \this_ppu.un1_M_surface_y_d_cry_6 ;
    wire bfn_14_22_0_;
    wire M_this_ppu_map_addr_9;
    wire \this_ppu.M_screen_y_q_esr_RNI563Q6Z0Z_2 ;
    wire M_this_oam_ram_read_data_23;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_23 ;
    wire M_this_oam_ram_read_data_1;
    wire \this_ppu.oam_cache.N_581_0 ;
    wire M_this_data_tmp_qZ0Z_13;
    wire bfn_14_24_0_;
    wire M_this_data_count_q_cry_0;
    wire M_this_data_count_q_cry_1;
    wire M_this_data_count_q_cry_2;
    wire M_this_data_count_q_cry_3;
    wire M_this_data_count_q_cry_4;
    wire M_this_data_count_q_cry_5;
    wire M_this_data_count_q_cry_6;
    wire M_this_data_count_q_cry_7;
    wire bfn_14_25_0_;
    wire M_this_data_count_q_cry_8;
    wire M_this_data_count_q_cry_9;
    wire M_this_data_count_q_cry_10;
    wire M_this_data_count_q_cry_11;
    wire M_this_data_count_q_cry_12;
    wire M_this_oam_address_qZ0Z_7;
    wire IO_port_data_write_i_m2_i_m2_0;
    wire GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO;
    wire \this_ppu.M_state_qZ0Z_8 ;
    wire \this_ppu.N_762_0 ;
    wire \this_ppu.N_91_0 ;
    wire \this_ppu.N_91_0_cascade_ ;
    wire \this_ppu.un1_M_surface_x_q_c3 ;
    wire \this_ppu.un1_M_surface_x_q_c3_cascade_ ;
    wire \this_ppu.un1_M_surface_x_q_c6 ;
    wire \this_ppu.N_1202 ;
    wire \this_ppu.M_state_qZ0Z_1 ;
    wire M_this_status_flags_qZ0Z_0;
    wire \this_ppu.N_1201 ;
    wire \this_ppu.M_state_qZ0Z_4 ;
    wire \this_ppu.M_state_q_srsts_1_8 ;
    wire \this_ppu.N_1145 ;
    wire \this_ppu.M_screen_y_qZ0Z_7 ;
    wire \this_ppu.M_screen_y_qZ0Z_1 ;
    wire \this_ppu.un3_M_screen_y_d_0_c2 ;
    wire \this_ppu.un3_M_screen_y_d_0_c2_cascade_ ;
    wire \this_ppu.un3_M_screen_y_d_0_c4_cascade_ ;
    wire \this_ppu.un3_M_screen_y_d_0_c6 ;
    wire N_861_0_cascade_;
    wire \this_ppu.M_screen_y_qZ0Z_2 ;
    wire \this_ppu.un3_M_screen_y_d_a_2 ;
    wire M_this_ppu_vram_addr_7;
    wire \this_ppu.M_screen_y_q_RNIQ9FQ6Z0Z_0 ;
    wire \this_ppu.un1_M_screen_x_q_c4_cascade_ ;
    wire \this_ppu.un1_M_screen_x_q_c4 ;
    wire M_this_ppu_vram_addr_4;
    wire \this_ppu.un1_M_screen_x_q_c5_cascade_ ;
    wire M_this_ppu_vram_addr_5;
    wire M_this_ppu_vram_addr_6;
    wire M_this_ppu_vram_addr_2;
    wire M_this_scroll_qZ0Z_0;
    wire M_this_scroll_qZ0Z_1;
    wire M_this_scroll_qZ0Z_2;
    wire M_this_scroll_qZ0Z_4;
    wire M_this_scroll_qZ0Z_7;
    wire this_vga_signals_vsync_1_i;
    wire M_this_data_count_qZ0Z_0;
    wire M_this_data_count_q_cry_0_THRU_CO;
    wire M_this_data_count_qZ0Z_1;
    wire M_this_data_count_q_cry_1_THRU_CO;
    wire M_this_data_count_qZ0Z_2;
    wire M_this_data_count_q_cry_2_THRU_CO;
    wire M_this_data_count_qZ0Z_3;
    wire M_this_data_count_q_cry_3_THRU_CO;
    wire M_this_data_count_q_cry_4_THRU_CO;
    wire M_this_data_count_q_cry_5_THRU_CO;
    wire M_this_data_count_q_cry_10_THRU_CO;
    wire M_this_data_count_q_s_10;
    wire M_this_data_count_q_cry_11_THRU_CO;
    wire M_this_data_count_q_s_13;
    wire M_this_data_count_qZ0Z_12;
    wire M_this_data_count_qZ0Z_11;
    wire M_this_data_count_qZ0Z_13;
    wire M_this_data_count_qZ0Z_10;
    wire M_this_data_count_q_s_8;
    wire M_this_data_count_qZ0Z_8;
    wire M_this_data_count_qZ0Z_5;
    wire M_this_data_count_qZ0Z_4;
    wire un1_M_this_oam_address_q_c6;
    wire \this_vga_signals.g0_1 ;
    wire \this_vga_signals.N_3_0 ;
    wire \this_vga_signals.M_pcounter_q_i_2_1 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO ;
    wire \this_ppu.M_oam_cache_cnt_qZ0Z_2 ;
    wire \this_vga_signals.M_lcounter_q_e_1_0_cascade_ ;
    wire N_26;
    wire \this_ppu.N_1198 ;
    wire \this_ppu.N_1198_cascade_ ;
    wire M_this_ppu_map_addr_1;
    wire \this_ppu.un1_M_surface_x_q_c2_cascade_ ;
    wire \this_ppu.un1_M_surface_x_q_c5_cascade_ ;
    wire M_this_ppu_map_addr_2;
    wire \this_ppu.un1_M_surface_x_q_c2 ;
    wire \this_ppu.offset_x ;
    wire \this_ppu.un1_M_surface_x_q_c1 ;
    wire M_this_ppu_map_addr_0;
    wire \this_ppu.M_surface_x_qZ0Z_2 ;
    wire \this_ppu.un1_M_surface_x_q_c1_cascade_ ;
    wire \this_ppu.M_surface_x_qZ0Z_1 ;
    wire \this_ppu.un1_M_surface_x_q_c4 ;
    wire \this_ppu.M_state_qZ0Z_2 ;
    wire \this_ppu.M_state_qZ0Z_10 ;
    wire M_this_ppu_vram_addr_3;
    wire \this_ppu.N_798_0_cascade_ ;
    wire M_this_ppu_vram_data_0;
    wire \this_ppu.N_1182_1 ;
    wire \this_ppu.M_state_qZ0Z_5 ;
    wire \this_vga_signals.g0_2 ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_cascade_ ;
    wire M_this_vga_signals_address_7;
    wire \this_ppu.M_state_qZ0Z_6 ;
    wire \this_ppu.N_82_0 ;
    wire \this_ppu.N_1659_0 ;
    wire \this_ppu.M_screen_y_qZ0Z_3 ;
    wire M_this_scroll_qZ0Z_3;
    wire \this_ppu.M_screen_y_q_esr_RNIF77F7Z0Z_3 ;
    wire \this_ppu.M_state_qZ0Z_9 ;
    wire \this_ppu.M_state_qZ0Z_7 ;
    wire \this_ppu.N_61_0 ;
    wire M_this_ppu_vram_addr_1;
    wire \this_ppu.N_61_0_cascade_ ;
    wire M_this_ppu_vram_addr_0;
    wire \this_ppu.un1_M_screen_x_q_c2 ;
    wire \this_ppu.M_state_d30_i_i_o2_3 ;
    wire \this_ppu.N_79_0 ;
    wire \this_ppu.N_79_0_cascade_ ;
    wire \this_ppu.M_pixel_cnt_q_600_1 ;
    wire \this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_i_0_0 ;
    wire \this_ppu.N_999_0 ;
    wire \this_ppu.N_838_0 ;
    wire \this_ppu.M_state_qZ0Z_0 ;
    wire \this_ppu.N_1042_0 ;
    wire \this_ppu.M_state_qZ0Z_11 ;
    wire \this_ppu.M_state_qZ0Z_3 ;
    wire \this_ppu.N_1042_0_cascade_ ;
    wire \this_ppu.un30_0_a2_i_0 ;
    wire \this_ppu.M_pixel_cnt_qZ0Z_0 ;
    wire bfn_16_23_0_;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1 ;
    wire \this_ppu.M_pixel_cnt_qZ0Z_3 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_CO ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1 ;
    wire CONSTANT_ONE_NET;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1 ;
    wire \this_ppu.M_pixel_cnt_qZ0Z_7 ;
    wire \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_6_s1 ;
    wire \this_ppu.N_1205 ;
    wire \this_ppu.M_state_d30_i_i_o2_4 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_CO ;
    wire \this_ppu.M_pixel_cnt_qZ0Z_1 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_CO ;
    wire \this_ppu.M_pixel_cnt_qZ0Z_2 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_CO ;
    wire \this_ppu.M_pixel_cnt_qZ0Z_5 ;
    wire \this_ppu.N_1301_cascade_ ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_CO ;
    wire \this_ppu.M_pixel_cnt_qZ0Z_6 ;
    wire \this_ppu.N_1730_0 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_CO ;
    wire \this_ppu.N_677_0 ;
    wire \this_ppu.M_pixel_cnt_qZ0Z_4 ;
    wire M_this_data_count_q_cry_6_THRU_CO;
    wire M_this_data_count_q_cry_8_THRU_CO;
    wire M_this_data_count_qZ0Z_9;
    wire N_231;
    wire M_this_data_tmp_qZ0Z_2;
    wire M_this_oam_ram_write_data_2;
    wire M_this_data_count_qZ0Z_7;
    wire M_this_data_count_qZ0Z_6;
    wire \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_16 ;
    wire N_1709_0;
    wire N_1693_0;
    wire \this_vga_signals.M_vcounter_q_esr_RNI01JU6Z0Z_9 ;
    wire \this_ppu.N_1269_cascade_ ;
    wire \this_ppu.N_1006_0 ;
    wire \this_vga_signals.N_1264_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x0 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x1 ;
    wire M_this_scroll_qZ0Z_10;
    wire M_this_scroll_qZ0Z_11;
    wire M_this_scroll_qZ0Z_12;
    wire M_this_scroll_qZ0Z_13;
    wire M_this_scroll_qZ0Z_14;
    wire M_this_scroll_qZ0Z_15;
    wire M_this_scroll_qZ0Z_8;
    wire M_this_scroll_qZ0Z_9;
    wire \this_vga_signals.mult1_un61_sum_c3_0_2_cascade_ ;
    wire \this_vga_signals.N_4_0 ;
    wire \this_vga_signals.if_m1_0_x2_1 ;
    wire \this_vga_signals.r_N_2_i_0 ;
    wire \this_vga_signals.N_836_0 ;
    wire \this_vga_signals.N_1043_cascade_ ;
    wire this_vga_signals_M_lcounter_q_0;
    wire N_792_0;
    wire this_vga_signals_M_lcounter_q_1;
    wire \this_ppu.M_last_q_0 ;
    wire N_771_0;
    wire N_771_0_cascade_;
    wire \this_ppu.N_774_0 ;
    wire \this_vga_signals.g1_0_0_cascade_ ;
    wire \this_vga_signals.if_N_6_0_0_0 ;
    wire \this_vga_signals.g1_0_0 ;
    wire \this_vga_signals.N_27_0_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_1_0_cascade_ ;
    wire M_this_reset_cond_out_0;
    wire N_782_0;
    wire N_1725_0;
    wire N_1717_0;
    wire \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_12 ;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_16 ;
    wire \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_16 ;
    wire \this_ppu.M_this_state_q_srsts_i_a2_10Z0Z_16 ;
    wire N_778_0_cascade_;
    wire N_1701_0;
    wire un1_M_this_oam_address_q_c5;
    wire M_this_oam_address_qZ0Z_5;
    wire un1_M_this_oam_address_q_c5_cascade_;
    wire M_this_oam_address_qZ0Z_6;
    wire un1_M_this_oam_address_q_c2;
    wire M_this_oam_address_qZ0Z_2;
    wire M_this_oam_address_qZ0Z_3;
    wire un1_M_this_oam_address_q_c3;
    wire M_this_oam_address_qZ0Z_4;
    wire M_this_oam_address_qZ0Z_1;
    wire M_this_oam_address_qZ0Z_0;
    wire N_778_0;
    wire M_this_oam_ram_write_data_0_sqmuxa;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb2_i ;
    wire \this_vga_signals.mult1_un54_sum_2_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0 ;
    wire \this_ppu.N_1115 ;
    wire \this_vga_signals.g0_33_N_3L4 ;
    wire \this_vga_signals.g0_33_N_4L6 ;
    wire \this_vga_signals.g0_33_N_5L8 ;
    wire \this_vga_signals.M_hcounter_d7_0_i_0_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire bfn_18_21_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire G_535;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire bfn_18_22_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.g0_0_0 ;
    wire \this_vga_signals.IO_port_data_write_0_a2_i_o2_2Z0Z_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.vsync_1_0_a3_0_a3_5 ;
    wire M_this_state_qZ0Z_12;
    wire \this_ppu.N_430_1_0_cascade_ ;
    wire M_this_state_q_fastZ0Z_13;
    wire \this_vga_signals.N_38_i_0_a2_3Z0Z_0_cascade_ ;
    wire \this_vga_signals.N_38_i_0_a2_3_xZ0Z1_cascade_ ;
    wire \this_vga_signals.N_38_i_0_a2_3_cascade_ ;
    wire \this_vga_signals.N_38_i_0_a2_0_3 ;
    wire port_enb_c;
    wire this_start_data_delay_M_last_q;
    wire M_this_delay_clk_out_0;
    wire N_765_0_cascade_;
    wire \this_ppu.N_229_1_0 ;
    wire \this_ppu.N_229_1_0_cascade_ ;
    wire N_229;
    wire N_1423;
    wire \this_vga_signals.SUM_2_i_i_1_0_3_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_x0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_x1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_0_ns_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_1_0 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_1_1 ;
    wire \this_vga_signals.if_m5_s_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_cascade_ ;
    wire \this_vga_signals.if_m5_d ;
    wire \this_vga_signals.if_m5_d_cascade_ ;
    wire \this_vga_signals.N_2840_0_0 ;
    wire \this_vga_signals.N_27_0_0 ;
    wire \this_vga_signals.vaddress_7_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c2_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3 ;
    wire \this_vga_signals.g1_2_0_cascade_ ;
    wire \this_vga_signals.if_m6_i_x2_3 ;
    wire \this_vga_signals.g1_3 ;
    wire this_vga_signals_CO0_0_i_i;
    wire this_vga_signals_CO0_0_i_i_cascade_;
    wire \this_vga_signals.vaddress_8 ;
    wire \this_vga_signals.g1 ;
    wire \this_vga_signals.N_39_0 ;
    wire \this_vga_signals.vaddress_7 ;
    wire \this_vga_signals.N_38_i_0_a2_0_4Z0Z_1 ;
    wire \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_17_cascade_ ;
    wire M_this_state_qZ0Z_17;
    wire \this_vga_signals.vsync_1_0_a3_0_a3_0 ;
    wire M_this_state_qZ0Z_18;
    wire this_ppu_M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0;
    wire \this_ppu.N_1322_cascade_ ;
    wire M_this_spr_ram_write_data_0;
    wire \this_vga_signals.N_1247 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0_cascade_ ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_9 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_1_1_1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.M_vcounter_q_5_repZ0Z1 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c2_0_cascade_ ;
    wire \this_vga_signals.g0_4 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_4_3 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_x1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_3 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1 ;
    wire \this_vga_signals.N_27_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_x0 ;
    wire \this_vga_signals.if_N_7_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_d_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_1_3 ;
    wire \this_vga_signals.mult1_un54_sum_1_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c ;
    wire \this_vga_signals.mult1_un54_sum_0_3_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_d ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0 ;
    wire \this_vga_signals.N_3_1_0_1 ;
    wire \this_vga_signals.g0_2_1 ;
    wire \this_vga_signals.g0_5 ;
    wire \this_vga_signals.mult1_un61_sum_axb1_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire \this_vga_signals.g0_1_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0 ;
    wire \this_vga_signals.mult1_un68_sum_c2_0_cascade_ ;
    wire \this_vga_signals.g0_0_3_1 ;
    wire \this_vga_signals.g0_0_3 ;
    wire \this_vga_signals.g1_1 ;
    wire \this_vga_signals.mult1_un54_sum_0_1 ;
    wire \this_vga_signals.g0_2_0 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_0 ;
    wire \this_vga_signals.vaddress_9 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_1 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_i ;
    wire \this_vga_signals.g0_0_x2 ;
    wire \this_vga_signals.if_m5_i_0_0_0 ;
    wire \this_ppu.N_1002_0 ;
    wire \this_ppu.N_235_2_0 ;
    wire \this_ppu.N_235_2_0_cascade_ ;
    wire M_this_state_qZ0Z_7;
    wire \this_ppu.N_1162 ;
    wire M_this_state_qZ0Z_9;
    wire M_this_state_qZ0Z_11;
    wire \this_ppu.N_1301 ;
    wire \this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_15 ;
    wire M_this_state_qZ0Z_15;
    wire \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_7 ;
    wire \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_11 ;
    wire \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_8 ;
    wire \this_ppu.N_807_0_cascade_ ;
    wire \this_ppu.N_1341 ;
    wire M_this_spr_ram_write_data_2;
    wire \this_ppu.oam_cache.mem_5 ;
    wire \this_vga_signals.mult1_un54_sum_1_3 ;
    wire \this_vga_signals.mult1_un47_sum_0_3_cascade_ ;
    wire \this_vga_signals.N_7 ;
    wire \this_vga_signals.mult1_un47_sum_2_3 ;
    wire \this_vga_signals.mult1_un47_sum_3_3_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_2_0_3 ;
    wire \this_ppu.m18_i_o2_0 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_0_3_0_0 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0 ;
    wire N_814_0_cascade_;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_2_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_2_2_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_c3_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_2_2 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_0_2_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_x1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_x0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_1 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0 ;
    wire \this_vga_signals.mult1_un47_sum_c2_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3 ;
    wire \this_vga_signals.g1_0 ;
    wire \this_vga_signals.g0_0_1 ;
    wire \this_vga_signals.g0_3_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un54_sum_c2_0 ;
    wire \this_vga_signals.M_vcounter_q_9_repZ0Z1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0 ;
    wire \this_vga_signals.M_vcounter_q_8_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_7_repZ0Z1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_3_cascade_ ;
    wire \this_vga_signals.g1_0_0_0_cascade_ ;
    wire \this_vga_signals.SUM_2_i_i_1_0_3 ;
    wire \this_vga_signals.N_5_0_0 ;
    wire \this_vga_signals.g1_0_1 ;
    wire \this_vga_signals.N_39_0_0 ;
    wire \this_vga_signals.g1_3_0_0_cascade_ ;
    wire \this_vga_signals.N_4_1 ;
    wire \this_vga_signals.g3_cascade_ ;
    wire \this_vga_signals.N_5_1 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_0_0_1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_0_0_1 ;
    wire \this_vga_signals.N_1264 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire this_vga_signals_M_vcounter_q_8;
    wire N_1001_0;
    wire N_814_0;
    wire N_1001_0_cascade_;
    wire this_vga_signals_M_vcounter_q_9;
    wire \this_vga_signals.g4 ;
    wire \this_ppu.N_1278_cascade_ ;
    wire \this_ppu.N_767_0 ;
    wire \this_ppu.N_1425 ;
    wire \this_ppu.N_1149_cascade_ ;
    wire \this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1Z0Z_0 ;
    wire \this_ppu.M_this_state_q_srsts_0_0_0_tz_0_0 ;
    wire M_this_state_qZ0Z_8;
    wire N_815_0;
    wire led_c_7;
    wire \this_ppu.N_807_0 ;
    wire M_this_state_qZ0Z_16;
    wire N_1415;
    wire N_1415_cascade_;
    wire \this_ppu.N_1278 ;
    wire \this_ppu.N_1166 ;
    wire \this_ppu.N_1263_cascade_ ;
    wire \this_ppu.N_1176_1 ;
    wire \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_3 ;
    wire \this_ppu.N_893 ;
    wire \this_ppu.N_969 ;
    wire un1_M_this_state_q_11_0_0_cascade_;
    wire \this_ppu.un1_M_this_state_q_11_0_0Z0Z_0_cascade_ ;
    wire \this_ppu.un1_M_this_state_q_11_0_0Z0Z_1 ;
    wire \this_ppu.N_430_1_0 ;
    wire \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_2 ;
    wire \this_ppu.N_1158_cascade_ ;
    wire \this_ppu.N_1263 ;
    wire port_address_in_4;
    wire port_address_in_0;
    wire port_rw_in;
    wire N_1422;
    wire M_this_spr_address_qZ0Z_0;
    wire bfn_22_14_0_;
    wire M_this_spr_address_qZ0Z_1;
    wire un1_M_this_spr_address_q_cry_0;
    wire M_this_spr_address_qZ0Z_2;
    wire un1_M_this_spr_address_q_cry_1;
    wire M_this_spr_address_qZ0Z_3;
    wire un1_M_this_spr_address_q_cry_2;
    wire M_this_spr_address_qZ0Z_4;
    wire un1_M_this_spr_address_q_cry_3;
    wire M_this_spr_address_qZ0Z_5;
    wire un1_M_this_spr_address_q_cry_4;
    wire M_this_spr_address_qZ0Z_6;
    wire un1_M_this_spr_address_q_cry_5;
    wire M_this_spr_address_qZ0Z_7;
    wire un1_M_this_spr_address_q_cry_6;
    wire un1_M_this_spr_address_q_cry_7;
    wire M_this_spr_address_qZ0Z_8;
    wire bfn_22_15_0_;
    wire M_this_spr_address_qZ0Z_9;
    wire un1_M_this_spr_address_q_cry_8;
    wire M_this_spr_address_qZ0Z_10;
    wire un1_M_this_spr_address_q_cry_9;
    wire un1_M_this_spr_address_q_cry_10;
    wire un1_M_this_spr_address_q_cry_11;
    wire N_1005_0;
    wire un1_M_this_spr_address_q_cry_12;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_5 ;
    wire \this_ppu.oam_cache.mem_6 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_6 ;
    wire \this_spr_ram.mem_out_bus4_2 ;
    wire \this_spr_ram.mem_out_bus0_2 ;
    wire \this_spr_ram.mem_mem_0_1_RNIM6VFZ0_cascade_ ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ;
    wire M_this_spr_ram_read_data_2_cascade_;
    wire M_this_ppu_vram_data_2;
    wire \this_spr_ram.mem_out_bus5_0 ;
    wire \this_spr_ram.mem_out_bus1_0 ;
    wire \this_spr_ram.mem_out_bus4_1 ;
    wire \this_spr_ram.mem_out_bus0_1 ;
    wire \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0_cascade_ ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ;
    wire M_this_spr_ram_read_data_2;
    wire M_this_spr_ram_read_data_1_cascade_;
    wire \this_ppu.N_1000_0 ;
    wire M_this_spr_ram_read_data_1;
    wire M_this_ppu_vram_data_1;
    wire \this_spr_ram.mem_mem_1_0_RNIMA1GZ0 ;
    wire M_this_spr_ram_read_data_0;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire \this_vga_signals.N_1307_0_g ;
    wire \this_vga_signals.N_1637_g ;
    wire \this_vga_signals.N_5_i_0 ;
    wire \this_vga_signals.N_5_i_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_0_1 ;
    wire \this_vga_signals.g0_21_1 ;
    wire \this_vga_signals.mult1_un47_sum_axb1 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_ns ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_3 ;
    wire \this_vga_signals.mult1_un47_sum_1_1 ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.vaddress_5 ;
    wire \this_vga_signals.g2_1_0 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_4 ;
    wire \this_vga_signals.mult1_un47_sum_2_1 ;
    wire \this_vga_signals.mult1_un54_sum_axb1 ;
    wire \this_vga_signals.if_N_7_0_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0 ;
    wire this_vga_signals_M_vcounter_q_4;
    wire this_vga_signals_M_vcounter_q_7;
    wire this_vga_signals_M_vcounter_q_5;
    wire this_vga_signals_M_vcounter_q_6;
    wire \this_vga_signals.vaddress_0_0_7 ;
    wire M_this_scroll_qZ0Z_6;
    wire \this_ppu.M_screen_y_q_esr_RNILD7F7Z0Z_6 ;
    wire M_this_spr_ram_write_data_3;
    wire \this_ppu.M_this_state_q_srsts_0_0_a2_1_xZ0Z_0 ;
    wire \this_ppu.N_798_0 ;
    wire \this_ppu.N_1426 ;
    wire M_this_ppu_vram_data_3;
    wire \this_ppu.N_1257 ;
    wire \this_ppu.N_1322 ;
    wire M_this_spr_ram_write_data_1;
    wire led_c_1;
    wire N_1416_cascade_;
    wire N_1151_3;
    wire \this_ppu.N_787_0 ;
    wire \this_ppu.M_this_state_q_srsts_0_0_a2_1_sxZ0Z_0 ;
    wire M_this_state_qZ0Z_14;
    wire M_this_state_qZ0Z_13;
    wire M_this_spr_ram_write_en_0_i_1_0;
    wire M_this_state_qZ0Z_3;
    wire port_address_in_2;
    wire port_address_in_1;
    wire M_this_substate_qZ0;
    wire this_ppu_M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1;
    wire M_this_map_address_qc_3_0_cascade_;
    wire M_this_state_qZ0Z_10;
    wire N_169_0;
    wire N_1048_i;
    wire \this_spr_ram.mem_out_bus5_1 ;
    wire \this_spr_ram.mem_out_bus1_1 ;
    wire \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0 ;
    wire \this_spr_ram.mem_out_bus5_2 ;
    wire \this_spr_ram.mem_out_bus1_2 ;
    wire \this_spr_ram.mem_mem_1_1_RNIOA1GZ0 ;
    wire \this_spr_ram.mem_out_bus6_0 ;
    wire \this_spr_ram.mem_out_bus2_0 ;
    wire \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_ ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0 ;
    wire \this_spr_ram.mem_WE_0 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7 ;
    wire \this_spr_ram.mem_out_bus6_2 ;
    wire \this_spr_ram.mem_out_bus2_2 ;
    wire \this_spr_ram.mem_mem_2_1_RNIQE3GZ0 ;
    wire \this_spr_ram.mem_out_bus4_3 ;
    wire \this_spr_ram.mem_out_bus0_3 ;
    wire \this_ppu.N_753_0 ;
    wire \this_ppu.M_screen_y_qZ0Z_6 ;
    wire \this_ppu.M_screen_y_qZ0Z_4 ;
    wire \this_ppu.un3_M_screen_y_d_0_c4 ;
    wire N_861_0;
    wire \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_0 ;
    wire \this_ppu.M_screen_y_qZ0Z_5 ;
    wire M_this_scroll_qZ0Z_5;
    wire \this_ppu.M_screen_y_q_esr_RNIJB7F7Z0Z_5 ;
    wire \this_spr_ram.mem_radregZ0Z_12 ;
    wire \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0 ;
    wire \this_spr_ram.mem_radregZ0Z_11 ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ;
    wire M_this_spr_ram_read_data_3;
    wire \this_spr_ram.mem_out_bus5_3 ;
    wire \this_spr_ram.mem_out_bus1_3 ;
    wire \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0 ;
    wire \this_spr_ram.mem_out_bus6_3 ;
    wire \this_spr_ram.mem_out_bus2_3 ;
    wire \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0 ;
    wire \this_spr_ram.mem_out_bus7_0 ;
    wire \this_spr_ram.mem_out_bus3_0 ;
    wire \this_spr_ram.mem_mem_3_0_RNIQI5GZ0 ;
    wire \this_spr_ram.mem_out_bus7_1 ;
    wire \this_spr_ram.mem_out_bus3_1 ;
    wire \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0 ;
    wire \this_spr_ram.mem_out_bus7_2 ;
    wire \this_spr_ram.mem_out_bus3_2 ;
    wire \this_spr_ram.mem_mem_3_1_RNISI5GZ0 ;
    wire \this_spr_ram.mem_out_bus7_3 ;
    wire \this_spr_ram.mem_out_bus3_3 ;
    wire \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0 ;
    wire M_this_ctrl_flags_qZ0Z_7;
    wire M_this_state_qZ0Z_2;
    wire N_38_i_0;
    wire N_38_i_0_i;
    wire \this_ppu.N_856_0 ;
    wire this_ppu_un1_M_this_state_q_7_i_0_0_0_cascade_;
    wire N_816_0;
    wire N_1416;
    wire M_this_state_qZ0Z_5;
    wire led_c_6;
    wire M_this_state_qZ0Z_6;
    wire this_ppu_un1_M_this_state_q_7_i_0_0_0;
    wire un1_M_this_state_q_7_i_0_a3_0_0_cascade_;
    wire \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0 ;
    wire M_this_map_ram_read_data_0;
    wire \this_ppu.N_785_0 ;
    wire read_data_RNI4PFJ1_0;
    wire N_1058;
    wire N_1062_cascade_;
    wire M_this_map_address_qc_5_0;
    wire N_1066;
    wire M_this_map_address_qc_6_0_cascade_;
    wire M_this_state_qZ0Z_4;
    wire N_794_0;
    wire M_this_map_address_qc_4_0;
    wire N_918_0;
    wire m5_i_a2_i_o3_i_a3;
    wire N_1048_i_0;
    wire \this_spr_ram.mem_WE_12 ;
    wire \this_spr_ram.mem_WE_8 ;
    wire \this_spr_ram.mem_WE_14 ;
    wire \this_spr_ram.mem_WE_10 ;
    wire \this_spr_ram.mem_out_bus4_0 ;
    wire \this_spr_ram.mem_out_bus0_0 ;
    wire \this_spr_ram.mem_mem_0_0_RNIK6VFZ0 ;
    wire \this_spr_ram.mem_out_bus2_1 ;
    wire \this_spr_ram.mem_radregZ0Z_13 ;
    wire \this_spr_ram.mem_out_bus6_1 ;
    wire \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0 ;
    wire M_this_map_ram_read_data_7;
    wire IO_port_data_write_i_m2_i_m2_7;
    wire \this_spr_ram.mem_WE_6 ;
    wire \this_spr_ram.mem_WE_4 ;
    wire M_this_spr_address_qZ0Z_12;
    wire M_this_spr_address_qZ0Z_11;
    wire M_this_spr_address_qZ0Z_13;
    wire M_this_spr_ram_write_en_0_i_1_0_0;
    wire \this_spr_ram.mem_WE_2 ;
    wire N_842_0;
    wire M_this_status_flags_qZ0Z_7;
    wire M_this_map_address_qc_3_1;
    wire un1_M_this_map_address_q_cry_0_c_RNOZ0;
    wire bfn_24_23_0_;
    wire M_this_map_address_qZ0Z_1;
    wire un1_M_this_map_address_q_cry_0_THRU_CO;
    wire un1_M_this_map_address_q_cry_0;
    wire M_this_map_address_qZ0Z_2;
    wire M_this_map_address_q_RNO_1Z0Z_2;
    wire un1_M_this_map_address_q_cry_1;
    wire M_this_map_address_qZ0Z_3;
    wire M_this_map_address_q_RNO_1Z0Z_3;
    wire un1_M_this_map_address_q_cry_2;
    wire M_this_map_address_qZ0Z_4;
    wire M_this_map_address_q_RNO_1Z0Z_4;
    wire un1_M_this_map_address_q_cry_3;
    wire un1_M_this_state_q_7_i_0_a3_0_0;
    wire un1_M_this_map_address_q_cry_4;
    wire un1_M_this_map_address_q_cry_5;
    wire un1_M_this_map_address_q_cry_6;
    wire un1_M_this_map_address_q_cry_7;
    wire bfn_24_24_0_;
    wire un1_M_this_map_address_q_cry_8;
    wire un1_M_this_map_address_q_cry_5_THRU_CO;
    wire port_data_in_1;
    wire M_this_map_address_qc_8_1_cascade_;
    wire M_this_map_address_qZ0Z_6;
    wire un1_M_this_map_address_q_cry_7_THRU_CO;
    wire un1_M_this_map_address_q_axb_0;
    wire M_this_map_address_qc_2_0;
    wire N_1097;
    wire M_this_map_address_qZ0Z_0;
    wire N_921_0;
    wire N_919_0;
    wire N_923_0;
    wire N_920_0;
    wire N_922_0;
    wire N_296_0;
    wire N_924_0;
    wire port_data_in_5;
    wire M_this_ctrl_flags_qZ0Z_5;
    wire port_data_in_7;
    wire M_this_ctrl_flags_qZ0Z_6;
    wire port_data_in_6;
    wire N_247;
    wire M_this_ext_address_qZ0Z_0;
    wire bfn_26_21_0_;
    wire un1_M_this_ext_address_q_cry_0;
    wire M_this_ext_address_qZ0Z_2;
    wire un1_M_this_ext_address_q_cry_1_THRU_CO;
    wire un1_M_this_ext_address_q_cry_1;
    wire un1_M_this_ext_address_q_cry_2;
    wire un1_M_this_ext_address_q_cry_3;
    wire un1_M_this_ext_address_q_cry_4;
    wire un1_M_this_ext_address_q_cry_5;
    wire un1_M_this_ext_address_q_cry_6;
    wire un1_M_this_ext_address_q_cry_7;
    wire bfn_26_22_0_;
    wire M_this_ext_address_qZ0Z_9;
    wire un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0;
    wire un1_M_this_ext_address_q_cry_8;
    wire un1_M_this_ext_address_q_cry_9;
    wire un1_M_this_ext_address_q_cry_10;
    wire un1_M_this_ext_address_q_cry_11;
    wire M_this_ext_address_qZ0Z_13;
    wire un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0;
    wire un1_M_this_ext_address_q_cry_12;
    wire M_this_ext_address_qZ0Z_14;
    wire un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0;
    wire un1_M_this_ext_address_q_cry_13;
    wire M_this_ext_address_qZ0Z_15;
    wire un1_M_this_ext_address_q_cry_14;
    wire un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0;
    wire un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0;
    wire M_this_ext_address_qZ0Z_10;
    wire un1_M_this_ext_address_q_cry_6_THRU_CO;
    wire M_this_ext_address_qZ0Z_7;
    wire un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0;
    wire M_this_ext_address_qZ0Z_11;
    wire un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0;
    wire M_this_ext_address_qZ0Z_12;
    wire M_this_state_qZ0Z_1;
    wire M_this_ctrl_flags_qZ0Z_4;
    wire M_this_map_address_qZ0Z_9;
    wire port_data_in_4;
    wire N_1081_cascade_;
    wire M_this_map_address_qc_1_1;
    wire M_this_map_address_qZ0Z_8;
    wire port_data_in_3;
    wire N_1078_cascade_;
    wire M_this_map_address_qc_0_1;
    wire M_this_map_ram_read_data_2;
    wire N_726_0;
    wire un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0;
    wire M_this_ext_address_qZ0Z_8;
    wire un1_M_this_ext_address_q_cry_0_THRU_CO;
    wire M_this_ext_address_qZ0Z_1;
    wire un1_M_this_ext_address_q_cry_2_THRU_CO;
    wire M_this_ext_address_qZ0Z_3;
    wire un1_M_this_ext_address_q_cry_3_THRU_CO;
    wire M_this_ext_address_qZ0Z_4;
    wire un1_M_this_ext_address_q_cry_4_THRU_CO;
    wire M_this_ext_address_qZ0Z_5;
    wire N_773_0;
    wire N_765_0;
    wire un1_M_this_ext_address_q_cry_5_THRU_CO;
    wire M_this_ext_address_qZ0Z_6;
    wire M_this_reset_cond_out_g_0;
    wire un1_M_this_map_address_q_cry_6_THRU_CO;
    wire M_this_map_address_qZ0Z_7;
    wire N_801_0;
    wire port_data_in_2;
    wire N_1075_cascade_;
    wire M_this_map_address_qc_1_0;
    wire port_address_in_3;
    wire N_459_0;
    wire N_1276;
    wire N_1242;
    wire port_data_in_0;
    wire N_1068;
    wire M_this_map_address_qc_7_1;
    wire M_this_map_address_q_RNO_1Z0Z_5;
    wire N_1258;
    wire M_this_map_address_qZ0Z_5;
    wire clk_0_c_g;
    wire N_620_g;
    wire M_this_map_ram_read_data_6;
    wire N_734_0;
    wire M_this_map_ram_read_data_5;
    wire N_996_0;
    wire port_address_in_6;
    wire port_address_in_5;
    wire port_address_in_7;
    wire M_this_substate_d_0_sqmuxa_3_0_o2_x;
    wire M_this_map_ram_read_data_4;
    wire N_730_0;
    wire \this_vga_signals.N_834_0 ;
    wire M_this_map_ram_read_data_3;
    wire N_728_0;
    wire _gnd_net_;

    defparam \this_map_ram.mem_mem_0_0_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_0_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,M_this_map_ram_read_data_3,dangling_wire_2,dangling_wire_3,dangling_wire_4,M_this_map_ram_read_data_2,dangling_wire_5,dangling_wire_6,dangling_wire_7,M_this_map_ram_read_data_1,dangling_wire_8,dangling_wire_9,dangling_wire_10,M_this_map_ram_read_data_0,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__21724,N__21343,N__21388,N__21427,N__21475,N__21187,N__21259,N__22924,N__23008,N__23416}),
            .WADDR({dangling_wire_13,N__40825,N__41560,N__42886,N__39646,N__42190,N__39244,N__39289,N__39331,N__39388,N__39574}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__40171,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__40186,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__38494,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__36076,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__42140),
            .RE(N__25236),
            .WCLKE(N__40149),
            .WCLK(N__42141),
            .WE(N__25255));
    defparam \this_map_ram.mem_mem_0_1_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_1_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_42,dangling_wire_43,M_this_map_ram_read_data_7,dangling_wire_44,dangling_wire_45,dangling_wire_46,M_this_map_ram_read_data_6,dangling_wire_47,dangling_wire_48,dangling_wire_49,M_this_map_ram_read_data_5,dangling_wire_50,dangling_wire_51,dangling_wire_52,M_this_map_ram_read_data_4,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__21718,N__21337,N__21382,N__21420,N__21469,N__21181,N__21253,N__22918,N__23001,N__23410}),
            .WADDR({dangling_wire_55,N__40819,N__41554,N__42880,N__39640,N__42184,N__39238,N__39283,N__39325,N__39382,N__39568}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__40075,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__40180,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__40165,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__39520,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__42144),
            .RE(N__25259),
            .WCLKE(N__40156),
            .WCLK(N__42145),
            .WE(N__25264));
    defparam \this_oam_ram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_0_physical  (
            .RDATA({M_this_oam_ram_read_data_15,M_this_oam_ram_read_data_14,M_this_oam_ram_read_data_13,M_this_oam_ram_read_data_12,M_this_oam_ram_read_data_11,M_this_oam_ram_read_data_10,M_this_oam_ram_read_data_9,M_this_oam_ram_read_data_8,M_this_oam_ram_read_data_7,M_this_oam_ram_read_data_6,M_this_oam_ram_read_data_5,M_this_oam_ram_read_data_4,M_this_oam_ram_read_data_3,M_this_oam_ram_read_data_2,M_this_oam_ram_read_data_1,M_this_oam_ram_read_data_0}),
            .RADDR({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,N__16678,N__15631,N__15757,N__15694,N__15451,N__16639}),
            .WADDR({dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,N__21814,N__26470,N__26521,N__26932,N__26998,N__26413}),
            .MASK({dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109}),
            .WDATA({N__17098,N__19276,N__19285,N__19294,N__19303,N__16318,N__16549,N__16519,N__17029,N__17050,N__16147,N__18010,N__18028,N__25327,N__18190,N__17230}),
            .RCLKE(),
            .RCLK(N__42117),
            .RE(N__24986),
            .WCLKE(N__26758),
            .WCLK(N__42118),
            .WE(N__24991));
    defparam \this_oam_ram.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_1_physical  (
            .RDATA({M_this_oam_ram_read_data_31,M_this_oam_ram_read_data_30,M_this_oam_ram_read_data_29,M_this_oam_ram_read_data_28,M_this_oam_ram_read_data_27,M_this_oam_ram_read_data_26,M_this_oam_ram_read_data_25,M_this_oam_ram_read_data_24,M_this_oam_ram_read_data_23,M_this_oam_ram_read_data_22,M_this_oam_ram_read_data_21,M_this_oam_ram_read_data_20,M_this_oam_ram_read_data_19,M_this_oam_ram_read_data_18,M_this_oam_ram_read_data_17,M_this_oam_ram_read_data_16}),
            .RADDR({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,N__16672,N__15625,N__15751,N__15688,N__15445,N__16633}),
            .WADDR({dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,N__21808,N__26464,N__26515,N__26926,N__26992,N__26407}),
            .MASK({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .WDATA({N__16507,N__17113,N__17980,N__16528,N__17122,N__17131,N__18178,N__16489,N__15373,N__20221,N__17971,N__15367,N__15361,N__15205,N__15355,N__16498}),
            .RCLKE(),
            .RCLK(N__42127),
            .RE(N__24987),
            .WCLKE(N__26757),
            .WCLK(N__42128),
            .WE(N__25133));
    defparam \this_ppu.oam_cache.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_ppu.oam_cache.mem_mem_0_0_physical  (
            .RDATA({\this_ppu.oam_cache.mem_15 ,\this_ppu.oam_cache.mem_14 ,\this_ppu.oam_cache.mem_13 ,\this_ppu.oam_cache.mem_12 ,\this_ppu.oam_cache.mem_11 ,\this_ppu.oam_cache.mem_10 ,\this_ppu.oam_cache.mem_9 ,\this_ppu.oam_cache.mem_8 ,\this_ppu.oam_cache.mem_7 ,\this_ppu.oam_cache.mem_6 ,\this_ppu.oam_cache.mem_5 ,\this_ppu.oam_cache.mem_4 ,\this_ppu.oam_cache.mem_3 ,\this_ppu.oam_cache.mem_2 ,\this_ppu.oam_cache.mem_1 ,\this_ppu.oam_cache.mem_0 }),
            .RADDR({dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,N__14788,N__14809,N__14824,N__14875}),
            .WADDR({dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,N__15535,N__22657,N__15805,N__16060}),
            .MASK({dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165}),
            .WDATA({N__14737,N__16450,N__13990,N__14614,N__17476,N__14668,N__14689,N__14707,N__14530,N__14725,N__16765,N__16732,N__14731,N__14602,N__21613,N__15301}),
            .RCLKE(),
            .RCLK(N__42060),
            .RE(N__24833),
            .WCLKE(N__24184),
            .WCLK(N__42061),
            .WE(N__24906));
    defparam \this_ppu.oam_cache.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \this_ppu.oam_cache.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,\this_ppu.oam_cache.mem_18 ,\this_ppu.oam_cache.mem_17 ,\this_ppu.oam_cache.mem_16 }),
            .RADDR({dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,N__14782,N__14803,N__14818,N__14869}),
            .WADDR({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,N__15529,N__22650,N__15799,N__16054}),
            .MASK({dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208}),
            .WDATA({N__16363,N__18964,N__16420,N__16282,N__16888,N__14578,N__14974,N__15946,N__21655,N__15031,N__15037,N__17566,N__16351,N__16159,N__16987,N__14662}),
            .RCLKE(),
            .RCLK(N__42084),
            .RE(N__24852),
            .WCLKE(N__24141),
            .WCLK(N__42085),
            .WE(N__24907));
    defparam \this_spr_ram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,\this_spr_ram.mem_out_bus0_1 ,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,\this_spr_ram.mem_out_bus0_0 ,dangling_wire_220,dangling_wire_221,dangling_wire_222}),
            .RADDR({N__19517,N__19715,N__19939,N__18921,N__38080,N__14283,N__14482,N__20129,N__20653,N__20878,N__21111}),
            .WADDR({N__33419,N__33607,N__33891,N__31338,N__31544,N__31713,N__31971,N__32172,N__32390,N__32601,N__32845}),
            .MASK({dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238}),
            .WDATA({dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,N__35965,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,N__28126,dangling_wire_250,dangling_wire_251,dangling_wire_252}),
            .RCLKE(),
            .RCLK(N__41984),
            .RE(N__25263),
            .WCLKE(N__38323),
            .WCLK(N__41985),
            .WE(N__25262));
    defparam \this_spr_ram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,\this_spr_ram.mem_out_bus0_3 ,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,\this_spr_ram.mem_out_bus0_2 ,dangling_wire_264,dangling_wire_265,dangling_wire_266}),
            .RADDR({N__19516,N__19714,N__19938,N__18922,N__38079,N__14284,N__14466,N__20128,N__20605,N__20874,N__21112}),
            .WADDR({N__33443,N__33673,N__33881,N__31337,N__31543,N__31712,N__31962,N__32171,N__32380,N__32602,N__32839}),
            .MASK({dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282}),
            .WDATA({dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,N__34577,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,N__29428,dangling_wire_294,dangling_wire_295,dangling_wire_296}),
            .RCLKE(),
            .RCLK(N__41986),
            .RE(N__25261),
            .WCLKE(N__38322),
            .WCLK(N__41987),
            .WE(N__25247));
    defparam \this_spr_ram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,\this_spr_ram.mem_out_bus1_1 ,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,\this_spr_ram.mem_out_bus1_0 ,dangling_wire_308,dangling_wire_309,dangling_wire_310}),
            .RADDR({N__19501,N__19717,N__19929,N__18917,N__38105,N__14282,N__14409,N__20140,N__20665,N__20867,N__21132}),
            .WADDR({N__33386,N__33658,N__33860,N__31316,N__31526,N__31735,N__31945,N__32150,N__32365,N__32631,N__32823}),
            .MASK({dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326}),
            .WDATA({dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,N__35960,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,N__28122,dangling_wire_338,dangling_wire_339,dangling_wire_340}),
            .RCLKE(),
            .RCLK(N__41988),
            .RE(N__25251),
            .WCLKE(N__38365),
            .WCLK(N__41989),
            .WE(N__25243));
    defparam \this_spr_ram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,\this_spr_ram.mem_out_bus1_3 ,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,\this_spr_ram.mem_out_bus1_2 ,dangling_wire_352,dangling_wire_353,dangling_wire_354}),
            .RADDR({N__19500,N__19713,N__19928,N__18906,N__38104,N__14280,N__14494,N__20139,N__20661,N__20857,N__21103}),
            .WADDR({N__33423,N__33633,N__33830,N__31315,N__31525,N__31708,N__31921,N__32149,N__32342,N__32632,N__32796}),
            .MASK({dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370}),
            .WDATA({dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,N__34576,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,N__29423,dangling_wire_382,dangling_wire_383,dangling_wire_384}),
            .RCLKE(),
            .RCLK(N__41996),
            .RE(N__25138),
            .WCLKE(N__38364),
            .WCLK(N__41995),
            .WE(N__25220));
    defparam \this_spr_ram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,\this_spr_ram.mem_out_bus2_1 ,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,\this_spr_ram.mem_out_bus2_0 ,dangling_wire_396,dangling_wire_397,dangling_wire_398}),
            .RADDR({N__19522,N__19709,N__19905,N__18905,N__38090,N__14269,N__14490,N__20132,N__20654,N__20845,N__21104}),
            .WADDR({N__33372,N__33597,N__33794,N__31282,N__31492,N__31707,N__31888,N__32116,N__32313,N__32579,N__32761}),
            .MASK({dangling_wire_399,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414}),
            .WDATA({dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,N__35950,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,N__28115,dangling_wire_426,dangling_wire_427,dangling_wire_428}),
            .RCLKE(),
            .RCLK(N__42013),
            .RE(N__25206),
            .WCLKE(N__39184),
            .WCLK(N__42014),
            .WE(N__25219));
    defparam \this_spr_ram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,\this_spr_ram.mem_out_bus2_3 ,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,\this_spr_ram.mem_out_bus2_2 ,dangling_wire_440,dangling_wire_441,dangling_wire_442}),
            .RADDR({N__19499,N__19685,N__19869,N__18904,N__38053,N__14268,N__14483,N__20118,N__20642,N__20833,N__21134}),
            .WADDR({N__33432,N__33616,N__33813,N__31241,N__31424,N__31648,N__31830,N__32055,N__32259,N__32537,N__32702}),
            .MASK({dangling_wire_443,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458}),
            .WDATA({dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,N__34553,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,N__29411,dangling_wire_470,dangling_wire_471,dangling_wire_472}),
            .RCLKE(),
            .RCLK(N__42029),
            .RE(N__25205),
            .WCLKE(N__39180),
            .WCLK(N__42030),
            .WE(N__25164));
    defparam \this_spr_ram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,\this_spr_ram.mem_out_bus3_1 ,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,\this_spr_ram.mem_out_bus3_0 ,dangling_wire_484,dangling_wire_485,dangling_wire_486}),
            .RADDR({N__19518,N__19684,N__19937,N__18903,N__38069,N__14267,N__14470,N__20117,N__20620,N__20817,N__21133}),
            .WADDR({N__33403,N__33576,N__33773,N__31242,N__31475,N__31694,N__31869,N__32099,N__32296,N__32613,N__32742}),
            .MASK({dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502}),
            .WDATA({dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,N__35936,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,N__28105,dangling_wire_514,dangling_wire_515,dangling_wire_516}),
            .RCLKE(),
            .RCLK(N__42047),
            .RE(N__25083),
            .WCLKE(N__38346),
            .WCLK(N__42048),
            .WE(N__25142));
    defparam \this_spr_ram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,\this_spr_ram.mem_out_bus3_3 ,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,dangling_wire_526,dangling_wire_527,\this_spr_ram.mem_out_bus3_2 ,dangling_wire_528,dangling_wire_529,dangling_wire_530}),
            .RADDR({N__19498,N__19683,N__19924,N__18916,N__38040,N__14276,N__14446,N__20116,N__20609,N__20790,N__21126}),
            .WADDR({N__33433,N__33649,N__33814,N__31258,N__31476,N__31727,N__31909,N__32100,N__32297,N__32633,N__32782}),
            .MASK({dangling_wire_531,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546}),
            .WDATA({dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,N__34565,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,N__29427,dangling_wire_558,dangling_wire_559,dangling_wire_560}),
            .RCLKE(),
            .RCLK(N__42071),
            .RE(N__25076),
            .WCLKE(N__38347),
            .WCLK(N__42072),
            .WE(N__25084));
    defparam \this_spr_ram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,\this_spr_ram.mem_out_bus4_1 ,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,dangling_wire_570,dangling_wire_571,\this_spr_ram.mem_out_bus4_0 ,dangling_wire_572,dangling_wire_573,dangling_wire_574}),
            .RADDR({N__19509,N__19682,N__19922,N__18899,N__38039,N__14262,N__14364,N__20115,N__20572,N__20757,N__21116}),
            .WADDR({N__33402,N__33620,N__33849,N__31295,N__31514,N__31728,N__31910,N__32138,N__32331,N__32609,N__32783}),
            .MASK({dangling_wire_575,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590}),
            .WDATA({dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,N__35918,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,N__28093,dangling_wire_602,dangling_wire_603,dangling_wire_604}),
            .RCLKE(),
            .RCLK(N__42094),
            .RE(N__25203),
            .WCLKE(N__38961),
            .WCLK(N__42095),
            .WE(N__25110));
    defparam \this_spr_ram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,\this_spr_ram.mem_out_bus4_3 ,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,dangling_wire_614,dangling_wire_615,\this_spr_ram.mem_out_bus4_2 ,dangling_wire_616,dangling_wire_617,dangling_wire_618}),
            .RADDR({N__19485,N__19681,N__19886,N__18895,N__38037,N__14263,N__14458,N__20111,N__20610,N__20802,N__21135}),
            .WADDR({N__33431,N__33650,N__33876,N__31296,N__31515,N__31746,N__31911,N__32139,N__32332,N__32641,N__32815}),
            .MASK({dangling_wire_619,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634}),
            .WDATA({dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,N__34528,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,N__29418,dangling_wire_646,dangling_wire_647,dangling_wire_648}),
            .RCLKE(),
            .RCLK(N__42110),
            .RE(N__25204),
            .WCLKE(N__38962),
            .WCLK(N__42111),
            .WE(N__25176));
    defparam \this_spr_ram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,\this_spr_ram.mem_out_bus5_1 ,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,dangling_wire_658,dangling_wire_659,\this_spr_ram.mem_out_bus5_0 ,dangling_wire_660,dangling_wire_661,dangling_wire_662}),
            .RADDR({N__19486,N__19692,N__19918,N__18896,N__37997,N__14264,N__14459,N__20112,N__20639,N__20803,N__21084}),
            .WADDR({N__33430,N__33651,N__33856,N__31323,N__31538,N__31747,N__31940,N__32166,N__32360,N__32637,N__32816}),
            .MASK({dangling_wire_663,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678}),
            .WDATA({dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,N__35914,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,N__28081,dangling_wire_690,dangling_wire_691,dangling_wire_692}),
            .RCLKE(),
            .RCLK(N__42121),
            .RE(N__25059),
            .WCLKE(N__38943),
            .WCLK(N__42122),
            .WE(N__25177));
    defparam \this_spr_ram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,\this_spr_ram.mem_out_bus5_3 ,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,dangling_wire_702,dangling_wire_703,\this_spr_ram.mem_out_bus5_2 ,dangling_wire_704,dangling_wire_705,dangling_wire_706}),
            .RADDR({N__19496,N__19693,N__19923,N__18897,N__38038,N__14265,N__14480,N__20113,N__20640,N__20829,N__21083}),
            .WADDR({N__33453,N__33669,N__33890,N__31324,N__31539,N__31714,N__31941,N__32170,N__32361,N__32630,N__32837}),
            .MASK({dangling_wire_707,dangling_wire_708,dangling_wire_709,dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722}),
            .WDATA({dangling_wire_723,dangling_wire_724,dangling_wire_725,dangling_wire_726,N__34566,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,N__29375,dangling_wire_734,dangling_wire_735,dangling_wire_736}),
            .RCLKE(),
            .RCLK(N__42130),
            .RE(N__25060),
            .WCLKE(N__38944),
            .WCLK(N__42131),
            .WE(N__25227));
    defparam \this_spr_ram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,\this_spr_ram.mem_out_bus6_1 ,dangling_wire_741,dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,dangling_wire_746,dangling_wire_747,\this_spr_ram.mem_out_bus6_0 ,dangling_wire_748,dangling_wire_749,dangling_wire_750}),
            .RADDR({N__19497,N__19694,N__19936,N__18898,N__38068,N__14266,N__14481,N__20114,N__20641,N__20830,N__21082}),
            .WADDR({N__33444,N__33678,N__33880,N__31339,N__31546,N__31736,N__31961,N__32182,N__32379,N__32623,N__32838}),
            .MASK({dangling_wire_751,dangling_wire_752,dangling_wire_753,dangling_wire_754,dangling_wire_755,dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766}),
            .WDATA({dangling_wire_767,dangling_wire_768,dangling_wire_769,dangling_wire_770,N__35949,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,N__28080,dangling_wire_778,dangling_wire_779,dangling_wire_780}),
            .RCLKE(),
            .RCLK(N__42135),
            .RE(N__25235),
            .WCLKE(N__38646),
            .WCLK(N__42136),
            .WE(N__25228));
    defparam \this_spr_ram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,\this_spr_ram.mem_out_bus6_3 ,dangling_wire_785,dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,dangling_wire_790,dangling_wire_791,\this_spr_ram.mem_out_bus6_2 ,dangling_wire_792,dangling_wire_793,dangling_wire_794}),
            .RADDR({N__19480,N__19704,N__19843,N__18850,N__38097,N__14257,N__14385,N__20104,N__20632,N__20810,N__21127}),
            .WADDR({N__33452,N__33662,N__33885,N__31340,N__31533,N__31748,N__31966,N__32183,N__32372,N__32634,N__32830}),
            .MASK({dangling_wire_795,dangling_wire_796,dangling_wire_797,dangling_wire_798,dangling_wire_799,dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810}),
            .WDATA({dangling_wire_811,dangling_wire_812,dangling_wire_813,dangling_wire_814,N__34578,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,N__29407,dangling_wire_822,dangling_wire_823,dangling_wire_824}),
            .RCLKE(),
            .RCLK(N__42133),
            .RE(N__24999),
            .WCLKE(N__38650),
            .WCLK(N__42134),
            .WE(N__25134));
    defparam \this_spr_ram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,\this_spr_ram.mem_out_bus7_1 ,dangling_wire_829,dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,dangling_wire_834,dangling_wire_835,\this_spr_ram.mem_out_bus7_0 ,dangling_wire_836,dangling_wire_837,dangling_wire_838}),
            .RADDR({N__19481,N__19705,N__19844,N__18894,N__38106,N__14258,N__14386,N__20130,N__20565,N__20831,N__21128}),
            .WADDR({N__33448,N__33674,N__33886,N__31347,N__31534,N__31755,N__31970,N__32187,N__32391,N__32635,N__32843}),
            .MASK({dangling_wire_839,dangling_wire_840,dangling_wire_841,dangling_wire_842,dangling_wire_843,dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854}),
            .WDATA({dangling_wire_855,dangling_wire_856,dangling_wire_857,dangling_wire_858,N__35964,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,N__28114,dangling_wire_866,dangling_wire_867,dangling_wire_868}),
            .RCLKE(),
            .RCLK(N__42138),
            .RE(N__25061),
            .WCLKE(N__36702),
            .WCLK(N__42139),
            .WE(N__25071));
    defparam \this_spr_ram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_869,dangling_wire_870,dangling_wire_871,dangling_wire_872,\this_spr_ram.mem_out_bus7_3 ,dangling_wire_873,dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,dangling_wire_878,dangling_wire_879,\this_spr_ram.mem_out_bus7_2 ,dangling_wire_880,dangling_wire_881,dangling_wire_882}),
            .RADDR({N__19508,N__19716,N__19885,N__18854,N__38107,N__14281,N__14416,N__20131,N__20652,N__20832,N__21139}),
            .WADDR({N__33454,N__33679,N__33892,N__31348,N__31545,N__31756,N__31972,N__32188,N__32395,N__32636,N__32844}),
            .MASK({dangling_wire_883,dangling_wire_884,dangling_wire_885,dangling_wire_886,dangling_wire_887,dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898}),
            .WDATA({dangling_wire_899,dangling_wire_900,dangling_wire_901,dangling_wire_902,N__34582,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,N__29422,dangling_wire_910,dangling_wire_911,dangling_wire_912}),
            .RCLKE(),
            .RCLK(N__42142),
            .RE(N__25072),
            .WCLKE(N__36706),
            .WCLK(N__42143),
            .WE(N__25199));
    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_913,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917,dangling_wire_918,dangling_wire_919,dangling_wire_920,dangling_wire_921,dangling_wire_922,dangling_wire_923,dangling_wire_924,M_this_vram_read_data_3,M_this_vram_read_data_2,M_this_vram_read_data_1,M_this_vram_read_data_0}),
            .RADDR({dangling_wire_925,dangling_wire_926,dangling_wire_927,N__23854,N__15466,N__18043,N__17539,N__16012,N__14839,N__16078,N__15883}),
            .WADDR({dangling_wire_928,dangling_wire_929,dangling_wire_930,N__22411,N__22267,N__22294,N__22330,N__23179,N__22243,N__23545,N__23512}),
            .MASK({dangling_wire_931,dangling_wire_932,dangling_wire_933,dangling_wire_934,dangling_wire_935,dangling_wire_936,dangling_wire_937,dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,dangling_wire_943,dangling_wire_944,dangling_wire_945,dangling_wire_946}),
            .WDATA({dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953,dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,dangling_wire_958,N__34405,N__33979,N__34330,N__23125}),
            .RCLKE(),
            .RCLK(N__42103),
            .RE(N__24923),
            .WCLKE(N__23035),
            .WCLK(N__42104),
            .WE(N__24870));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__44414),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__44416),
            .DIN(N__44415),
            .DOUT(N__44414),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__44416),
            .PADOUT(N__44415),
            .PADIN(N__44414),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__44405),
            .DIN(N__44404),
            .DOUT(N__44403),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__44405),
            .PADOUT(N__44404),
            .PADIN(N__44403),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__44396),
            .DIN(N__44395),
            .DOUT(N__44394),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__44396),
            .PADOUT(N__44395),
            .PADIN(N__44394),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__44387),
            .DIN(N__44386),
            .DOUT(N__44385),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__44387),
            .PADOUT(N__44386),
            .PADIN(N__44385),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14569),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__44378),
            .DIN(N__44377),
            .DOUT(N__44376),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__44378),
            .PADOUT(N__44377),
            .PADIN(N__44376),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__16306),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_0_iopad (
            .OE(N__44369),
            .DIN(N__44368),
            .DOUT(N__44367),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__44369),
            .PADOUT(N__44368),
            .PADIN(N__44367),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__25260),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_1_iopad (
            .OE(N__44360),
            .DIN(N__44359),
            .DOUT(N__44358),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__44360),
            .PADOUT(N__44359),
            .PADIN(N__44358),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__35863),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_2_iopad (
            .OE(N__44351),
            .DIN(N__44350),
            .DOUT(N__44349),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__44351),
            .PADOUT(N__44350),
            .PADIN(N__44349),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_3_iopad (
            .OE(N__44342),
            .DIN(N__44341),
            .DOUT(N__44340),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__44342),
            .PADOUT(N__44341),
            .PADIN(N__44340),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_4_iopad (
            .OE(N__44333),
            .DIN(N__44332),
            .DOUT(N__44331),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__44333),
            .PADOUT(N__44332),
            .PADIN(N__44331),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_5_iopad (
            .OE(N__44324),
            .DIN(N__44323),
            .DOUT(N__44322),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__44324),
            .PADOUT(N__44323),
            .PADIN(N__44322),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__36064),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_6_iopad (
            .OE(N__44315),
            .DIN(N__44314),
            .DOUT(N__44313),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__44315),
            .PADOUT(N__44314),
            .PADIN(N__44313),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37360),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_7_iopad (
            .OE(N__44306),
            .DIN(N__44305),
            .DOUT(N__44304),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__44306),
            .PADOUT(N__44305),
            .PADIN(N__44304),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__30871),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__44297),
            .DIN(N__44296),
            .DOUT(N__44295),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__44297),
            .PADOUT(N__44296),
            .PADIN(N__44295),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__40291),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37607));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__44288),
            .DIN(N__44287),
            .DOUT(N__44286),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__44288),
            .PADOUT(N__44287),
            .PADIN(N__44286),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__41305),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37585));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__44279),
            .DIN(N__44278),
            .DOUT(N__44277),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__44279),
            .PADOUT(N__44278),
            .PADIN(N__44277),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__40246),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37576));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__44270),
            .DIN(N__44269),
            .DOUT(N__44268),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__44270),
            .PADOUT(N__44269),
            .PADIN(N__44268),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__41266),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37622));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__44261),
            .DIN(N__44260),
            .DOUT(N__44259),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__44261),
            .PADOUT(N__44260),
            .PADIN(N__44259),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__41227),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37611));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__44252),
            .DIN(N__44251),
            .DOUT(N__44250),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__44252),
            .PADOUT(N__44251),
            .PADIN(N__44250),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__41191),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37561));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__44243),
            .DIN(N__44242),
            .DOUT(N__44241),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__44243),
            .PADOUT(N__44242),
            .PADIN(N__44241),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__43279),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37606));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__44234),
            .DIN(N__44233),
            .DOUT(N__44232),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__44234),
            .PADOUT(N__44233),
            .PADIN(N__44232),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__40984),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37639));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__44225),
            .DIN(N__44224),
            .DOUT(N__44223),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__44225),
            .PADOUT(N__44224),
            .PADIN(N__44223),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__41020),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37577));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__44216),
            .DIN(N__44215),
            .DOUT(N__44214),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__44216),
            .PADOUT(N__44215),
            .PADIN(N__44214),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__40942),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37609));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__44207),
            .DIN(N__44206),
            .DOUT(N__44205),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__44207),
            .PADOUT(N__44206),
            .PADIN(N__44205),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__40912),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37612));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__44198),
            .DIN(N__44197),
            .DOUT(N__44196),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__44198),
            .PADOUT(N__44197),
            .PADIN(N__44196),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__40582),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37562));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__44189),
            .DIN(N__44188),
            .DOUT(N__44187),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__44189),
            .PADOUT(N__44188),
            .PADIN(N__44187),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__40543),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37623));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__44180),
            .DIN(N__44179),
            .DOUT(N__44178),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__44180),
            .PADOUT(N__44179),
            .PADIN(N__44178),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__40507),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37635));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__44171),
            .DIN(N__44170),
            .DOUT(N__44169),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__44171),
            .PADOUT(N__44170),
            .PADIN(N__44169),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__41335),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37608));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__44162),
            .DIN(N__44161),
            .DOUT(N__44160),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__44162),
            .PADOUT(N__44161),
            .PADIN(N__44160),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__40636),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37584));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__44153),
            .DIN(N__44152),
            .DOUT(N__44151),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__44153),
            .PADOUT(N__44152),
            .PADIN(N__44151),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_iobuf_0_iopad (
            .OE(N__44144),
            .DIN(N__44143),
            .DOUT(N__44142),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_data_iobuf_0_preio (
            .PADOEN(N__44144),
            .PADOUT(N__44143),
            .PADIN(N__44142),
            .CLOCKENABLE(),
            .DIN0(port_data_in_0),
            .DIN1(),
            .DOUT0(N__21787),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38437));
    IO_PAD port_data_iobuf_1_iopad (
            .OE(N__44135),
            .DIN(N__44134),
            .DOUT(N__44133),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_data_iobuf_1_preio (
            .PADOEN(N__44135),
            .PADOUT(N__44134),
            .PADIN(N__44133),
            .CLOCKENABLE(),
            .DIN0(port_data_in_1),
            .DIN1(),
            .DOUT0(N__20173),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38438));
    IO_PAD port_data_iobuf_2_iopad (
            .OE(N__44126),
            .DIN(N__44125),
            .DOUT(N__44124),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_data_iobuf_2_preio (
            .PADOEN(N__44126),
            .PADOUT(N__44125),
            .PADIN(N__44124),
            .CLOCKENABLE(),
            .DIN0(port_data_in_2),
            .DIN1(),
            .DOUT0(N__41350),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38401));
    IO_PAD port_data_iobuf_3_iopad (
            .OE(N__44117),
            .DIN(N__44116),
            .DOUT(N__44115),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_data_iobuf_3_preio (
            .PADOEN(N__44117),
            .PADOUT(N__44116),
            .PADIN(N__44115),
            .CLOCKENABLE(),
            .DIN0(port_data_in_3),
            .DIN1(),
            .DOUT0(N__43588),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38413));
    IO_PAD port_data_iobuf_4_iopad (
            .OE(N__44108),
            .DIN(N__44107),
            .DOUT(N__44106),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_data_iobuf_4_preio (
            .PADOEN(N__44108),
            .PADOUT(N__44107),
            .PADIN(N__44106),
            .CLOCKENABLE(),
            .DIN0(port_data_in_4),
            .DIN1(),
            .DOUT0(N__43714),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38431));
    IO_PAD port_data_iobuf_5_iopad (
            .OE(N__44099),
            .DIN(N__44098),
            .DOUT(N__44097),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_data_iobuf_5_preio (
            .PADOEN(N__44099),
            .PADOUT(N__44098),
            .PADIN(N__44097),
            .CLOCKENABLE(),
            .DIN0(port_data_in_5),
            .DIN1(),
            .DOUT0(N__43903),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38445));
    IO_PAD port_data_iobuf_6_iopad (
            .OE(N__44090),
            .DIN(N__44089),
            .DOUT(N__44088),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_data_iobuf_6_preio (
            .PADOEN(N__44090),
            .PADOUT(N__44089),
            .PADIN(N__44088),
            .CLOCKENABLE(),
            .DIN0(port_data_in_6),
            .DIN1(),
            .DOUT0(N__41575),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38457));
    IO_PAD port_data_iobuf_7_iopad (
            .OE(N__44081),
            .DIN(N__44080),
            .DOUT(N__44079),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_data_iobuf_7_preio (
            .PADOEN(N__44081),
            .PADOUT(N__44080),
            .PADIN(N__44079),
            .CLOCKENABLE(),
            .DIN0(port_data_in_7),
            .DIN1(),
            .DOUT0(N__38983),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38461));
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__44072),
            .DIN(N__44071),
            .DOUT(N__44070),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__44072),
            .PADOUT(N__44071),
            .PADIN(N__44070),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14062),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__44063),
            .DIN(N__44062),
            .DOUT(N__44061),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__44063),
            .PADOUT(N__44062),
            .PADIN(N__44061),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37762),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__44054),
            .DIN(N__44053),
            .DOUT(N__44052),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__44054),
            .PADOUT(N__44053),
            .PADIN(N__44052),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__44045),
            .DIN(N__44044),
            .DOUT(N__44043),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__44045),
            .PADOUT(N__44044),
            .PADIN(N__44043),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14020),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__44036),
            .DIN(N__44035),
            .DOUT(N__44034),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__44036),
            .PADOUT(N__44035),
            .PADIN(N__44034),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__24869),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__37610));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__44027),
            .DIN(N__44026),
            .DOUT(N__44025),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__44027),
            .PADOUT(N__44026),
            .PADIN(N__44025),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14770),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__44018),
            .DIN(N__44017),
            .DOUT(N__44016),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__44018),
            .PADOUT(N__44017),
            .PADIN(N__44016),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__15349),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__44009),
            .DIN(N__44008),
            .DOUT(N__44007),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__44009),
            .PADOUT(N__44008),
            .PADIN(N__44007),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13978),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__44000),
            .DIN(N__43999),
            .DOUT(N__43998),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__44000),
            .PADOUT(N__43999),
            .PADIN(N__43998),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__16699),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__43991),
            .DIN(N__43990),
            .DOUT(N__43989),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__43991),
            .PADOUT(N__43990),
            .PADIN(N__43989),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14044),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__43982),
            .DIN(N__43981),
            .DOUT(N__43980),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__43982),
            .PADOUT(N__43981),
            .PADIN(N__43980),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14551),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__43973),
            .DIN(N__43972),
            .DOUT(N__43971),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__43973),
            .PADOUT(N__43972),
            .PADIN(N__43971),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__43964),
            .DIN(N__43963),
            .DOUT(N__43962),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__43964),
            .PADOUT(N__43963),
            .PADIN(N__43962),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14056),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__43955),
            .DIN(N__43954),
            .DOUT(N__43953),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__43955),
            .PADOUT(N__43954),
            .PADIN(N__43953),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22441),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__11033 (
            .O(N__43936),
            .I(N__43932));
    InMux I__11032 (
            .O(N__43935),
            .I(N__43929));
    LocalMux I__11031 (
            .O(N__43932),
            .I(N__43926));
    LocalMux I__11030 (
            .O(N__43929),
            .I(N__43923));
    Span4Mux_v I__11029 (
            .O(N__43926),
            .I(N__43920));
    Span4Mux_h I__11028 (
            .O(N__43923),
            .I(N__43917));
    Span4Mux_h I__11027 (
            .O(N__43920),
            .I(N__43912));
    Span4Mux_v I__11026 (
            .O(N__43917),
            .I(N__43912));
    Span4Mux_v I__11025 (
            .O(N__43912),
            .I(N__43909));
    Span4Mux_v I__11024 (
            .O(N__43909),
            .I(N__43906));
    Odrv4 I__11023 (
            .O(N__43906),
            .I(M_this_map_ram_read_data_5));
    IoInMux I__11022 (
            .O(N__43903),
            .I(N__43900));
    LocalMux I__11021 (
            .O(N__43900),
            .I(N__43897));
    Odrv12 I__11020 (
            .O(N__43897),
            .I(N_996_0));
    CascadeMux I__11019 (
            .O(N__43894),
            .I(N__43891));
    InMux I__11018 (
            .O(N__43891),
            .I(N__43888));
    LocalMux I__11017 (
            .O(N__43888),
            .I(N__43884));
    CascadeMux I__11016 (
            .O(N__43887),
            .I(N__43881));
    Span4Mux_h I__11015 (
            .O(N__43884),
            .I(N__43878));
    InMux I__11014 (
            .O(N__43881),
            .I(N__43875));
    Span4Mux_h I__11013 (
            .O(N__43878),
            .I(N__43869));
    LocalMux I__11012 (
            .O(N__43875),
            .I(N__43869));
    InMux I__11011 (
            .O(N__43874),
            .I(N__43866));
    Sp12to4 I__11010 (
            .O(N__43869),
            .I(N__43861));
    LocalMux I__11009 (
            .O(N__43866),
            .I(N__43861));
    Span12Mux_v I__11008 (
            .O(N__43861),
            .I(N__43858));
    Odrv12 I__11007 (
            .O(N__43858),
            .I(port_address_in_6));
    InMux I__11006 (
            .O(N__43855),
            .I(N__43851));
    InMux I__11005 (
            .O(N__43854),
            .I(N__43848));
    LocalMux I__11004 (
            .O(N__43851),
            .I(N__43844));
    LocalMux I__11003 (
            .O(N__43848),
            .I(N__43841));
    InMux I__11002 (
            .O(N__43847),
            .I(N__43838));
    Span4Mux_v I__11001 (
            .O(N__43844),
            .I(N__43835));
    Span4Mux_v I__11000 (
            .O(N__43841),
            .I(N__43832));
    LocalMux I__10999 (
            .O(N__43838),
            .I(N__43829));
    Sp12to4 I__10998 (
            .O(N__43835),
            .I(N__43826));
    Span4Mux_h I__10997 (
            .O(N__43832),
            .I(N__43823));
    Span4Mux_v I__10996 (
            .O(N__43829),
            .I(N__43820));
    Odrv12 I__10995 (
            .O(N__43826),
            .I(port_address_in_5));
    Odrv4 I__10994 (
            .O(N__43823),
            .I(port_address_in_5));
    Odrv4 I__10993 (
            .O(N__43820),
            .I(port_address_in_5));
    InMux I__10992 (
            .O(N__43813),
            .I(N__43810));
    LocalMux I__10991 (
            .O(N__43810),
            .I(N__43807));
    Span4Mux_v I__10990 (
            .O(N__43807),
            .I(N__43803));
    InMux I__10989 (
            .O(N__43806),
            .I(N__43800));
    Span4Mux_h I__10988 (
            .O(N__43803),
            .I(N__43796));
    LocalMux I__10987 (
            .O(N__43800),
            .I(N__43793));
    InMux I__10986 (
            .O(N__43799),
            .I(N__43790));
    Span4Mux_v I__10985 (
            .O(N__43796),
            .I(N__43787));
    Span4Mux_h I__10984 (
            .O(N__43793),
            .I(N__43784));
    LocalMux I__10983 (
            .O(N__43790),
            .I(N__43781));
    Sp12to4 I__10982 (
            .O(N__43787),
            .I(N__43778));
    Sp12to4 I__10981 (
            .O(N__43784),
            .I(N__43775));
    Span12Mux_v I__10980 (
            .O(N__43781),
            .I(N__43772));
    Span12Mux_s2_h I__10979 (
            .O(N__43778),
            .I(N__43767));
    Span12Mux_v I__10978 (
            .O(N__43775),
            .I(N__43767));
    Span12Mux_v I__10977 (
            .O(N__43772),
            .I(N__43764));
    Span12Mux_v I__10976 (
            .O(N__43767),
            .I(N__43761));
    Odrv12 I__10975 (
            .O(N__43764),
            .I(port_address_in_7));
    Odrv12 I__10974 (
            .O(N__43761),
            .I(port_address_in_7));
    InMux I__10973 (
            .O(N__43756),
            .I(N__43753));
    LocalMux I__10972 (
            .O(N__43753),
            .I(N__43750));
    Odrv12 I__10971 (
            .O(N__43750),
            .I(M_this_substate_d_0_sqmuxa_3_0_o2_x));
    InMux I__10970 (
            .O(N__43747),
            .I(N__43743));
    InMux I__10969 (
            .O(N__43746),
            .I(N__43740));
    LocalMux I__10968 (
            .O(N__43743),
            .I(N__43737));
    LocalMux I__10967 (
            .O(N__43740),
            .I(N__43734));
    Span4Mux_h I__10966 (
            .O(N__43737),
            .I(N__43731));
    Span4Mux_v I__10965 (
            .O(N__43734),
            .I(N__43728));
    Sp12to4 I__10964 (
            .O(N__43731),
            .I(N__43725));
    Span4Mux_v I__10963 (
            .O(N__43728),
            .I(N__43722));
    Span12Mux_v I__10962 (
            .O(N__43725),
            .I(N__43719));
    Odrv4 I__10961 (
            .O(N__43722),
            .I(M_this_map_ram_read_data_4));
    Odrv12 I__10960 (
            .O(N__43719),
            .I(M_this_map_ram_read_data_4));
    IoInMux I__10959 (
            .O(N__43714),
            .I(N__43711));
    LocalMux I__10958 (
            .O(N__43711),
            .I(N__43708));
    Odrv12 I__10957 (
            .O(N__43708),
            .I(N_730_0));
    InMux I__10956 (
            .O(N__43705),
            .I(N__43700));
    InMux I__10955 (
            .O(N__43704),
            .I(N__43697));
    InMux I__10954 (
            .O(N__43703),
            .I(N__43692));
    LocalMux I__10953 (
            .O(N__43700),
            .I(N__43687));
    LocalMux I__10952 (
            .O(N__43697),
            .I(N__43687));
    InMux I__10951 (
            .O(N__43696),
            .I(N__43682));
    InMux I__10950 (
            .O(N__43695),
            .I(N__43682));
    LocalMux I__10949 (
            .O(N__43692),
            .I(N__43678));
    Span4Mux_v I__10948 (
            .O(N__43687),
            .I(N__43675));
    LocalMux I__10947 (
            .O(N__43682),
            .I(N__43672));
    InMux I__10946 (
            .O(N__43681),
            .I(N__43669));
    Span4Mux_v I__10945 (
            .O(N__43678),
            .I(N__43666));
    Span4Mux_v I__10944 (
            .O(N__43675),
            .I(N__43659));
    Span4Mux_v I__10943 (
            .O(N__43672),
            .I(N__43659));
    LocalMux I__10942 (
            .O(N__43669),
            .I(N__43656));
    Span4Mux_h I__10941 (
            .O(N__43666),
            .I(N__43653));
    InMux I__10940 (
            .O(N__43665),
            .I(N__43650));
    InMux I__10939 (
            .O(N__43664),
            .I(N__43647));
    Span4Mux_h I__10938 (
            .O(N__43659),
            .I(N__43642));
    Span4Mux_v I__10937 (
            .O(N__43656),
            .I(N__43642));
    Span4Mux_h I__10936 (
            .O(N__43653),
            .I(N__43639));
    LocalMux I__10935 (
            .O(N__43650),
            .I(N__43636));
    LocalMux I__10934 (
            .O(N__43647),
            .I(N__43633));
    Sp12to4 I__10933 (
            .O(N__43642),
            .I(N__43630));
    Span4Mux_h I__10932 (
            .O(N__43639),
            .I(N__43623));
    Span4Mux_v I__10931 (
            .O(N__43636),
            .I(N__43623));
    Span4Mux_v I__10930 (
            .O(N__43633),
            .I(N__43623));
    Span12Mux_h I__10929 (
            .O(N__43630),
            .I(N__43620));
    Span4Mux_v I__10928 (
            .O(N__43623),
            .I(N__43617));
    Odrv12 I__10927 (
            .O(N__43620),
            .I(\this_vga_signals.N_834_0 ));
    Odrv4 I__10926 (
            .O(N__43617),
            .I(\this_vga_signals.N_834_0 ));
    InMux I__10925 (
            .O(N__43612),
            .I(N__43609));
    LocalMux I__10924 (
            .O(N__43609),
            .I(N__43605));
    InMux I__10923 (
            .O(N__43608),
            .I(N__43602));
    Span12Mux_v I__10922 (
            .O(N__43605),
            .I(N__43599));
    LocalMux I__10921 (
            .O(N__43602),
            .I(N__43596));
    Span12Mux_h I__10920 (
            .O(N__43599),
            .I(N__43593));
    Odrv4 I__10919 (
            .O(N__43596),
            .I(M_this_map_ram_read_data_3));
    Odrv12 I__10918 (
            .O(N__43593),
            .I(M_this_map_ram_read_data_3));
    IoInMux I__10917 (
            .O(N__43588),
            .I(N__43585));
    LocalMux I__10916 (
            .O(N__43585),
            .I(N__43582));
    Span4Mux_s1_v I__10915 (
            .O(N__43582),
            .I(N__43579));
    Odrv4 I__10914 (
            .O(N__43579),
            .I(N_728_0));
    CascadeMux I__10913 (
            .O(N__43576),
            .I(N__43569));
    CascadeMux I__10912 (
            .O(N__43575),
            .I(N__43558));
    CascadeMux I__10911 (
            .O(N__43574),
            .I(N__43555));
    CascadeMux I__10910 (
            .O(N__43573),
            .I(N__43552));
    CascadeMux I__10909 (
            .O(N__43572),
            .I(N__43549));
    InMux I__10908 (
            .O(N__43569),
            .I(N__43530));
    InMux I__10907 (
            .O(N__43568),
            .I(N__43530));
    InMux I__10906 (
            .O(N__43567),
            .I(N__43530));
    InMux I__10905 (
            .O(N__43566),
            .I(N__43530));
    InMux I__10904 (
            .O(N__43565),
            .I(N__43530));
    InMux I__10903 (
            .O(N__43564),
            .I(N__43530));
    InMux I__10902 (
            .O(N__43563),
            .I(N__43517));
    InMux I__10901 (
            .O(N__43562),
            .I(N__43517));
    InMux I__10900 (
            .O(N__43561),
            .I(N__43517));
    InMux I__10899 (
            .O(N__43558),
            .I(N__43517));
    InMux I__10898 (
            .O(N__43555),
            .I(N__43517));
    InMux I__10897 (
            .O(N__43552),
            .I(N__43504));
    InMux I__10896 (
            .O(N__43549),
            .I(N__43504));
    InMux I__10895 (
            .O(N__43548),
            .I(N__43504));
    InMux I__10894 (
            .O(N__43547),
            .I(N__43504));
    InMux I__10893 (
            .O(N__43546),
            .I(N__43504));
    InMux I__10892 (
            .O(N__43545),
            .I(N__43504));
    InMux I__10891 (
            .O(N__43544),
            .I(N__43496));
    InMux I__10890 (
            .O(N__43543),
            .I(N__43493));
    LocalMux I__10889 (
            .O(N__43530),
            .I(N__43490));
    CascadeMux I__10888 (
            .O(N__43529),
            .I(N__43481));
    InMux I__10887 (
            .O(N__43528),
            .I(N__43478));
    LocalMux I__10886 (
            .O(N__43517),
            .I(N__43475));
    LocalMux I__10885 (
            .O(N__43504),
            .I(N__43472));
    InMux I__10884 (
            .O(N__43503),
            .I(N__43467));
    InMux I__10883 (
            .O(N__43502),
            .I(N__43464));
    InMux I__10882 (
            .O(N__43501),
            .I(N__43461));
    InMux I__10881 (
            .O(N__43500),
            .I(N__43457));
    InMux I__10880 (
            .O(N__43499),
            .I(N__43454));
    LocalMux I__10879 (
            .O(N__43496),
            .I(N__43447));
    LocalMux I__10878 (
            .O(N__43493),
            .I(N__43447));
    Span4Mux_h I__10877 (
            .O(N__43490),
            .I(N__43447));
    InMux I__10876 (
            .O(N__43489),
            .I(N__43440));
    InMux I__10875 (
            .O(N__43488),
            .I(N__43440));
    InMux I__10874 (
            .O(N__43487),
            .I(N__43440));
    InMux I__10873 (
            .O(N__43486),
            .I(N__43433));
    InMux I__10872 (
            .O(N__43485),
            .I(N__43433));
    InMux I__10871 (
            .O(N__43484),
            .I(N__43433));
    InMux I__10870 (
            .O(N__43481),
            .I(N__43428));
    LocalMux I__10869 (
            .O(N__43478),
            .I(N__43425));
    Span4Mux_v I__10868 (
            .O(N__43475),
            .I(N__43420));
    Span4Mux_h I__10867 (
            .O(N__43472),
            .I(N__43420));
    InMux I__10866 (
            .O(N__43471),
            .I(N__43417));
    InMux I__10865 (
            .O(N__43470),
            .I(N__43412));
    LocalMux I__10864 (
            .O(N__43467),
            .I(N__43405));
    LocalMux I__10863 (
            .O(N__43464),
            .I(N__43405));
    LocalMux I__10862 (
            .O(N__43461),
            .I(N__43405));
    InMux I__10861 (
            .O(N__43460),
            .I(N__43402));
    LocalMux I__10860 (
            .O(N__43457),
            .I(N__43398));
    LocalMux I__10859 (
            .O(N__43454),
            .I(N__43389));
    Span4Mux_v I__10858 (
            .O(N__43447),
            .I(N__43389));
    LocalMux I__10857 (
            .O(N__43440),
            .I(N__43389));
    LocalMux I__10856 (
            .O(N__43433),
            .I(N__43389));
    InMux I__10855 (
            .O(N__43432),
            .I(N__43384));
    InMux I__10854 (
            .O(N__43431),
            .I(N__43384));
    LocalMux I__10853 (
            .O(N__43428),
            .I(N__43381));
    Span4Mux_v I__10852 (
            .O(N__43425),
            .I(N__43378));
    Span4Mux_h I__10851 (
            .O(N__43420),
            .I(N__43373));
    LocalMux I__10850 (
            .O(N__43417),
            .I(N__43373));
    InMux I__10849 (
            .O(N__43416),
            .I(N__43366));
    InMux I__10848 (
            .O(N__43415),
            .I(N__43366));
    LocalMux I__10847 (
            .O(N__43412),
            .I(N__43362));
    Span4Mux_v I__10846 (
            .O(N__43405),
            .I(N__43357));
    LocalMux I__10845 (
            .O(N__43402),
            .I(N__43357));
    InMux I__10844 (
            .O(N__43401),
            .I(N__43351));
    Span4Mux_v I__10843 (
            .O(N__43398),
            .I(N__43344));
    Span4Mux_v I__10842 (
            .O(N__43389),
            .I(N__43344));
    LocalMux I__10841 (
            .O(N__43384),
            .I(N__43344));
    Span4Mux_v I__10840 (
            .O(N__43381),
            .I(N__43341));
    Span4Mux_h I__10839 (
            .O(N__43378),
            .I(N__43338));
    Span4Mux_h I__10838 (
            .O(N__43373),
            .I(N__43335));
    InMux I__10837 (
            .O(N__43372),
            .I(N__43332));
    InMux I__10836 (
            .O(N__43371),
            .I(N__43329));
    LocalMux I__10835 (
            .O(N__43366),
            .I(N__43326));
    InMux I__10834 (
            .O(N__43365),
            .I(N__43323));
    Span4Mux_h I__10833 (
            .O(N__43362),
            .I(N__43318));
    Span4Mux_h I__10832 (
            .O(N__43357),
            .I(N__43318));
    InMux I__10831 (
            .O(N__43356),
            .I(N__43311));
    InMux I__10830 (
            .O(N__43355),
            .I(N__43311));
    InMux I__10829 (
            .O(N__43354),
            .I(N__43311));
    LocalMux I__10828 (
            .O(N__43351),
            .I(N__43306));
    Span4Mux_h I__10827 (
            .O(N__43344),
            .I(N__43306));
    Odrv4 I__10826 (
            .O(N__43341),
            .I(N_765_0));
    Odrv4 I__10825 (
            .O(N__43338),
            .I(N_765_0));
    Odrv4 I__10824 (
            .O(N__43335),
            .I(N_765_0));
    LocalMux I__10823 (
            .O(N__43332),
            .I(N_765_0));
    LocalMux I__10822 (
            .O(N__43329),
            .I(N_765_0));
    Odrv4 I__10821 (
            .O(N__43326),
            .I(N_765_0));
    LocalMux I__10820 (
            .O(N__43323),
            .I(N_765_0));
    Odrv4 I__10819 (
            .O(N__43318),
            .I(N_765_0));
    LocalMux I__10818 (
            .O(N__43311),
            .I(N_765_0));
    Odrv4 I__10817 (
            .O(N__43306),
            .I(N_765_0));
    InMux I__10816 (
            .O(N__43285),
            .I(N__43282));
    LocalMux I__10815 (
            .O(N__43282),
            .I(un1_M_this_ext_address_q_cry_5_THRU_CO));
    IoInMux I__10814 (
            .O(N__43279),
            .I(N__43276));
    LocalMux I__10813 (
            .O(N__43276),
            .I(N__43272));
    CascadeMux I__10812 (
            .O(N__43275),
            .I(N__43268));
    Span12Mux_s5_h I__10811 (
            .O(N__43272),
            .I(N__43265));
    InMux I__10810 (
            .O(N__43271),
            .I(N__43262));
    InMux I__10809 (
            .O(N__43268),
            .I(N__43259));
    Odrv12 I__10808 (
            .O(N__43265),
            .I(M_this_ext_address_qZ0Z_6));
    LocalMux I__10807 (
            .O(N__43262),
            .I(M_this_ext_address_qZ0Z_6));
    LocalMux I__10806 (
            .O(N__43259),
            .I(M_this_ext_address_qZ0Z_6));
    CascadeMux I__10805 (
            .O(N__43252),
            .I(N__43245));
    CascadeMux I__10804 (
            .O(N__43251),
            .I(N__43229));
    InMux I__10803 (
            .O(N__43250),
            .I(N__43212));
    InMux I__10802 (
            .O(N__43249),
            .I(N__43212));
    InMux I__10801 (
            .O(N__43248),
            .I(N__43209));
    InMux I__10800 (
            .O(N__43245),
            .I(N__43206));
    InMux I__10799 (
            .O(N__43244),
            .I(N__43203));
    InMux I__10798 (
            .O(N__43243),
            .I(N__43200));
    InMux I__10797 (
            .O(N__43242),
            .I(N__43197));
    InMux I__10796 (
            .O(N__43241),
            .I(N__43194));
    InMux I__10795 (
            .O(N__43240),
            .I(N__43191));
    InMux I__10794 (
            .O(N__43239),
            .I(N__43186));
    InMux I__10793 (
            .O(N__43238),
            .I(N__43186));
    InMux I__10792 (
            .O(N__43237),
            .I(N__43183));
    InMux I__10791 (
            .O(N__43236),
            .I(N__43180));
    InMux I__10790 (
            .O(N__43235),
            .I(N__43177));
    InMux I__10789 (
            .O(N__43234),
            .I(N__43174));
    InMux I__10788 (
            .O(N__43233),
            .I(N__43171));
    InMux I__10787 (
            .O(N__43232),
            .I(N__43166));
    InMux I__10786 (
            .O(N__43229),
            .I(N__43166));
    InMux I__10785 (
            .O(N__43228),
            .I(N__43163));
    InMux I__10784 (
            .O(N__43227),
            .I(N__43158));
    InMux I__10783 (
            .O(N__43226),
            .I(N__43158));
    InMux I__10782 (
            .O(N__43225),
            .I(N__43153));
    InMux I__10781 (
            .O(N__43224),
            .I(N__43153));
    InMux I__10780 (
            .O(N__43223),
            .I(N__43150));
    InMux I__10779 (
            .O(N__43222),
            .I(N__43147));
    InMux I__10778 (
            .O(N__43221),
            .I(N__43144));
    InMux I__10777 (
            .O(N__43220),
            .I(N__43141));
    InMux I__10776 (
            .O(N__43219),
            .I(N__43138));
    InMux I__10775 (
            .O(N__43218),
            .I(N__43135));
    InMux I__10774 (
            .O(N__43217),
            .I(N__43132));
    LocalMux I__10773 (
            .O(N__43212),
            .I(N__43094));
    LocalMux I__10772 (
            .O(N__43209),
            .I(N__43091));
    LocalMux I__10771 (
            .O(N__43206),
            .I(N__43088));
    LocalMux I__10770 (
            .O(N__43203),
            .I(N__43085));
    LocalMux I__10769 (
            .O(N__43200),
            .I(N__43082));
    LocalMux I__10768 (
            .O(N__43197),
            .I(N__43079));
    LocalMux I__10767 (
            .O(N__43194),
            .I(N__43076));
    LocalMux I__10766 (
            .O(N__43191),
            .I(N__43073));
    LocalMux I__10765 (
            .O(N__43186),
            .I(N__43070));
    LocalMux I__10764 (
            .O(N__43183),
            .I(N__43067));
    LocalMux I__10763 (
            .O(N__43180),
            .I(N__43064));
    LocalMux I__10762 (
            .O(N__43177),
            .I(N__43061));
    LocalMux I__10761 (
            .O(N__43174),
            .I(N__43058));
    LocalMux I__10760 (
            .O(N__43171),
            .I(N__43055));
    LocalMux I__10759 (
            .O(N__43166),
            .I(N__43052));
    LocalMux I__10758 (
            .O(N__43163),
            .I(N__43049));
    LocalMux I__10757 (
            .O(N__43158),
            .I(N__43046));
    LocalMux I__10756 (
            .O(N__43153),
            .I(N__43043));
    LocalMux I__10755 (
            .O(N__43150),
            .I(N__43040));
    LocalMux I__10754 (
            .O(N__43147),
            .I(N__43037));
    LocalMux I__10753 (
            .O(N__43144),
            .I(N__43034));
    LocalMux I__10752 (
            .O(N__43141),
            .I(N__43031));
    LocalMux I__10751 (
            .O(N__43138),
            .I(N__43028));
    LocalMux I__10750 (
            .O(N__43135),
            .I(N__43025));
    LocalMux I__10749 (
            .O(N__43132),
            .I(N__43022));
    SRMux I__10748 (
            .O(N__43131),
            .I(N__42901));
    SRMux I__10747 (
            .O(N__43130),
            .I(N__42901));
    SRMux I__10746 (
            .O(N__43129),
            .I(N__42901));
    SRMux I__10745 (
            .O(N__43128),
            .I(N__42901));
    SRMux I__10744 (
            .O(N__43127),
            .I(N__42901));
    SRMux I__10743 (
            .O(N__43126),
            .I(N__42901));
    SRMux I__10742 (
            .O(N__43125),
            .I(N__42901));
    SRMux I__10741 (
            .O(N__43124),
            .I(N__42901));
    SRMux I__10740 (
            .O(N__43123),
            .I(N__42901));
    SRMux I__10739 (
            .O(N__43122),
            .I(N__42901));
    SRMux I__10738 (
            .O(N__43121),
            .I(N__42901));
    SRMux I__10737 (
            .O(N__43120),
            .I(N__42901));
    SRMux I__10736 (
            .O(N__43119),
            .I(N__42901));
    SRMux I__10735 (
            .O(N__43118),
            .I(N__42901));
    SRMux I__10734 (
            .O(N__43117),
            .I(N__42901));
    SRMux I__10733 (
            .O(N__43116),
            .I(N__42901));
    SRMux I__10732 (
            .O(N__43115),
            .I(N__42901));
    SRMux I__10731 (
            .O(N__43114),
            .I(N__42901));
    SRMux I__10730 (
            .O(N__43113),
            .I(N__42901));
    SRMux I__10729 (
            .O(N__43112),
            .I(N__42901));
    SRMux I__10728 (
            .O(N__43111),
            .I(N__42901));
    SRMux I__10727 (
            .O(N__43110),
            .I(N__42901));
    SRMux I__10726 (
            .O(N__43109),
            .I(N__42901));
    SRMux I__10725 (
            .O(N__43108),
            .I(N__42901));
    SRMux I__10724 (
            .O(N__43107),
            .I(N__42901));
    SRMux I__10723 (
            .O(N__43106),
            .I(N__42901));
    SRMux I__10722 (
            .O(N__43105),
            .I(N__42901));
    SRMux I__10721 (
            .O(N__43104),
            .I(N__42901));
    SRMux I__10720 (
            .O(N__43103),
            .I(N__42901));
    SRMux I__10719 (
            .O(N__43102),
            .I(N__42901));
    SRMux I__10718 (
            .O(N__43101),
            .I(N__42901));
    SRMux I__10717 (
            .O(N__43100),
            .I(N__42901));
    SRMux I__10716 (
            .O(N__43099),
            .I(N__42901));
    SRMux I__10715 (
            .O(N__43098),
            .I(N__42901));
    SRMux I__10714 (
            .O(N__43097),
            .I(N__42901));
    Glb2LocalMux I__10713 (
            .O(N__43094),
            .I(N__42901));
    Glb2LocalMux I__10712 (
            .O(N__43091),
            .I(N__42901));
    Glb2LocalMux I__10711 (
            .O(N__43088),
            .I(N__42901));
    Glb2LocalMux I__10710 (
            .O(N__43085),
            .I(N__42901));
    Glb2LocalMux I__10709 (
            .O(N__43082),
            .I(N__42901));
    Glb2LocalMux I__10708 (
            .O(N__43079),
            .I(N__42901));
    Glb2LocalMux I__10707 (
            .O(N__43076),
            .I(N__42901));
    Glb2LocalMux I__10706 (
            .O(N__43073),
            .I(N__42901));
    Glb2LocalMux I__10705 (
            .O(N__43070),
            .I(N__42901));
    Glb2LocalMux I__10704 (
            .O(N__43067),
            .I(N__42901));
    Glb2LocalMux I__10703 (
            .O(N__43064),
            .I(N__42901));
    Glb2LocalMux I__10702 (
            .O(N__43061),
            .I(N__42901));
    Glb2LocalMux I__10701 (
            .O(N__43058),
            .I(N__42901));
    Glb2LocalMux I__10700 (
            .O(N__43055),
            .I(N__42901));
    Glb2LocalMux I__10699 (
            .O(N__43052),
            .I(N__42901));
    Glb2LocalMux I__10698 (
            .O(N__43049),
            .I(N__42901));
    Glb2LocalMux I__10697 (
            .O(N__43046),
            .I(N__42901));
    Glb2LocalMux I__10696 (
            .O(N__43043),
            .I(N__42901));
    Glb2LocalMux I__10695 (
            .O(N__43040),
            .I(N__42901));
    Glb2LocalMux I__10694 (
            .O(N__43037),
            .I(N__42901));
    Glb2LocalMux I__10693 (
            .O(N__43034),
            .I(N__42901));
    Glb2LocalMux I__10692 (
            .O(N__43031),
            .I(N__42901));
    Glb2LocalMux I__10691 (
            .O(N__43028),
            .I(N__42901));
    Glb2LocalMux I__10690 (
            .O(N__43025),
            .I(N__42901));
    Glb2LocalMux I__10689 (
            .O(N__43022),
            .I(N__42901));
    GlobalMux I__10688 (
            .O(N__42901),
            .I(N__42898));
    gio2CtrlBuf I__10687 (
            .O(N__42898),
            .I(M_this_reset_cond_out_g_0));
    InMux I__10686 (
            .O(N__42895),
            .I(N__42892));
    LocalMux I__10685 (
            .O(N__42892),
            .I(N__42889));
    Odrv12 I__10684 (
            .O(N__42889),
            .I(un1_M_this_map_address_q_cry_6_THRU_CO));
    CascadeMux I__10683 (
            .O(N__42886),
            .I(N__42883));
    CascadeBuf I__10682 (
            .O(N__42883),
            .I(N__42880));
    CascadeMux I__10681 (
            .O(N__42880),
            .I(N__42877));
    InMux I__10680 (
            .O(N__42877),
            .I(N__42874));
    LocalMux I__10679 (
            .O(N__42874),
            .I(N__42871));
    Span4Mux_h I__10678 (
            .O(N__42871),
            .I(N__42866));
    CascadeMux I__10677 (
            .O(N__42870),
            .I(N__42863));
    InMux I__10676 (
            .O(N__42869),
            .I(N__42860));
    Span4Mux_v I__10675 (
            .O(N__42866),
            .I(N__42856));
    InMux I__10674 (
            .O(N__42863),
            .I(N__42853));
    LocalMux I__10673 (
            .O(N__42860),
            .I(N__42850));
    InMux I__10672 (
            .O(N__42859),
            .I(N__42847));
    Span4Mux_v I__10671 (
            .O(N__42856),
            .I(N__42844));
    LocalMux I__10670 (
            .O(N__42853),
            .I(M_this_map_address_qZ0Z_7));
    Odrv4 I__10669 (
            .O(N__42850),
            .I(M_this_map_address_qZ0Z_7));
    LocalMux I__10668 (
            .O(N__42847),
            .I(M_this_map_address_qZ0Z_7));
    Odrv4 I__10667 (
            .O(N__42844),
            .I(M_this_map_address_qZ0Z_7));
    InMux I__10666 (
            .O(N__42835),
            .I(N__42831));
    InMux I__10665 (
            .O(N__42834),
            .I(N__42825));
    LocalMux I__10664 (
            .O(N__42831),
            .I(N__42822));
    InMux I__10663 (
            .O(N__42830),
            .I(N__42817));
    InMux I__10662 (
            .O(N__42829),
            .I(N__42817));
    InMux I__10661 (
            .O(N__42828),
            .I(N__42814));
    LocalMux I__10660 (
            .O(N__42825),
            .I(N__42807));
    Span4Mux_v I__10659 (
            .O(N__42822),
            .I(N__42807));
    LocalMux I__10658 (
            .O(N__42817),
            .I(N__42807));
    LocalMux I__10657 (
            .O(N__42814),
            .I(N__42804));
    Span4Mux_h I__10656 (
            .O(N__42807),
            .I(N__42801));
    Odrv12 I__10655 (
            .O(N__42804),
            .I(N_801_0));
    Odrv4 I__10654 (
            .O(N__42801),
            .I(N_801_0));
    InMux I__10653 (
            .O(N__42796),
            .I(N__42793));
    LocalMux I__10652 (
            .O(N__42793),
            .I(N__42788));
    InMux I__10651 (
            .O(N__42792),
            .I(N__42785));
    InMux I__10650 (
            .O(N__42791),
            .I(N__42782));
    Span4Mux_h I__10649 (
            .O(N__42788),
            .I(N__42775));
    LocalMux I__10648 (
            .O(N__42785),
            .I(N__42775));
    LocalMux I__10647 (
            .O(N__42782),
            .I(N__42775));
    Span4Mux_v I__10646 (
            .O(N__42775),
            .I(N__42769));
    InMux I__10645 (
            .O(N__42774),
            .I(N__42766));
    InMux I__10644 (
            .O(N__42773),
            .I(N__42761));
    InMux I__10643 (
            .O(N__42772),
            .I(N__42758));
    Span4Mux_h I__10642 (
            .O(N__42769),
            .I(N__42754));
    LocalMux I__10641 (
            .O(N__42766),
            .I(N__42751));
    InMux I__10640 (
            .O(N__42765),
            .I(N__42747));
    InMux I__10639 (
            .O(N__42764),
            .I(N__42744));
    LocalMux I__10638 (
            .O(N__42761),
            .I(N__42741));
    LocalMux I__10637 (
            .O(N__42758),
            .I(N__42738));
    CascadeMux I__10636 (
            .O(N__42757),
            .I(N__42735));
    Span4Mux_h I__10635 (
            .O(N__42754),
            .I(N__42732));
    Span4Mux_v I__10634 (
            .O(N__42751),
            .I(N__42729));
    InMux I__10633 (
            .O(N__42750),
            .I(N__42726));
    LocalMux I__10632 (
            .O(N__42747),
            .I(N__42723));
    LocalMux I__10631 (
            .O(N__42744),
            .I(N__42720));
    Span4Mux_v I__10630 (
            .O(N__42741),
            .I(N__42717));
    Span4Mux_v I__10629 (
            .O(N__42738),
            .I(N__42714));
    InMux I__10628 (
            .O(N__42735),
            .I(N__42711));
    Span4Mux_h I__10627 (
            .O(N__42732),
            .I(N__42703));
    Span4Mux_v I__10626 (
            .O(N__42729),
            .I(N__42703));
    LocalMux I__10625 (
            .O(N__42726),
            .I(N__42703));
    Span12Mux_v I__10624 (
            .O(N__42723),
            .I(N__42698));
    Span12Mux_h I__10623 (
            .O(N__42720),
            .I(N__42698));
    IoSpan4Mux I__10622 (
            .O(N__42717),
            .I(N__42695));
    Sp12to4 I__10621 (
            .O(N__42714),
            .I(N__42692));
    LocalMux I__10620 (
            .O(N__42711),
            .I(N__42689));
    InMux I__10619 (
            .O(N__42710),
            .I(N__42686));
    Span4Mux_h I__10618 (
            .O(N__42703),
            .I(N__42683));
    Span12Mux_h I__10617 (
            .O(N__42698),
            .I(N__42680));
    IoSpan4Mux I__10616 (
            .O(N__42695),
            .I(N__42677));
    Span12Mux_h I__10615 (
            .O(N__42692),
            .I(N__42670));
    Sp12to4 I__10614 (
            .O(N__42689),
            .I(N__42670));
    LocalMux I__10613 (
            .O(N__42686),
            .I(N__42670));
    Span4Mux_v I__10612 (
            .O(N__42683),
            .I(N__42667));
    Odrv12 I__10611 (
            .O(N__42680),
            .I(port_data_in_2));
    Odrv4 I__10610 (
            .O(N__42677),
            .I(port_data_in_2));
    Odrv12 I__10609 (
            .O(N__42670),
            .I(port_data_in_2));
    Odrv4 I__10608 (
            .O(N__42667),
            .I(port_data_in_2));
    CascadeMux I__10607 (
            .O(N__42658),
            .I(N_1075_cascade_));
    InMux I__10606 (
            .O(N__42655),
            .I(N__42652));
    LocalMux I__10605 (
            .O(N__42652),
            .I(M_this_map_address_qc_1_0));
    InMux I__10604 (
            .O(N__42649),
            .I(N__42645));
    InMux I__10603 (
            .O(N__42648),
            .I(N__42642));
    LocalMux I__10602 (
            .O(N__42645),
            .I(N__42637));
    LocalMux I__10601 (
            .O(N__42642),
            .I(N__42637));
    Span4Mux_v I__10600 (
            .O(N__42637),
            .I(N__42633));
    InMux I__10599 (
            .O(N__42636),
            .I(N__42630));
    Span4Mux_h I__10598 (
            .O(N__42633),
            .I(N__42625));
    LocalMux I__10597 (
            .O(N__42630),
            .I(N__42625));
    Span4Mux_h I__10596 (
            .O(N__42625),
            .I(N__42622));
    Span4Mux_v I__10595 (
            .O(N__42622),
            .I(N__42619));
    Odrv4 I__10594 (
            .O(N__42619),
            .I(port_address_in_3));
    InMux I__10593 (
            .O(N__42616),
            .I(N__42611));
    InMux I__10592 (
            .O(N__42615),
            .I(N__42608));
    InMux I__10591 (
            .O(N__42614),
            .I(N__42605));
    LocalMux I__10590 (
            .O(N__42611),
            .I(N__42598));
    LocalMux I__10589 (
            .O(N__42608),
            .I(N__42598));
    LocalMux I__10588 (
            .O(N__42605),
            .I(N__42598));
    Odrv12 I__10587 (
            .O(N__42598),
            .I(N_459_0));
    InMux I__10586 (
            .O(N__42595),
            .I(N__42589));
    InMux I__10585 (
            .O(N__42594),
            .I(N__42585));
    InMux I__10584 (
            .O(N__42593),
            .I(N__42582));
    InMux I__10583 (
            .O(N__42592),
            .I(N__42579));
    LocalMux I__10582 (
            .O(N__42589),
            .I(N__42576));
    InMux I__10581 (
            .O(N__42588),
            .I(N__42573));
    LocalMux I__10580 (
            .O(N__42585),
            .I(N__42568));
    LocalMux I__10579 (
            .O(N__42582),
            .I(N__42568));
    LocalMux I__10578 (
            .O(N__42579),
            .I(N__42565));
    Span4Mux_h I__10577 (
            .O(N__42576),
            .I(N__42562));
    LocalMux I__10576 (
            .O(N__42573),
            .I(N__42555));
    Span4Mux_v I__10575 (
            .O(N__42568),
            .I(N__42555));
    Span4Mux_h I__10574 (
            .O(N__42565),
            .I(N__42555));
    Span4Mux_h I__10573 (
            .O(N__42562),
            .I(N__42552));
    Span4Mux_h I__10572 (
            .O(N__42555),
            .I(N__42549));
    Odrv4 I__10571 (
            .O(N__42552),
            .I(N_1276));
    Odrv4 I__10570 (
            .O(N__42549),
            .I(N_1276));
    InMux I__10569 (
            .O(N__42544),
            .I(N__42536));
    InMux I__10568 (
            .O(N__42543),
            .I(N__42533));
    CascadeMux I__10567 (
            .O(N__42542),
            .I(N__42530));
    InMux I__10566 (
            .O(N__42541),
            .I(N__42526));
    InMux I__10565 (
            .O(N__42540),
            .I(N__42523));
    InMux I__10564 (
            .O(N__42539),
            .I(N__42520));
    LocalMux I__10563 (
            .O(N__42536),
            .I(N__42517));
    LocalMux I__10562 (
            .O(N__42533),
            .I(N__42514));
    InMux I__10561 (
            .O(N__42530),
            .I(N__42509));
    InMux I__10560 (
            .O(N__42529),
            .I(N__42509));
    LocalMux I__10559 (
            .O(N__42526),
            .I(N__42500));
    LocalMux I__10558 (
            .O(N__42523),
            .I(N__42500));
    LocalMux I__10557 (
            .O(N__42520),
            .I(N__42500));
    Span12Mux_v I__10556 (
            .O(N__42517),
            .I(N__42496));
    Span4Mux_v I__10555 (
            .O(N__42514),
            .I(N__42493));
    LocalMux I__10554 (
            .O(N__42509),
            .I(N__42490));
    InMux I__10553 (
            .O(N__42508),
            .I(N__42487));
    InMux I__10552 (
            .O(N__42507),
            .I(N__42484));
    Span12Mux_s10_h I__10551 (
            .O(N__42500),
            .I(N__42481));
    InMux I__10550 (
            .O(N__42499),
            .I(N__42478));
    Odrv12 I__10549 (
            .O(N__42496),
            .I(N_1242));
    Odrv4 I__10548 (
            .O(N__42493),
            .I(N_1242));
    Odrv4 I__10547 (
            .O(N__42490),
            .I(N_1242));
    LocalMux I__10546 (
            .O(N__42487),
            .I(N_1242));
    LocalMux I__10545 (
            .O(N__42484),
            .I(N_1242));
    Odrv12 I__10544 (
            .O(N__42481),
            .I(N_1242));
    LocalMux I__10543 (
            .O(N__42478),
            .I(N_1242));
    CascadeMux I__10542 (
            .O(N__42463),
            .I(N__42460));
    InMux I__10541 (
            .O(N__42460),
            .I(N__42456));
    CascadeMux I__10540 (
            .O(N__42459),
            .I(N__42453));
    LocalMux I__10539 (
            .O(N__42456),
            .I(N__42450));
    InMux I__10538 (
            .O(N__42453),
            .I(N__42446));
    Span4Mux_h I__10537 (
            .O(N__42450),
            .I(N__42440));
    InMux I__10536 (
            .O(N__42449),
            .I(N__42436));
    LocalMux I__10535 (
            .O(N__42446),
            .I(N__42433));
    InMux I__10534 (
            .O(N__42445),
            .I(N__42430));
    InMux I__10533 (
            .O(N__42444),
            .I(N__42426));
    InMux I__10532 (
            .O(N__42443),
            .I(N__42423));
    Span4Mux_h I__10531 (
            .O(N__42440),
            .I(N__42420));
    InMux I__10530 (
            .O(N__42439),
            .I(N__42417));
    LocalMux I__10529 (
            .O(N__42436),
            .I(N__42412));
    Span4Mux_h I__10528 (
            .O(N__42433),
            .I(N__42407));
    LocalMux I__10527 (
            .O(N__42430),
            .I(N__42407));
    InMux I__10526 (
            .O(N__42429),
            .I(N__42404));
    LocalMux I__10525 (
            .O(N__42426),
            .I(N__42401));
    LocalMux I__10524 (
            .O(N__42423),
            .I(N__42398));
    Span4Mux_h I__10523 (
            .O(N__42420),
            .I(N__42393));
    LocalMux I__10522 (
            .O(N__42417),
            .I(N__42393));
    InMux I__10521 (
            .O(N__42416),
            .I(N__42390));
    InMux I__10520 (
            .O(N__42415),
            .I(N__42387));
    Span4Mux_v I__10519 (
            .O(N__42412),
            .I(N__42384));
    Span4Mux_h I__10518 (
            .O(N__42407),
            .I(N__42381));
    LocalMux I__10517 (
            .O(N__42404),
            .I(N__42378));
    Span4Mux_h I__10516 (
            .O(N__42401),
            .I(N__42374));
    Span4Mux_v I__10515 (
            .O(N__42398),
            .I(N__42371));
    Span4Mux_h I__10514 (
            .O(N__42393),
            .I(N__42368));
    LocalMux I__10513 (
            .O(N__42390),
            .I(N__42363));
    LocalMux I__10512 (
            .O(N__42387),
            .I(N__42363));
    Span4Mux_v I__10511 (
            .O(N__42384),
            .I(N__42358));
    Span4Mux_h I__10510 (
            .O(N__42381),
            .I(N__42358));
    Span4Mux_v I__10509 (
            .O(N__42378),
            .I(N__42355));
    InMux I__10508 (
            .O(N__42377),
            .I(N__42352));
    Span4Mux_v I__10507 (
            .O(N__42374),
            .I(N__42347));
    Span4Mux_h I__10506 (
            .O(N__42371),
            .I(N__42347));
    Span4Mux_v I__10505 (
            .O(N__42368),
            .I(N__42342));
    Span4Mux_h I__10504 (
            .O(N__42363),
            .I(N__42342));
    Span4Mux_h I__10503 (
            .O(N__42358),
            .I(N__42339));
    Sp12to4 I__10502 (
            .O(N__42355),
            .I(N__42334));
    LocalMux I__10501 (
            .O(N__42352),
            .I(N__42334));
    Span4Mux_h I__10500 (
            .O(N__42347),
            .I(N__42329));
    Span4Mux_v I__10499 (
            .O(N__42342),
            .I(N__42329));
    Sp12to4 I__10498 (
            .O(N__42339),
            .I(N__42324));
    Span12Mux_h I__10497 (
            .O(N__42334),
            .I(N__42324));
    Odrv4 I__10496 (
            .O(N__42329),
            .I(port_data_in_0));
    Odrv12 I__10495 (
            .O(N__42324),
            .I(port_data_in_0));
    InMux I__10494 (
            .O(N__42319),
            .I(N__42316));
    LocalMux I__10493 (
            .O(N__42316),
            .I(N_1068));
    InMux I__10492 (
            .O(N__42313),
            .I(N__42310));
    LocalMux I__10491 (
            .O(N__42310),
            .I(M_this_map_address_qc_7_1));
    InMux I__10490 (
            .O(N__42307),
            .I(N__42304));
    LocalMux I__10489 (
            .O(N__42304),
            .I(N__42301));
    Span4Mux_h I__10488 (
            .O(N__42301),
            .I(N__42298));
    Odrv4 I__10487 (
            .O(N__42298),
            .I(M_this_map_address_q_RNO_1Z0Z_5));
    CascadeMux I__10486 (
            .O(N__42295),
            .I(N__42290));
    InMux I__10485 (
            .O(N__42294),
            .I(N__42285));
    InMux I__10484 (
            .O(N__42293),
            .I(N__42280));
    InMux I__10483 (
            .O(N__42290),
            .I(N__42277));
    InMux I__10482 (
            .O(N__42289),
            .I(N__42274));
    InMux I__10481 (
            .O(N__42288),
            .I(N__42271));
    LocalMux I__10480 (
            .O(N__42285),
            .I(N__42268));
    InMux I__10479 (
            .O(N__42284),
            .I(N__42263));
    InMux I__10478 (
            .O(N__42283),
            .I(N__42263));
    LocalMux I__10477 (
            .O(N__42280),
            .I(N__42255));
    LocalMux I__10476 (
            .O(N__42277),
            .I(N__42250));
    LocalMux I__10475 (
            .O(N__42274),
            .I(N__42250));
    LocalMux I__10474 (
            .O(N__42271),
            .I(N__42247));
    Span4Mux_v I__10473 (
            .O(N__42268),
            .I(N__42244));
    LocalMux I__10472 (
            .O(N__42263),
            .I(N__42241));
    InMux I__10471 (
            .O(N__42262),
            .I(N__42237));
    CascadeMux I__10470 (
            .O(N__42261),
            .I(N__42234));
    InMux I__10469 (
            .O(N__42260),
            .I(N__42227));
    InMux I__10468 (
            .O(N__42259),
            .I(N__42227));
    InMux I__10467 (
            .O(N__42258),
            .I(N__42227));
    Span4Mux_h I__10466 (
            .O(N__42255),
            .I(N__42220));
    Span4Mux_v I__10465 (
            .O(N__42250),
            .I(N__42220));
    Span4Mux_v I__10464 (
            .O(N__42247),
            .I(N__42220));
    Span4Mux_h I__10463 (
            .O(N__42244),
            .I(N__42217));
    Span4Mux_h I__10462 (
            .O(N__42241),
            .I(N__42214));
    InMux I__10461 (
            .O(N__42240),
            .I(N__42211));
    LocalMux I__10460 (
            .O(N__42237),
            .I(N__42208));
    InMux I__10459 (
            .O(N__42234),
            .I(N__42205));
    LocalMux I__10458 (
            .O(N__42227),
            .I(N_1258));
    Odrv4 I__10457 (
            .O(N__42220),
            .I(N_1258));
    Odrv4 I__10456 (
            .O(N__42217),
            .I(N_1258));
    Odrv4 I__10455 (
            .O(N__42214),
            .I(N_1258));
    LocalMux I__10454 (
            .O(N__42211),
            .I(N_1258));
    Odrv12 I__10453 (
            .O(N__42208),
            .I(N_1258));
    LocalMux I__10452 (
            .O(N__42205),
            .I(N_1258));
    CascadeMux I__10451 (
            .O(N__42190),
            .I(N__42187));
    CascadeBuf I__10450 (
            .O(N__42187),
            .I(N__42184));
    CascadeMux I__10449 (
            .O(N__42184),
            .I(N__42180));
    CascadeMux I__10448 (
            .O(N__42183),
            .I(N__42177));
    InMux I__10447 (
            .O(N__42180),
            .I(N__42174));
    InMux I__10446 (
            .O(N__42177),
            .I(N__42171));
    LocalMux I__10445 (
            .O(N__42174),
            .I(N__42168));
    LocalMux I__10444 (
            .O(N__42171),
            .I(N__42164));
    Span4Mux_s2_v I__10443 (
            .O(N__42168),
            .I(N__42161));
    InMux I__10442 (
            .O(N__42167),
            .I(N__42158));
    Span4Mux_h I__10441 (
            .O(N__42164),
            .I(N__42155));
    Span4Mux_v I__10440 (
            .O(N__42161),
            .I(N__42152));
    LocalMux I__10439 (
            .O(N__42158),
            .I(M_this_map_address_qZ0Z_5));
    Odrv4 I__10438 (
            .O(N__42155),
            .I(M_this_map_address_qZ0Z_5));
    Odrv4 I__10437 (
            .O(N__42152),
            .I(M_this_map_address_qZ0Z_5));
    ClkMux I__10436 (
            .O(N__42145),
            .I(N__41659));
    ClkMux I__10435 (
            .O(N__42144),
            .I(N__41659));
    ClkMux I__10434 (
            .O(N__42143),
            .I(N__41659));
    ClkMux I__10433 (
            .O(N__42142),
            .I(N__41659));
    ClkMux I__10432 (
            .O(N__42141),
            .I(N__41659));
    ClkMux I__10431 (
            .O(N__42140),
            .I(N__41659));
    ClkMux I__10430 (
            .O(N__42139),
            .I(N__41659));
    ClkMux I__10429 (
            .O(N__42138),
            .I(N__41659));
    ClkMux I__10428 (
            .O(N__42137),
            .I(N__41659));
    ClkMux I__10427 (
            .O(N__42136),
            .I(N__41659));
    ClkMux I__10426 (
            .O(N__42135),
            .I(N__41659));
    ClkMux I__10425 (
            .O(N__42134),
            .I(N__41659));
    ClkMux I__10424 (
            .O(N__42133),
            .I(N__41659));
    ClkMux I__10423 (
            .O(N__42132),
            .I(N__41659));
    ClkMux I__10422 (
            .O(N__42131),
            .I(N__41659));
    ClkMux I__10421 (
            .O(N__42130),
            .I(N__41659));
    ClkMux I__10420 (
            .O(N__42129),
            .I(N__41659));
    ClkMux I__10419 (
            .O(N__42128),
            .I(N__41659));
    ClkMux I__10418 (
            .O(N__42127),
            .I(N__41659));
    ClkMux I__10417 (
            .O(N__42126),
            .I(N__41659));
    ClkMux I__10416 (
            .O(N__42125),
            .I(N__41659));
    ClkMux I__10415 (
            .O(N__42124),
            .I(N__41659));
    ClkMux I__10414 (
            .O(N__42123),
            .I(N__41659));
    ClkMux I__10413 (
            .O(N__42122),
            .I(N__41659));
    ClkMux I__10412 (
            .O(N__42121),
            .I(N__41659));
    ClkMux I__10411 (
            .O(N__42120),
            .I(N__41659));
    ClkMux I__10410 (
            .O(N__42119),
            .I(N__41659));
    ClkMux I__10409 (
            .O(N__42118),
            .I(N__41659));
    ClkMux I__10408 (
            .O(N__42117),
            .I(N__41659));
    ClkMux I__10407 (
            .O(N__42116),
            .I(N__41659));
    ClkMux I__10406 (
            .O(N__42115),
            .I(N__41659));
    ClkMux I__10405 (
            .O(N__42114),
            .I(N__41659));
    ClkMux I__10404 (
            .O(N__42113),
            .I(N__41659));
    ClkMux I__10403 (
            .O(N__42112),
            .I(N__41659));
    ClkMux I__10402 (
            .O(N__42111),
            .I(N__41659));
    ClkMux I__10401 (
            .O(N__42110),
            .I(N__41659));
    ClkMux I__10400 (
            .O(N__42109),
            .I(N__41659));
    ClkMux I__10399 (
            .O(N__42108),
            .I(N__41659));
    ClkMux I__10398 (
            .O(N__42107),
            .I(N__41659));
    ClkMux I__10397 (
            .O(N__42106),
            .I(N__41659));
    ClkMux I__10396 (
            .O(N__42105),
            .I(N__41659));
    ClkMux I__10395 (
            .O(N__42104),
            .I(N__41659));
    ClkMux I__10394 (
            .O(N__42103),
            .I(N__41659));
    ClkMux I__10393 (
            .O(N__42102),
            .I(N__41659));
    ClkMux I__10392 (
            .O(N__42101),
            .I(N__41659));
    ClkMux I__10391 (
            .O(N__42100),
            .I(N__41659));
    ClkMux I__10390 (
            .O(N__42099),
            .I(N__41659));
    ClkMux I__10389 (
            .O(N__42098),
            .I(N__41659));
    ClkMux I__10388 (
            .O(N__42097),
            .I(N__41659));
    ClkMux I__10387 (
            .O(N__42096),
            .I(N__41659));
    ClkMux I__10386 (
            .O(N__42095),
            .I(N__41659));
    ClkMux I__10385 (
            .O(N__42094),
            .I(N__41659));
    ClkMux I__10384 (
            .O(N__42093),
            .I(N__41659));
    ClkMux I__10383 (
            .O(N__42092),
            .I(N__41659));
    ClkMux I__10382 (
            .O(N__42091),
            .I(N__41659));
    ClkMux I__10381 (
            .O(N__42090),
            .I(N__41659));
    ClkMux I__10380 (
            .O(N__42089),
            .I(N__41659));
    ClkMux I__10379 (
            .O(N__42088),
            .I(N__41659));
    ClkMux I__10378 (
            .O(N__42087),
            .I(N__41659));
    ClkMux I__10377 (
            .O(N__42086),
            .I(N__41659));
    ClkMux I__10376 (
            .O(N__42085),
            .I(N__41659));
    ClkMux I__10375 (
            .O(N__42084),
            .I(N__41659));
    ClkMux I__10374 (
            .O(N__42083),
            .I(N__41659));
    ClkMux I__10373 (
            .O(N__42082),
            .I(N__41659));
    ClkMux I__10372 (
            .O(N__42081),
            .I(N__41659));
    ClkMux I__10371 (
            .O(N__42080),
            .I(N__41659));
    ClkMux I__10370 (
            .O(N__42079),
            .I(N__41659));
    ClkMux I__10369 (
            .O(N__42078),
            .I(N__41659));
    ClkMux I__10368 (
            .O(N__42077),
            .I(N__41659));
    ClkMux I__10367 (
            .O(N__42076),
            .I(N__41659));
    ClkMux I__10366 (
            .O(N__42075),
            .I(N__41659));
    ClkMux I__10365 (
            .O(N__42074),
            .I(N__41659));
    ClkMux I__10364 (
            .O(N__42073),
            .I(N__41659));
    ClkMux I__10363 (
            .O(N__42072),
            .I(N__41659));
    ClkMux I__10362 (
            .O(N__42071),
            .I(N__41659));
    ClkMux I__10361 (
            .O(N__42070),
            .I(N__41659));
    ClkMux I__10360 (
            .O(N__42069),
            .I(N__41659));
    ClkMux I__10359 (
            .O(N__42068),
            .I(N__41659));
    ClkMux I__10358 (
            .O(N__42067),
            .I(N__41659));
    ClkMux I__10357 (
            .O(N__42066),
            .I(N__41659));
    ClkMux I__10356 (
            .O(N__42065),
            .I(N__41659));
    ClkMux I__10355 (
            .O(N__42064),
            .I(N__41659));
    ClkMux I__10354 (
            .O(N__42063),
            .I(N__41659));
    ClkMux I__10353 (
            .O(N__42062),
            .I(N__41659));
    ClkMux I__10352 (
            .O(N__42061),
            .I(N__41659));
    ClkMux I__10351 (
            .O(N__42060),
            .I(N__41659));
    ClkMux I__10350 (
            .O(N__42059),
            .I(N__41659));
    ClkMux I__10349 (
            .O(N__42058),
            .I(N__41659));
    ClkMux I__10348 (
            .O(N__42057),
            .I(N__41659));
    ClkMux I__10347 (
            .O(N__42056),
            .I(N__41659));
    ClkMux I__10346 (
            .O(N__42055),
            .I(N__41659));
    ClkMux I__10345 (
            .O(N__42054),
            .I(N__41659));
    ClkMux I__10344 (
            .O(N__42053),
            .I(N__41659));
    ClkMux I__10343 (
            .O(N__42052),
            .I(N__41659));
    ClkMux I__10342 (
            .O(N__42051),
            .I(N__41659));
    ClkMux I__10341 (
            .O(N__42050),
            .I(N__41659));
    ClkMux I__10340 (
            .O(N__42049),
            .I(N__41659));
    ClkMux I__10339 (
            .O(N__42048),
            .I(N__41659));
    ClkMux I__10338 (
            .O(N__42047),
            .I(N__41659));
    ClkMux I__10337 (
            .O(N__42046),
            .I(N__41659));
    ClkMux I__10336 (
            .O(N__42045),
            .I(N__41659));
    ClkMux I__10335 (
            .O(N__42044),
            .I(N__41659));
    ClkMux I__10334 (
            .O(N__42043),
            .I(N__41659));
    ClkMux I__10333 (
            .O(N__42042),
            .I(N__41659));
    ClkMux I__10332 (
            .O(N__42041),
            .I(N__41659));
    ClkMux I__10331 (
            .O(N__42040),
            .I(N__41659));
    ClkMux I__10330 (
            .O(N__42039),
            .I(N__41659));
    ClkMux I__10329 (
            .O(N__42038),
            .I(N__41659));
    ClkMux I__10328 (
            .O(N__42037),
            .I(N__41659));
    ClkMux I__10327 (
            .O(N__42036),
            .I(N__41659));
    ClkMux I__10326 (
            .O(N__42035),
            .I(N__41659));
    ClkMux I__10325 (
            .O(N__42034),
            .I(N__41659));
    ClkMux I__10324 (
            .O(N__42033),
            .I(N__41659));
    ClkMux I__10323 (
            .O(N__42032),
            .I(N__41659));
    ClkMux I__10322 (
            .O(N__42031),
            .I(N__41659));
    ClkMux I__10321 (
            .O(N__42030),
            .I(N__41659));
    ClkMux I__10320 (
            .O(N__42029),
            .I(N__41659));
    ClkMux I__10319 (
            .O(N__42028),
            .I(N__41659));
    ClkMux I__10318 (
            .O(N__42027),
            .I(N__41659));
    ClkMux I__10317 (
            .O(N__42026),
            .I(N__41659));
    ClkMux I__10316 (
            .O(N__42025),
            .I(N__41659));
    ClkMux I__10315 (
            .O(N__42024),
            .I(N__41659));
    ClkMux I__10314 (
            .O(N__42023),
            .I(N__41659));
    ClkMux I__10313 (
            .O(N__42022),
            .I(N__41659));
    ClkMux I__10312 (
            .O(N__42021),
            .I(N__41659));
    ClkMux I__10311 (
            .O(N__42020),
            .I(N__41659));
    ClkMux I__10310 (
            .O(N__42019),
            .I(N__41659));
    ClkMux I__10309 (
            .O(N__42018),
            .I(N__41659));
    ClkMux I__10308 (
            .O(N__42017),
            .I(N__41659));
    ClkMux I__10307 (
            .O(N__42016),
            .I(N__41659));
    ClkMux I__10306 (
            .O(N__42015),
            .I(N__41659));
    ClkMux I__10305 (
            .O(N__42014),
            .I(N__41659));
    ClkMux I__10304 (
            .O(N__42013),
            .I(N__41659));
    ClkMux I__10303 (
            .O(N__42012),
            .I(N__41659));
    ClkMux I__10302 (
            .O(N__42011),
            .I(N__41659));
    ClkMux I__10301 (
            .O(N__42010),
            .I(N__41659));
    ClkMux I__10300 (
            .O(N__42009),
            .I(N__41659));
    ClkMux I__10299 (
            .O(N__42008),
            .I(N__41659));
    ClkMux I__10298 (
            .O(N__42007),
            .I(N__41659));
    ClkMux I__10297 (
            .O(N__42006),
            .I(N__41659));
    ClkMux I__10296 (
            .O(N__42005),
            .I(N__41659));
    ClkMux I__10295 (
            .O(N__42004),
            .I(N__41659));
    ClkMux I__10294 (
            .O(N__42003),
            .I(N__41659));
    ClkMux I__10293 (
            .O(N__42002),
            .I(N__41659));
    ClkMux I__10292 (
            .O(N__42001),
            .I(N__41659));
    ClkMux I__10291 (
            .O(N__42000),
            .I(N__41659));
    ClkMux I__10290 (
            .O(N__41999),
            .I(N__41659));
    ClkMux I__10289 (
            .O(N__41998),
            .I(N__41659));
    ClkMux I__10288 (
            .O(N__41997),
            .I(N__41659));
    ClkMux I__10287 (
            .O(N__41996),
            .I(N__41659));
    ClkMux I__10286 (
            .O(N__41995),
            .I(N__41659));
    ClkMux I__10285 (
            .O(N__41994),
            .I(N__41659));
    ClkMux I__10284 (
            .O(N__41993),
            .I(N__41659));
    ClkMux I__10283 (
            .O(N__41992),
            .I(N__41659));
    ClkMux I__10282 (
            .O(N__41991),
            .I(N__41659));
    ClkMux I__10281 (
            .O(N__41990),
            .I(N__41659));
    ClkMux I__10280 (
            .O(N__41989),
            .I(N__41659));
    ClkMux I__10279 (
            .O(N__41988),
            .I(N__41659));
    ClkMux I__10278 (
            .O(N__41987),
            .I(N__41659));
    ClkMux I__10277 (
            .O(N__41986),
            .I(N__41659));
    ClkMux I__10276 (
            .O(N__41985),
            .I(N__41659));
    ClkMux I__10275 (
            .O(N__41984),
            .I(N__41659));
    GlobalMux I__10274 (
            .O(N__41659),
            .I(N__41656));
    gio2CtrlBuf I__10273 (
            .O(N__41656),
            .I(clk_0_c_g));
    SRMux I__10272 (
            .O(N__41653),
            .I(N__41608));
    SRMux I__10271 (
            .O(N__41652),
            .I(N__41608));
    SRMux I__10270 (
            .O(N__41651),
            .I(N__41608));
    SRMux I__10269 (
            .O(N__41650),
            .I(N__41608));
    SRMux I__10268 (
            .O(N__41649),
            .I(N__41608));
    SRMux I__10267 (
            .O(N__41648),
            .I(N__41608));
    SRMux I__10266 (
            .O(N__41647),
            .I(N__41608));
    SRMux I__10265 (
            .O(N__41646),
            .I(N__41608));
    SRMux I__10264 (
            .O(N__41645),
            .I(N__41608));
    SRMux I__10263 (
            .O(N__41644),
            .I(N__41608));
    SRMux I__10262 (
            .O(N__41643),
            .I(N__41608));
    SRMux I__10261 (
            .O(N__41642),
            .I(N__41608));
    SRMux I__10260 (
            .O(N__41641),
            .I(N__41608));
    SRMux I__10259 (
            .O(N__41640),
            .I(N__41608));
    SRMux I__10258 (
            .O(N__41639),
            .I(N__41608));
    GlobalMux I__10257 (
            .O(N__41608),
            .I(N__41605));
    gio2CtrlBuf I__10256 (
            .O(N__41605),
            .I(N_620_g));
    InMux I__10255 (
            .O(N__41602),
            .I(N__41598));
    InMux I__10254 (
            .O(N__41601),
            .I(N__41595));
    LocalMux I__10253 (
            .O(N__41598),
            .I(N__41592));
    LocalMux I__10252 (
            .O(N__41595),
            .I(N__41589));
    Span4Mux_v I__10251 (
            .O(N__41592),
            .I(N__41586));
    Span12Mux_s9_h I__10250 (
            .O(N__41589),
            .I(N__41581));
    Sp12to4 I__10249 (
            .O(N__41586),
            .I(N__41581));
    Span12Mux_v I__10248 (
            .O(N__41581),
            .I(N__41578));
    Odrv12 I__10247 (
            .O(N__41578),
            .I(M_this_map_ram_read_data_6));
    IoInMux I__10246 (
            .O(N__41575),
            .I(N__41572));
    LocalMux I__10245 (
            .O(N__41572),
            .I(N__41569));
    Span4Mux_s3_h I__10244 (
            .O(N__41569),
            .I(N__41566));
    Span4Mux_v I__10243 (
            .O(N__41566),
            .I(N__41563));
    Odrv4 I__10242 (
            .O(N__41563),
            .I(N_734_0));
    CascadeMux I__10241 (
            .O(N__41560),
            .I(N__41557));
    CascadeBuf I__10240 (
            .O(N__41557),
            .I(N__41554));
    CascadeMux I__10239 (
            .O(N__41554),
            .I(N__41551));
    InMux I__10238 (
            .O(N__41551),
            .I(N__41546));
    CascadeMux I__10237 (
            .O(N__41550),
            .I(N__41543));
    InMux I__10236 (
            .O(N__41549),
            .I(N__41539));
    LocalMux I__10235 (
            .O(N__41546),
            .I(N__41536));
    InMux I__10234 (
            .O(N__41543),
            .I(N__41533));
    InMux I__10233 (
            .O(N__41542),
            .I(N__41530));
    LocalMux I__10232 (
            .O(N__41539),
            .I(N__41527));
    Span4Mux_v I__10231 (
            .O(N__41536),
            .I(N__41524));
    LocalMux I__10230 (
            .O(N__41533),
            .I(M_this_map_address_qZ0Z_8));
    LocalMux I__10229 (
            .O(N__41530),
            .I(M_this_map_address_qZ0Z_8));
    Odrv4 I__10228 (
            .O(N__41527),
            .I(M_this_map_address_qZ0Z_8));
    Odrv4 I__10227 (
            .O(N__41524),
            .I(M_this_map_address_qZ0Z_8));
    InMux I__10226 (
            .O(N__41515),
            .I(N__41506));
    InMux I__10225 (
            .O(N__41514),
            .I(N__41503));
    InMux I__10224 (
            .O(N__41513),
            .I(N__41500));
    InMux I__10223 (
            .O(N__41512),
            .I(N__41497));
    InMux I__10222 (
            .O(N__41511),
            .I(N__41494));
    InMux I__10221 (
            .O(N__41510),
            .I(N__41491));
    InMux I__10220 (
            .O(N__41509),
            .I(N__41488));
    LocalMux I__10219 (
            .O(N__41506),
            .I(N__41485));
    LocalMux I__10218 (
            .O(N__41503),
            .I(N__41482));
    LocalMux I__10217 (
            .O(N__41500),
            .I(N__41475));
    LocalMux I__10216 (
            .O(N__41497),
            .I(N__41475));
    LocalMux I__10215 (
            .O(N__41494),
            .I(N__41475));
    LocalMux I__10214 (
            .O(N__41491),
            .I(N__41471));
    LocalMux I__10213 (
            .O(N__41488),
            .I(N__41467));
    Span4Mux_h I__10212 (
            .O(N__41485),
            .I(N__41461));
    Span4Mux_v I__10211 (
            .O(N__41482),
            .I(N__41461));
    Span4Mux_v I__10210 (
            .O(N__41475),
            .I(N__41458));
    InMux I__10209 (
            .O(N__41474),
            .I(N__41455));
    Span4Mux_h I__10208 (
            .O(N__41471),
            .I(N__41451));
    InMux I__10207 (
            .O(N__41470),
            .I(N__41448));
    Span4Mux_h I__10206 (
            .O(N__41467),
            .I(N__41445));
    InMux I__10205 (
            .O(N__41466),
            .I(N__41442));
    Span4Mux_v I__10204 (
            .O(N__41461),
            .I(N__41437));
    Span4Mux_h I__10203 (
            .O(N__41458),
            .I(N__41437));
    LocalMux I__10202 (
            .O(N__41455),
            .I(N__41434));
    InMux I__10201 (
            .O(N__41454),
            .I(N__41431));
    Span4Mux_v I__10200 (
            .O(N__41451),
            .I(N__41426));
    LocalMux I__10199 (
            .O(N__41448),
            .I(N__41426));
    Span4Mux_v I__10198 (
            .O(N__41445),
            .I(N__41421));
    LocalMux I__10197 (
            .O(N__41442),
            .I(N__41421));
    Sp12to4 I__10196 (
            .O(N__41437),
            .I(N__41418));
    Span12Mux_v I__10195 (
            .O(N__41434),
            .I(N__41413));
    LocalMux I__10194 (
            .O(N__41431),
            .I(N__41413));
    Span4Mux_h I__10193 (
            .O(N__41426),
            .I(N__41410));
    Span4Mux_v I__10192 (
            .O(N__41421),
            .I(N__41407));
    Span12Mux_h I__10191 (
            .O(N__41418),
            .I(N__41404));
    Span12Mux_h I__10190 (
            .O(N__41413),
            .I(N__41401));
    Span4Mux_v I__10189 (
            .O(N__41410),
            .I(N__41398));
    Span4Mux_h I__10188 (
            .O(N__41407),
            .I(N__41395));
    Odrv12 I__10187 (
            .O(N__41404),
            .I(port_data_in_3));
    Odrv12 I__10186 (
            .O(N__41401),
            .I(port_data_in_3));
    Odrv4 I__10185 (
            .O(N__41398),
            .I(port_data_in_3));
    Odrv4 I__10184 (
            .O(N__41395),
            .I(port_data_in_3));
    CascadeMux I__10183 (
            .O(N__41386),
            .I(N_1078_cascade_));
    InMux I__10182 (
            .O(N__41383),
            .I(N__41380));
    LocalMux I__10181 (
            .O(N__41380),
            .I(N__41377));
    Odrv4 I__10180 (
            .O(N__41377),
            .I(M_this_map_address_qc_0_1));
    InMux I__10179 (
            .O(N__41374),
            .I(N__41371));
    LocalMux I__10178 (
            .O(N__41371),
            .I(N__41368));
    Span4Mux_v I__10177 (
            .O(N__41368),
            .I(N__41365));
    Span4Mux_v I__10176 (
            .O(N__41365),
            .I(N__41361));
    InMux I__10175 (
            .O(N__41364),
            .I(N__41358));
    Sp12to4 I__10174 (
            .O(N__41361),
            .I(N__41355));
    LocalMux I__10173 (
            .O(N__41358),
            .I(M_this_map_ram_read_data_2));
    Odrv12 I__10172 (
            .O(N__41355),
            .I(M_this_map_ram_read_data_2));
    IoInMux I__10171 (
            .O(N__41350),
            .I(N__41347));
    LocalMux I__10170 (
            .O(N__41347),
            .I(N__41344));
    Odrv4 I__10169 (
            .O(N__41344),
            .I(N_726_0));
    InMux I__10168 (
            .O(N__41341),
            .I(N__41338));
    LocalMux I__10167 (
            .O(N__41338),
            .I(un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0));
    IoInMux I__10166 (
            .O(N__41335),
            .I(N__41332));
    LocalMux I__10165 (
            .O(N__41332),
            .I(N__41329));
    Span4Mux_s2_v I__10164 (
            .O(N__41329),
            .I(N__41326));
    Sp12to4 I__10163 (
            .O(N__41326),
            .I(N__41323));
    Span12Mux_h I__10162 (
            .O(N__41323),
            .I(N__41319));
    InMux I__10161 (
            .O(N__41322),
            .I(N__41316));
    Odrv12 I__10160 (
            .O(N__41319),
            .I(M_this_ext_address_qZ0Z_8));
    LocalMux I__10159 (
            .O(N__41316),
            .I(M_this_ext_address_qZ0Z_8));
    InMux I__10158 (
            .O(N__41311),
            .I(N__41308));
    LocalMux I__10157 (
            .O(N__41308),
            .I(un1_M_this_ext_address_q_cry_0_THRU_CO));
    IoInMux I__10156 (
            .O(N__41305),
            .I(N__41302));
    LocalMux I__10155 (
            .O(N__41302),
            .I(N__41299));
    Span4Mux_s2_v I__10154 (
            .O(N__41299),
            .I(N__41296));
    Span4Mux_v I__10153 (
            .O(N__41296),
            .I(N__41292));
    CascadeMux I__10152 (
            .O(N__41295),
            .I(N__41289));
    Span4Mux_v I__10151 (
            .O(N__41292),
            .I(N__41285));
    InMux I__10150 (
            .O(N__41289),
            .I(N__41282));
    InMux I__10149 (
            .O(N__41288),
            .I(N__41279));
    Odrv4 I__10148 (
            .O(N__41285),
            .I(M_this_ext_address_qZ0Z_1));
    LocalMux I__10147 (
            .O(N__41282),
            .I(M_this_ext_address_qZ0Z_1));
    LocalMux I__10146 (
            .O(N__41279),
            .I(M_this_ext_address_qZ0Z_1));
    InMux I__10145 (
            .O(N__41272),
            .I(N__41269));
    LocalMux I__10144 (
            .O(N__41269),
            .I(un1_M_this_ext_address_q_cry_2_THRU_CO));
    IoInMux I__10143 (
            .O(N__41266),
            .I(N__41263));
    LocalMux I__10142 (
            .O(N__41263),
            .I(N__41260));
    IoSpan4Mux I__10141 (
            .O(N__41260),
            .I(N__41257));
    Span4Mux_s3_h I__10140 (
            .O(N__41257),
            .I(N__41253));
    CascadeMux I__10139 (
            .O(N__41256),
            .I(N__41250));
    Span4Mux_v I__10138 (
            .O(N__41253),
            .I(N__41246));
    InMux I__10137 (
            .O(N__41250),
            .I(N__41243));
    InMux I__10136 (
            .O(N__41249),
            .I(N__41240));
    Odrv4 I__10135 (
            .O(N__41246),
            .I(M_this_ext_address_qZ0Z_3));
    LocalMux I__10134 (
            .O(N__41243),
            .I(M_this_ext_address_qZ0Z_3));
    LocalMux I__10133 (
            .O(N__41240),
            .I(M_this_ext_address_qZ0Z_3));
    InMux I__10132 (
            .O(N__41233),
            .I(N__41230));
    LocalMux I__10131 (
            .O(N__41230),
            .I(un1_M_this_ext_address_q_cry_3_THRU_CO));
    IoInMux I__10130 (
            .O(N__41227),
            .I(N__41224));
    LocalMux I__10129 (
            .O(N__41224),
            .I(N__41221));
    IoSpan4Mux I__10128 (
            .O(N__41221),
            .I(N__41218));
    Span4Mux_s0_h I__10127 (
            .O(N__41218),
            .I(N__41215));
    Span4Mux_h I__10126 (
            .O(N__41215),
            .I(N__41210));
    InMux I__10125 (
            .O(N__41214),
            .I(N__41207));
    InMux I__10124 (
            .O(N__41213),
            .I(N__41204));
    Odrv4 I__10123 (
            .O(N__41210),
            .I(M_this_ext_address_qZ0Z_4));
    LocalMux I__10122 (
            .O(N__41207),
            .I(M_this_ext_address_qZ0Z_4));
    LocalMux I__10121 (
            .O(N__41204),
            .I(M_this_ext_address_qZ0Z_4));
    InMux I__10120 (
            .O(N__41197),
            .I(N__41194));
    LocalMux I__10119 (
            .O(N__41194),
            .I(un1_M_this_ext_address_q_cry_4_THRU_CO));
    IoInMux I__10118 (
            .O(N__41191),
            .I(N__41188));
    LocalMux I__10117 (
            .O(N__41188),
            .I(N__41185));
    IoSpan4Mux I__10116 (
            .O(N__41185),
            .I(N__41181));
    CascadeMux I__10115 (
            .O(N__41184),
            .I(N__41178));
    Span4Mux_s2_h I__10114 (
            .O(N__41181),
            .I(N__41174));
    InMux I__10113 (
            .O(N__41178),
            .I(N__41171));
    InMux I__10112 (
            .O(N__41177),
            .I(N__41168));
    Odrv4 I__10111 (
            .O(N__41174),
            .I(M_this_ext_address_qZ0Z_5));
    LocalMux I__10110 (
            .O(N__41171),
            .I(M_this_ext_address_qZ0Z_5));
    LocalMux I__10109 (
            .O(N__41168),
            .I(M_this_ext_address_qZ0Z_5));
    CascadeMux I__10108 (
            .O(N__41161),
            .I(N__41157));
    CascadeMux I__10107 (
            .O(N__41160),
            .I(N__41154));
    InMux I__10106 (
            .O(N__41157),
            .I(N__41146));
    InMux I__10105 (
            .O(N__41154),
            .I(N__41146));
    CascadeMux I__10104 (
            .O(N__41153),
            .I(N__41142));
    InMux I__10103 (
            .O(N__41152),
            .I(N__41137));
    InMux I__10102 (
            .O(N__41151),
            .I(N__41137));
    LocalMux I__10101 (
            .O(N__41146),
            .I(N__41126));
    InMux I__10100 (
            .O(N__41145),
            .I(N__41123));
    InMux I__10099 (
            .O(N__41142),
            .I(N__41120));
    LocalMux I__10098 (
            .O(N__41137),
            .I(N__41117));
    InMux I__10097 (
            .O(N__41136),
            .I(N__41104));
    InMux I__10096 (
            .O(N__41135),
            .I(N__41104));
    InMux I__10095 (
            .O(N__41134),
            .I(N__41104));
    InMux I__10094 (
            .O(N__41133),
            .I(N__41104));
    InMux I__10093 (
            .O(N__41132),
            .I(N__41104));
    InMux I__10092 (
            .O(N__41131),
            .I(N__41104));
    CascadeMux I__10091 (
            .O(N__41130),
            .I(N__41101));
    CascadeMux I__10090 (
            .O(N__41129),
            .I(N__41098));
    Span4Mux_h I__10089 (
            .O(N__41126),
            .I(N__41092));
    LocalMux I__10088 (
            .O(N__41123),
            .I(N__41085));
    LocalMux I__10087 (
            .O(N__41120),
            .I(N__41085));
    Span4Mux_h I__10086 (
            .O(N__41117),
            .I(N__41085));
    LocalMux I__10085 (
            .O(N__41104),
            .I(N__41082));
    InMux I__10084 (
            .O(N__41101),
            .I(N__41079));
    InMux I__10083 (
            .O(N__41098),
            .I(N__41076));
    InMux I__10082 (
            .O(N__41097),
            .I(N__41069));
    InMux I__10081 (
            .O(N__41096),
            .I(N__41069));
    InMux I__10080 (
            .O(N__41095),
            .I(N__41069));
    Span4Mux_v I__10079 (
            .O(N__41092),
            .I(N__41062));
    Span4Mux_v I__10078 (
            .O(N__41085),
            .I(N__41062));
    Span4Mux_h I__10077 (
            .O(N__41082),
            .I(N__41062));
    LocalMux I__10076 (
            .O(N__41079),
            .I(N__41053));
    LocalMux I__10075 (
            .O(N__41076),
            .I(N__41053));
    LocalMux I__10074 (
            .O(N__41069),
            .I(N__41053));
    Span4Mux_h I__10073 (
            .O(N__41062),
            .I(N__41050));
    InMux I__10072 (
            .O(N__41061),
            .I(N__41045));
    InMux I__10071 (
            .O(N__41060),
            .I(N__41045));
    Odrv12 I__10070 (
            .O(N__41053),
            .I(N_773_0));
    Odrv4 I__10069 (
            .O(N__41050),
            .I(N_773_0));
    LocalMux I__10068 (
            .O(N__41045),
            .I(N_773_0));
    InMux I__10067 (
            .O(N__41038),
            .I(un1_M_this_ext_address_q_cry_14));
    InMux I__10066 (
            .O(N__41035),
            .I(N__41032));
    LocalMux I__10065 (
            .O(N__41032),
            .I(N__41029));
    Odrv12 I__10064 (
            .O(N__41029),
            .I(un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0));
    InMux I__10063 (
            .O(N__41026),
            .I(N__41023));
    LocalMux I__10062 (
            .O(N__41023),
            .I(un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0));
    IoInMux I__10061 (
            .O(N__41020),
            .I(N__41017));
    LocalMux I__10060 (
            .O(N__41017),
            .I(N__41014));
    Span4Mux_s1_v I__10059 (
            .O(N__41014),
            .I(N__41011));
    Span4Mux_v I__10058 (
            .O(N__41011),
            .I(N__41008));
    Span4Mux_v I__10057 (
            .O(N__41008),
            .I(N__41005));
    Span4Mux_h I__10056 (
            .O(N__41005),
            .I(N__41001));
    InMux I__10055 (
            .O(N__41004),
            .I(N__40998));
    Odrv4 I__10054 (
            .O(N__41001),
            .I(M_this_ext_address_qZ0Z_10));
    LocalMux I__10053 (
            .O(N__40998),
            .I(M_this_ext_address_qZ0Z_10));
    InMux I__10052 (
            .O(N__40993),
            .I(N__40990));
    LocalMux I__10051 (
            .O(N__40990),
            .I(N__40987));
    Odrv4 I__10050 (
            .O(N__40987),
            .I(un1_M_this_ext_address_q_cry_6_THRU_CO));
    IoInMux I__10049 (
            .O(N__40984),
            .I(N__40981));
    LocalMux I__10048 (
            .O(N__40981),
            .I(N__40978));
    Span4Mux_s2_h I__10047 (
            .O(N__40978),
            .I(N__40975));
    Span4Mux_h I__10046 (
            .O(N__40975),
            .I(N__40972));
    Sp12to4 I__10045 (
            .O(N__40972),
            .I(N__40968));
    InMux I__10044 (
            .O(N__40971),
            .I(N__40964));
    Span12Mux_s11_v I__10043 (
            .O(N__40968),
            .I(N__40961));
    InMux I__10042 (
            .O(N__40967),
            .I(N__40958));
    LocalMux I__10041 (
            .O(N__40964),
            .I(N__40955));
    Odrv12 I__10040 (
            .O(N__40961),
            .I(M_this_ext_address_qZ0Z_7));
    LocalMux I__10039 (
            .O(N__40958),
            .I(M_this_ext_address_qZ0Z_7));
    Odrv4 I__10038 (
            .O(N__40955),
            .I(M_this_ext_address_qZ0Z_7));
    InMux I__10037 (
            .O(N__40948),
            .I(N__40945));
    LocalMux I__10036 (
            .O(N__40945),
            .I(un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0));
    IoInMux I__10035 (
            .O(N__40942),
            .I(N__40939));
    LocalMux I__10034 (
            .O(N__40939),
            .I(N__40936));
    Span4Mux_s2_v I__10033 (
            .O(N__40936),
            .I(N__40933));
    Span4Mux_h I__10032 (
            .O(N__40933),
            .I(N__40930));
    Span4Mux_v I__10031 (
            .O(N__40930),
            .I(N__40926));
    InMux I__10030 (
            .O(N__40929),
            .I(N__40923));
    Odrv4 I__10029 (
            .O(N__40926),
            .I(M_this_ext_address_qZ0Z_11));
    LocalMux I__10028 (
            .O(N__40923),
            .I(M_this_ext_address_qZ0Z_11));
    InMux I__10027 (
            .O(N__40918),
            .I(N__40915));
    LocalMux I__10026 (
            .O(N__40915),
            .I(un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0));
    IoInMux I__10025 (
            .O(N__40912),
            .I(N__40909));
    LocalMux I__10024 (
            .O(N__40909),
            .I(N__40906));
    Span4Mux_s1_h I__10023 (
            .O(N__40906),
            .I(N__40903));
    Span4Mux_h I__10022 (
            .O(N__40903),
            .I(N__40899));
    InMux I__10021 (
            .O(N__40902),
            .I(N__40896));
    Odrv4 I__10020 (
            .O(N__40899),
            .I(M_this_ext_address_qZ0Z_12));
    LocalMux I__10019 (
            .O(N__40896),
            .I(M_this_ext_address_qZ0Z_12));
    InMux I__10018 (
            .O(N__40891),
            .I(N__40885));
    InMux I__10017 (
            .O(N__40890),
            .I(N__40885));
    LocalMux I__10016 (
            .O(N__40885),
            .I(N__40882));
    Span4Mux_v I__10015 (
            .O(N__40882),
            .I(N__40877));
    InMux I__10014 (
            .O(N__40881),
            .I(N__40874));
    InMux I__10013 (
            .O(N__40880),
            .I(N__40871));
    Span4Mux_v I__10012 (
            .O(N__40877),
            .I(N__40866));
    LocalMux I__10011 (
            .O(N__40874),
            .I(N__40866));
    LocalMux I__10010 (
            .O(N__40871),
            .I(N__40863));
    Span4Mux_h I__10009 (
            .O(N__40866),
            .I(N__40858));
    Span4Mux_h I__10008 (
            .O(N__40863),
            .I(N__40855));
    InMux I__10007 (
            .O(N__40862),
            .I(N__40852));
    InMux I__10006 (
            .O(N__40861),
            .I(N__40849));
    Odrv4 I__10005 (
            .O(N__40858),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__10004 (
            .O(N__40855),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__10003 (
            .O(N__40852),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__10002 (
            .O(N__40849),
            .I(M_this_state_qZ0Z_1));
    InMux I__10001 (
            .O(N__40840),
            .I(N__40836));
    InMux I__10000 (
            .O(N__40839),
            .I(N__40833));
    LocalMux I__9999 (
            .O(N__40836),
            .I(N__40830));
    LocalMux I__9998 (
            .O(N__40833),
            .I(M_this_ctrl_flags_qZ0Z_4));
    Odrv4 I__9997 (
            .O(N__40830),
            .I(M_this_ctrl_flags_qZ0Z_4));
    CascadeMux I__9996 (
            .O(N__40825),
            .I(N__40822));
    CascadeBuf I__9995 (
            .O(N__40822),
            .I(N__40819));
    CascadeMux I__9994 (
            .O(N__40819),
            .I(N__40816));
    InMux I__9993 (
            .O(N__40816),
            .I(N__40813));
    LocalMux I__9992 (
            .O(N__40813),
            .I(N__40809));
    InMux I__9991 (
            .O(N__40812),
            .I(N__40805));
    Span4Mux_s3_v I__9990 (
            .O(N__40809),
            .I(N__40802));
    InMux I__9989 (
            .O(N__40808),
            .I(N__40799));
    LocalMux I__9988 (
            .O(N__40805),
            .I(N__40796));
    Span4Mux_v I__9987 (
            .O(N__40802),
            .I(N__40793));
    LocalMux I__9986 (
            .O(N__40799),
            .I(M_this_map_address_qZ0Z_9));
    Odrv4 I__9985 (
            .O(N__40796),
            .I(M_this_map_address_qZ0Z_9));
    Odrv4 I__9984 (
            .O(N__40793),
            .I(M_this_map_address_qZ0Z_9));
    InMux I__9983 (
            .O(N__40786),
            .I(N__40779));
    InMux I__9982 (
            .O(N__40785),
            .I(N__40776));
    InMux I__9981 (
            .O(N__40784),
            .I(N__40773));
    InMux I__9980 (
            .O(N__40783),
            .I(N__40770));
    InMux I__9979 (
            .O(N__40782),
            .I(N__40767));
    LocalMux I__9978 (
            .O(N__40779),
            .I(N__40764));
    LocalMux I__9977 (
            .O(N__40776),
            .I(N__40760));
    LocalMux I__9976 (
            .O(N__40773),
            .I(N__40757));
    LocalMux I__9975 (
            .O(N__40770),
            .I(N__40752));
    LocalMux I__9974 (
            .O(N__40767),
            .I(N__40752));
    Span4Mux_v I__9973 (
            .O(N__40764),
            .I(N__40748));
    InMux I__9972 (
            .O(N__40763),
            .I(N__40744));
    Span4Mux_h I__9971 (
            .O(N__40760),
            .I(N__40739));
    Span4Mux_v I__9970 (
            .O(N__40757),
            .I(N__40739));
    Span4Mux_v I__9969 (
            .O(N__40752),
            .I(N__40736));
    InMux I__9968 (
            .O(N__40751),
            .I(N__40733));
    Span4Mux_v I__9967 (
            .O(N__40748),
            .I(N__40730));
    InMux I__9966 (
            .O(N__40747),
            .I(N__40727));
    LocalMux I__9965 (
            .O(N__40744),
            .I(N__40723));
    Span4Mux_v I__9964 (
            .O(N__40739),
            .I(N__40718));
    Span4Mux_h I__9963 (
            .O(N__40736),
            .I(N__40718));
    LocalMux I__9962 (
            .O(N__40733),
            .I(N__40715));
    Span4Mux_h I__9961 (
            .O(N__40730),
            .I(N__40710));
    LocalMux I__9960 (
            .O(N__40727),
            .I(N__40710));
    CascadeMux I__9959 (
            .O(N__40726),
            .I(N__40706));
    Span4Mux_v I__9958 (
            .O(N__40723),
            .I(N__40702));
    Span4Mux_h I__9957 (
            .O(N__40718),
            .I(N__40697));
    Span4Mux_v I__9956 (
            .O(N__40715),
            .I(N__40697));
    Span4Mux_h I__9955 (
            .O(N__40710),
            .I(N__40694));
    InMux I__9954 (
            .O(N__40709),
            .I(N__40689));
    InMux I__9953 (
            .O(N__40706),
            .I(N__40689));
    InMux I__9952 (
            .O(N__40705),
            .I(N__40686));
    Sp12to4 I__9951 (
            .O(N__40702),
            .I(N__40680));
    Sp12to4 I__9950 (
            .O(N__40697),
            .I(N__40680));
    Span4Mux_v I__9949 (
            .O(N__40694),
            .I(N__40677));
    LocalMux I__9948 (
            .O(N__40689),
            .I(N__40672));
    LocalMux I__9947 (
            .O(N__40686),
            .I(N__40672));
    InMux I__9946 (
            .O(N__40685),
            .I(N__40669));
    Span12Mux_h I__9945 (
            .O(N__40680),
            .I(N__40662));
    Sp12to4 I__9944 (
            .O(N__40677),
            .I(N__40662));
    Span12Mux_v I__9943 (
            .O(N__40672),
            .I(N__40662));
    LocalMux I__9942 (
            .O(N__40669),
            .I(N__40659));
    Odrv12 I__9941 (
            .O(N__40662),
            .I(port_data_in_4));
    Odrv12 I__9940 (
            .O(N__40659),
            .I(port_data_in_4));
    CascadeMux I__9939 (
            .O(N__40654),
            .I(N_1081_cascade_));
    InMux I__9938 (
            .O(N__40651),
            .I(N__40648));
    LocalMux I__9937 (
            .O(N__40648),
            .I(N__40645));
    Odrv4 I__9936 (
            .O(N__40645),
            .I(M_this_map_address_qc_1_1));
    InMux I__9935 (
            .O(N__40642),
            .I(un1_M_this_ext_address_q_cry_6));
    InMux I__9934 (
            .O(N__40639),
            .I(bfn_26_22_0_));
    IoInMux I__9933 (
            .O(N__40636),
            .I(N__40633));
    LocalMux I__9932 (
            .O(N__40633),
            .I(N__40630));
    IoSpan4Mux I__9931 (
            .O(N__40630),
            .I(N__40627));
    Span4Mux_s2_v I__9930 (
            .O(N__40627),
            .I(N__40623));
    InMux I__9929 (
            .O(N__40626),
            .I(N__40620));
    Span4Mux_v I__9928 (
            .O(N__40623),
            .I(N__40617));
    LocalMux I__9927 (
            .O(N__40620),
            .I(N__40614));
    Span4Mux_v I__9926 (
            .O(N__40617),
            .I(N__40609));
    Span4Mux_h I__9925 (
            .O(N__40614),
            .I(N__40609));
    Odrv4 I__9924 (
            .O(N__40609),
            .I(M_this_ext_address_qZ0Z_9));
    InMux I__9923 (
            .O(N__40606),
            .I(N__40603));
    LocalMux I__9922 (
            .O(N__40603),
            .I(N__40600));
    Span4Mux_h I__9921 (
            .O(N__40600),
            .I(N__40597));
    Odrv4 I__9920 (
            .O(N__40597),
            .I(un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0));
    InMux I__9919 (
            .O(N__40594),
            .I(un1_M_this_ext_address_q_cry_8));
    InMux I__9918 (
            .O(N__40591),
            .I(un1_M_this_ext_address_q_cry_9));
    InMux I__9917 (
            .O(N__40588),
            .I(un1_M_this_ext_address_q_cry_10));
    InMux I__9916 (
            .O(N__40585),
            .I(un1_M_this_ext_address_q_cry_11));
    IoInMux I__9915 (
            .O(N__40582),
            .I(N__40579));
    LocalMux I__9914 (
            .O(N__40579),
            .I(N__40576));
    IoSpan4Mux I__9913 (
            .O(N__40576),
            .I(N__40573));
    Span4Mux_s2_h I__9912 (
            .O(N__40573),
            .I(N__40569));
    InMux I__9911 (
            .O(N__40572),
            .I(N__40566));
    Span4Mux_h I__9910 (
            .O(N__40569),
            .I(N__40561));
    LocalMux I__9909 (
            .O(N__40566),
            .I(N__40561));
    Span4Mux_v I__9908 (
            .O(N__40561),
            .I(N__40558));
    Odrv4 I__9907 (
            .O(N__40558),
            .I(M_this_ext_address_qZ0Z_13));
    InMux I__9906 (
            .O(N__40555),
            .I(N__40552));
    LocalMux I__9905 (
            .O(N__40552),
            .I(N__40549));
    Odrv12 I__9904 (
            .O(N__40549),
            .I(un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0));
    InMux I__9903 (
            .O(N__40546),
            .I(un1_M_this_ext_address_q_cry_12));
    IoInMux I__9902 (
            .O(N__40543),
            .I(N__40540));
    LocalMux I__9901 (
            .O(N__40540),
            .I(N__40537));
    Span4Mux_s2_h I__9900 (
            .O(N__40537),
            .I(N__40533));
    InMux I__9899 (
            .O(N__40536),
            .I(N__40530));
    Span4Mux_h I__9898 (
            .O(N__40533),
            .I(N__40527));
    LocalMux I__9897 (
            .O(N__40530),
            .I(N__40524));
    Odrv4 I__9896 (
            .O(N__40527),
            .I(M_this_ext_address_qZ0Z_14));
    Odrv12 I__9895 (
            .O(N__40524),
            .I(M_this_ext_address_qZ0Z_14));
    InMux I__9894 (
            .O(N__40519),
            .I(N__40516));
    LocalMux I__9893 (
            .O(N__40516),
            .I(N__40513));
    Odrv12 I__9892 (
            .O(N__40513),
            .I(un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0));
    InMux I__9891 (
            .O(N__40510),
            .I(un1_M_this_ext_address_q_cry_13));
    IoInMux I__9890 (
            .O(N__40507),
            .I(N__40504));
    LocalMux I__9889 (
            .O(N__40504),
            .I(N__40500));
    InMux I__9888 (
            .O(N__40503),
            .I(N__40497));
    Span12Mux_s1_h I__9887 (
            .O(N__40500),
            .I(N__40494));
    LocalMux I__9886 (
            .O(N__40497),
            .I(N__40491));
    Span12Mux_v I__9885 (
            .O(N__40494),
            .I(N__40488));
    Span4Mux_v I__9884 (
            .O(N__40491),
            .I(N__40485));
    Odrv12 I__9883 (
            .O(N__40488),
            .I(M_this_ext_address_qZ0Z_15));
    Odrv4 I__9882 (
            .O(N__40485),
            .I(M_this_ext_address_qZ0Z_15));
    CascadeMux I__9881 (
            .O(N__40480),
            .I(N__40476));
    InMux I__9880 (
            .O(N__40479),
            .I(N__40473));
    InMux I__9879 (
            .O(N__40476),
            .I(N__40470));
    LocalMux I__9878 (
            .O(N__40473),
            .I(N__40467));
    LocalMux I__9877 (
            .O(N__40470),
            .I(N__40464));
    Span4Mux_v I__9876 (
            .O(N__40467),
            .I(N__40459));
    Span4Mux_v I__9875 (
            .O(N__40464),
            .I(N__40459));
    Span4Mux_h I__9874 (
            .O(N__40459),
            .I(N__40455));
    InMux I__9873 (
            .O(N__40458),
            .I(N__40452));
    Span4Mux_h I__9872 (
            .O(N__40455),
            .I(N__40449));
    LocalMux I__9871 (
            .O(N__40452),
            .I(M_this_ctrl_flags_qZ0Z_6));
    Odrv4 I__9870 (
            .O(N__40449),
            .I(M_this_ctrl_flags_qZ0Z_6));
    InMux I__9869 (
            .O(N__40444),
            .I(N__40440));
    InMux I__9868 (
            .O(N__40443),
            .I(N__40437));
    LocalMux I__9867 (
            .O(N__40440),
            .I(N__40430));
    LocalMux I__9866 (
            .O(N__40437),
            .I(N__40430));
    CascadeMux I__9865 (
            .O(N__40436),
            .I(N__40427));
    InMux I__9864 (
            .O(N__40435),
            .I(N__40424));
    Span4Mux_v I__9863 (
            .O(N__40430),
            .I(N__40421));
    InMux I__9862 (
            .O(N__40427),
            .I(N__40416));
    LocalMux I__9861 (
            .O(N__40424),
            .I(N__40412));
    Span4Mux_h I__9860 (
            .O(N__40421),
            .I(N__40408));
    InMux I__9859 (
            .O(N__40420),
            .I(N__40405));
    CascadeMux I__9858 (
            .O(N__40419),
            .I(N__40401));
    LocalMux I__9857 (
            .O(N__40416),
            .I(N__40398));
    InMux I__9856 (
            .O(N__40415),
            .I(N__40394));
    Span4Mux_v I__9855 (
            .O(N__40412),
            .I(N__40391));
    InMux I__9854 (
            .O(N__40411),
            .I(N__40388));
    Span4Mux_v I__9853 (
            .O(N__40408),
            .I(N__40383));
    LocalMux I__9852 (
            .O(N__40405),
            .I(N__40383));
    InMux I__9851 (
            .O(N__40404),
            .I(N__40378));
    InMux I__9850 (
            .O(N__40401),
            .I(N__40378));
    Span4Mux_v I__9849 (
            .O(N__40398),
            .I(N__40375));
    InMux I__9848 (
            .O(N__40397),
            .I(N__40372));
    LocalMux I__9847 (
            .O(N__40394),
            .I(N__40369));
    Span4Mux_h I__9846 (
            .O(N__40391),
            .I(N__40364));
    LocalMux I__9845 (
            .O(N__40388),
            .I(N__40364));
    Span4Mux_v I__9844 (
            .O(N__40383),
            .I(N__40361));
    LocalMux I__9843 (
            .O(N__40378),
            .I(N__40358));
    Span4Mux_h I__9842 (
            .O(N__40375),
            .I(N__40355));
    LocalMux I__9841 (
            .O(N__40372),
            .I(N__40352));
    Span12Mux_h I__9840 (
            .O(N__40369),
            .I(N__40347));
    Sp12to4 I__9839 (
            .O(N__40364),
            .I(N__40347));
    Span4Mux_v I__9838 (
            .O(N__40361),
            .I(N__40344));
    Span4Mux_v I__9837 (
            .O(N__40358),
            .I(N__40341));
    Sp12to4 I__9836 (
            .O(N__40355),
            .I(N__40336));
    Span12Mux_s9_v I__9835 (
            .O(N__40352),
            .I(N__40336));
    Span12Mux_v I__9834 (
            .O(N__40347),
            .I(N__40331));
    Sp12to4 I__9833 (
            .O(N__40344),
            .I(N__40331));
    Span4Mux_h I__9832 (
            .O(N__40341),
            .I(N__40328));
    Span12Mux_v I__9831 (
            .O(N__40336),
            .I(N__40325));
    Span12Mux_h I__9830 (
            .O(N__40331),
            .I(N__40322));
    Span4Mux_v I__9829 (
            .O(N__40328),
            .I(N__40319));
    Odrv12 I__9828 (
            .O(N__40325),
            .I(port_data_in_6));
    Odrv12 I__9827 (
            .O(N__40322),
            .I(port_data_in_6));
    Odrv4 I__9826 (
            .O(N__40319),
            .I(port_data_in_6));
    InMux I__9825 (
            .O(N__40312),
            .I(N__40308));
    InMux I__9824 (
            .O(N__40311),
            .I(N__40305));
    LocalMux I__9823 (
            .O(N__40308),
            .I(N__40300));
    LocalMux I__9822 (
            .O(N__40305),
            .I(N__40300));
    Span4Mux_h I__9821 (
            .O(N__40300),
            .I(N__40297));
    Span4Mux_h I__9820 (
            .O(N__40297),
            .I(N__40294));
    Odrv4 I__9819 (
            .O(N__40294),
            .I(N_247));
    IoInMux I__9818 (
            .O(N__40291),
            .I(N__40288));
    LocalMux I__9817 (
            .O(N__40288),
            .I(N__40285));
    IoSpan4Mux I__9816 (
            .O(N__40285),
            .I(N__40282));
    Span4Mux_s3_v I__9815 (
            .O(N__40282),
            .I(N__40277));
    CascadeMux I__9814 (
            .O(N__40281),
            .I(N__40274));
    CascadeMux I__9813 (
            .O(N__40280),
            .I(N__40271));
    Sp12to4 I__9812 (
            .O(N__40277),
            .I(N__40268));
    InMux I__9811 (
            .O(N__40274),
            .I(N__40265));
    InMux I__9810 (
            .O(N__40271),
            .I(N__40262));
    Span12Mux_s11_v I__9809 (
            .O(N__40268),
            .I(N__40259));
    LocalMux I__9808 (
            .O(N__40265),
            .I(N__40254));
    LocalMux I__9807 (
            .O(N__40262),
            .I(N__40254));
    Odrv12 I__9806 (
            .O(N__40259),
            .I(M_this_ext_address_qZ0Z_0));
    Odrv4 I__9805 (
            .O(N__40254),
            .I(M_this_ext_address_qZ0Z_0));
    InMux I__9804 (
            .O(N__40249),
            .I(un1_M_this_ext_address_q_cry_0));
    IoInMux I__9803 (
            .O(N__40246),
            .I(N__40243));
    LocalMux I__9802 (
            .O(N__40243),
            .I(N__40240));
    IoSpan4Mux I__9801 (
            .O(N__40240),
            .I(N__40237));
    Span4Mux_s3_v I__9800 (
            .O(N__40237),
            .I(N__40233));
    CascadeMux I__9799 (
            .O(N__40236),
            .I(N__40229));
    Span4Mux_v I__9798 (
            .O(N__40233),
            .I(N__40226));
    InMux I__9797 (
            .O(N__40232),
            .I(N__40223));
    InMux I__9796 (
            .O(N__40229),
            .I(N__40220));
    Span4Mux_v I__9795 (
            .O(N__40226),
            .I(N__40215));
    LocalMux I__9794 (
            .O(N__40223),
            .I(N__40215));
    LocalMux I__9793 (
            .O(N__40220),
            .I(M_this_ext_address_qZ0Z_2));
    Odrv4 I__9792 (
            .O(N__40215),
            .I(M_this_ext_address_qZ0Z_2));
    InMux I__9791 (
            .O(N__40210),
            .I(N__40207));
    LocalMux I__9790 (
            .O(N__40207),
            .I(N__40204));
    Odrv4 I__9789 (
            .O(N__40204),
            .I(un1_M_this_ext_address_q_cry_1_THRU_CO));
    InMux I__9788 (
            .O(N__40201),
            .I(un1_M_this_ext_address_q_cry_1));
    InMux I__9787 (
            .O(N__40198),
            .I(un1_M_this_ext_address_q_cry_2));
    InMux I__9786 (
            .O(N__40195),
            .I(un1_M_this_ext_address_q_cry_3));
    InMux I__9785 (
            .O(N__40192),
            .I(un1_M_this_ext_address_q_cry_4));
    InMux I__9784 (
            .O(N__40189),
            .I(un1_M_this_ext_address_q_cry_5));
    InMux I__9783 (
            .O(N__40186),
            .I(N__40183));
    LocalMux I__9782 (
            .O(N__40183),
            .I(N_919_0));
    InMux I__9781 (
            .O(N__40180),
            .I(N__40177));
    LocalMux I__9780 (
            .O(N__40177),
            .I(N__40174));
    Odrv4 I__9779 (
            .O(N__40174),
            .I(N_923_0));
    InMux I__9778 (
            .O(N__40171),
            .I(N__40168));
    LocalMux I__9777 (
            .O(N__40168),
            .I(N_920_0));
    InMux I__9776 (
            .O(N__40165),
            .I(N__40162));
    LocalMux I__9775 (
            .O(N__40162),
            .I(N__40159));
    Odrv4 I__9774 (
            .O(N__40159),
            .I(N_922_0));
    CEMux I__9773 (
            .O(N__40156),
            .I(N__40146));
    InMux I__9772 (
            .O(N__40155),
            .I(N__40141));
    InMux I__9771 (
            .O(N__40154),
            .I(N__40141));
    InMux I__9770 (
            .O(N__40153),
            .I(N__40136));
    InMux I__9769 (
            .O(N__40152),
            .I(N__40136));
    InMux I__9768 (
            .O(N__40151),
            .I(N__40133));
    InMux I__9767 (
            .O(N__40150),
            .I(N__40130));
    CEMux I__9766 (
            .O(N__40149),
            .I(N__40126));
    LocalMux I__9765 (
            .O(N__40146),
            .I(N__40123));
    LocalMux I__9764 (
            .O(N__40141),
            .I(N__40113));
    LocalMux I__9763 (
            .O(N__40136),
            .I(N__40113));
    LocalMux I__9762 (
            .O(N__40133),
            .I(N__40113));
    LocalMux I__9761 (
            .O(N__40130),
            .I(N__40113));
    InMux I__9760 (
            .O(N__40129),
            .I(N__40110));
    LocalMux I__9759 (
            .O(N__40126),
            .I(N__40107));
    Span4Mux_s2_v I__9758 (
            .O(N__40123),
            .I(N__40104));
    InMux I__9757 (
            .O(N__40122),
            .I(N__40101));
    Span4Mux_v I__9756 (
            .O(N__40113),
            .I(N__40096));
    LocalMux I__9755 (
            .O(N__40110),
            .I(N__40096));
    Span4Mux_h I__9754 (
            .O(N__40107),
            .I(N__40093));
    Span4Mux_h I__9753 (
            .O(N__40104),
            .I(N__40088));
    LocalMux I__9752 (
            .O(N__40101),
            .I(N__40088));
    Span4Mux_v I__9751 (
            .O(N__40096),
            .I(N__40085));
    Span4Mux_v I__9750 (
            .O(N__40093),
            .I(N__40080));
    Span4Mux_v I__9749 (
            .O(N__40088),
            .I(N__40080));
    Odrv4 I__9748 (
            .O(N__40085),
            .I(N_296_0));
    Odrv4 I__9747 (
            .O(N__40080),
            .I(N_296_0));
    InMux I__9746 (
            .O(N__40075),
            .I(N__40072));
    LocalMux I__9745 (
            .O(N__40072),
            .I(N_924_0));
    InMux I__9744 (
            .O(N__40069),
            .I(N__40065));
    InMux I__9743 (
            .O(N__40068),
            .I(N__40062));
    LocalMux I__9742 (
            .O(N__40065),
            .I(N__40053));
    LocalMux I__9741 (
            .O(N__40062),
            .I(N__40053));
    InMux I__9740 (
            .O(N__40061),
            .I(N__40049));
    InMux I__9739 (
            .O(N__40060),
            .I(N__40046));
    InMux I__9738 (
            .O(N__40059),
            .I(N__40043));
    InMux I__9737 (
            .O(N__40058),
            .I(N__40040));
    Span4Mux_v I__9736 (
            .O(N__40053),
            .I(N__40036));
    CascadeMux I__9735 (
            .O(N__40052),
            .I(N__40033));
    LocalMux I__9734 (
            .O(N__40049),
            .I(N__40029));
    LocalMux I__9733 (
            .O(N__40046),
            .I(N__40022));
    LocalMux I__9732 (
            .O(N__40043),
            .I(N__40022));
    LocalMux I__9731 (
            .O(N__40040),
            .I(N__40022));
    InMux I__9730 (
            .O(N__40039),
            .I(N__40019));
    Span4Mux_h I__9729 (
            .O(N__40036),
            .I(N__40016));
    InMux I__9728 (
            .O(N__40033),
            .I(N__40013));
    CascadeMux I__9727 (
            .O(N__40032),
            .I(N__40009));
    Span4Mux_v I__9726 (
            .O(N__40029),
            .I(N__40006));
    Span4Mux_v I__9725 (
            .O(N__40022),
            .I(N__40003));
    LocalMux I__9724 (
            .O(N__40019),
            .I(N__40000));
    Span4Mux_h I__9723 (
            .O(N__40016),
            .I(N__39995));
    LocalMux I__9722 (
            .O(N__40013),
            .I(N__39995));
    InMux I__9721 (
            .O(N__40012),
            .I(N__39990));
    InMux I__9720 (
            .O(N__40009),
            .I(N__39990));
    Span4Mux_v I__9719 (
            .O(N__40006),
            .I(N__39987));
    Span4Mux_v I__9718 (
            .O(N__40003),
            .I(N__39982));
    Span4Mux_v I__9717 (
            .O(N__40000),
            .I(N__39982));
    Span4Mux_v I__9716 (
            .O(N__39995),
            .I(N__39979));
    LocalMux I__9715 (
            .O(N__39990),
            .I(N__39976));
    Span4Mux_v I__9714 (
            .O(N__39987),
            .I(N__39973));
    Sp12to4 I__9713 (
            .O(N__39982),
            .I(N__39970));
    Span4Mux_h I__9712 (
            .O(N__39979),
            .I(N__39965));
    Span4Mux_v I__9711 (
            .O(N__39976),
            .I(N__39965));
    Sp12to4 I__9710 (
            .O(N__39973),
            .I(N__39960));
    Span12Mux_h I__9709 (
            .O(N__39970),
            .I(N__39960));
    Span4Mux_h I__9708 (
            .O(N__39965),
            .I(N__39957));
    Odrv12 I__9707 (
            .O(N__39960),
            .I(port_data_in_5));
    Odrv4 I__9706 (
            .O(N__39957),
            .I(port_data_in_5));
    CascadeMux I__9705 (
            .O(N__39952),
            .I(N__39949));
    InMux I__9704 (
            .O(N__39949),
            .I(N__39946));
    LocalMux I__9703 (
            .O(N__39946),
            .I(N__39942));
    InMux I__9702 (
            .O(N__39945),
            .I(N__39939));
    Span12Mux_h I__9701 (
            .O(N__39942),
            .I(N__39936));
    LocalMux I__9700 (
            .O(N__39939),
            .I(M_this_ctrl_flags_qZ0Z_5));
    Odrv12 I__9699 (
            .O(N__39936),
            .I(M_this_ctrl_flags_qZ0Z_5));
    InMux I__9698 (
            .O(N__39931),
            .I(N__39928));
    LocalMux I__9697 (
            .O(N__39928),
            .I(N__39923));
    InMux I__9696 (
            .O(N__39927),
            .I(N__39920));
    InMux I__9695 (
            .O(N__39926),
            .I(N__39917));
    Span4Mux_h I__9694 (
            .O(N__39923),
            .I(N__39910));
    LocalMux I__9693 (
            .O(N__39920),
            .I(N__39910));
    LocalMux I__9692 (
            .O(N__39917),
            .I(N__39910));
    Span4Mux_v I__9691 (
            .O(N__39910),
            .I(N__39907));
    Span4Mux_h I__9690 (
            .O(N__39907),
            .I(N__39902));
    InMux I__9689 (
            .O(N__39906),
            .I(N__39899));
    InMux I__9688 (
            .O(N__39905),
            .I(N__39894));
    Span4Mux_v I__9687 (
            .O(N__39902),
            .I(N__39889));
    LocalMux I__9686 (
            .O(N__39899),
            .I(N__39889));
    CascadeMux I__9685 (
            .O(N__39898),
            .I(N__39886));
    CascadeMux I__9684 (
            .O(N__39897),
            .I(N__39883));
    LocalMux I__9683 (
            .O(N__39894),
            .I(N__39880));
    Span4Mux_h I__9682 (
            .O(N__39889),
            .I(N__39877));
    InMux I__9681 (
            .O(N__39886),
            .I(N__39874));
    InMux I__9680 (
            .O(N__39883),
            .I(N__39871));
    Span4Mux_h I__9679 (
            .O(N__39880),
            .I(N__39867));
    Span4Mux_h I__9678 (
            .O(N__39877),
            .I(N__39860));
    LocalMux I__9677 (
            .O(N__39874),
            .I(N__39860));
    LocalMux I__9676 (
            .O(N__39871),
            .I(N__39860));
    InMux I__9675 (
            .O(N__39870),
            .I(N__39857));
    Span4Mux_v I__9674 (
            .O(N__39867),
            .I(N__39853));
    Span4Mux_v I__9673 (
            .O(N__39860),
            .I(N__39850));
    LocalMux I__9672 (
            .O(N__39857),
            .I(N__39847));
    InMux I__9671 (
            .O(N__39856),
            .I(N__39844));
    Span4Mux_v I__9670 (
            .O(N__39853),
            .I(N__39839));
    Span4Mux_h I__9669 (
            .O(N__39850),
            .I(N__39839));
    Span12Mux_s10_v I__9668 (
            .O(N__39847),
            .I(N__39835));
    LocalMux I__9667 (
            .O(N__39844),
            .I(N__39832));
    Sp12to4 I__9666 (
            .O(N__39839),
            .I(N__39829));
    InMux I__9665 (
            .O(N__39838),
            .I(N__39826));
    Span12Mux_v I__9664 (
            .O(N__39835),
            .I(N__39823));
    Span12Mux_h I__9663 (
            .O(N__39832),
            .I(N__39816));
    Span12Mux_s6_h I__9662 (
            .O(N__39829),
            .I(N__39816));
    LocalMux I__9661 (
            .O(N__39826),
            .I(N__39816));
    Span12Mux_h I__9660 (
            .O(N__39823),
            .I(N__39813));
    Span12Mux_v I__9659 (
            .O(N__39816),
            .I(N__39810));
    Odrv12 I__9658 (
            .O(N__39813),
            .I(port_data_in_7));
    Odrv12 I__9657 (
            .O(N__39810),
            .I(port_data_in_7));
    InMux I__9656 (
            .O(N__39805),
            .I(un1_M_this_map_address_q_cry_5));
    InMux I__9655 (
            .O(N__39802),
            .I(un1_M_this_map_address_q_cry_6));
    InMux I__9654 (
            .O(N__39799),
            .I(bfn_24_24_0_));
    InMux I__9653 (
            .O(N__39796),
            .I(un1_M_this_map_address_q_cry_8));
    InMux I__9652 (
            .O(N__39793),
            .I(N__39790));
    LocalMux I__9651 (
            .O(N__39790),
            .I(N__39787));
    Odrv4 I__9650 (
            .O(N__39787),
            .I(un1_M_this_map_address_q_cry_5_THRU_CO));
    InMux I__9649 (
            .O(N__39784),
            .I(N__39778));
    InMux I__9648 (
            .O(N__39783),
            .I(N__39774));
    InMux I__9647 (
            .O(N__39782),
            .I(N__39771));
    InMux I__9646 (
            .O(N__39781),
            .I(N__39768));
    LocalMux I__9645 (
            .O(N__39778),
            .I(N__39765));
    InMux I__9644 (
            .O(N__39777),
            .I(N__39762));
    LocalMux I__9643 (
            .O(N__39774),
            .I(N__39757));
    LocalMux I__9642 (
            .O(N__39771),
            .I(N__39754));
    LocalMux I__9641 (
            .O(N__39768),
            .I(N__39750));
    Span4Mux_v I__9640 (
            .O(N__39765),
            .I(N__39745));
    LocalMux I__9639 (
            .O(N__39762),
            .I(N__39745));
    InMux I__9638 (
            .O(N__39761),
            .I(N__39742));
    InMux I__9637 (
            .O(N__39760),
            .I(N__39739));
    Span4Mux_h I__9636 (
            .O(N__39757),
            .I(N__39736));
    Span4Mux_h I__9635 (
            .O(N__39754),
            .I(N__39733));
    InMux I__9634 (
            .O(N__39753),
            .I(N__39730));
    Span4Mux_v I__9633 (
            .O(N__39750),
            .I(N__39725));
    Span4Mux_v I__9632 (
            .O(N__39745),
            .I(N__39720));
    LocalMux I__9631 (
            .O(N__39742),
            .I(N__39720));
    LocalMux I__9630 (
            .O(N__39739),
            .I(N__39717));
    Span4Mux_h I__9629 (
            .O(N__39736),
            .I(N__39710));
    Span4Mux_v I__9628 (
            .O(N__39733),
            .I(N__39710));
    LocalMux I__9627 (
            .O(N__39730),
            .I(N__39710));
    InMux I__9626 (
            .O(N__39729),
            .I(N__39707));
    InMux I__9625 (
            .O(N__39728),
            .I(N__39704));
    Span4Mux_v I__9624 (
            .O(N__39725),
            .I(N__39701));
    Span4Mux_v I__9623 (
            .O(N__39720),
            .I(N__39698));
    Span4Mux_v I__9622 (
            .O(N__39717),
            .I(N__39695));
    Span4Mux_h I__9621 (
            .O(N__39710),
            .I(N__39690));
    LocalMux I__9620 (
            .O(N__39707),
            .I(N__39690));
    LocalMux I__9619 (
            .O(N__39704),
            .I(N__39687));
    Sp12to4 I__9618 (
            .O(N__39701),
            .I(N__39681));
    Sp12to4 I__9617 (
            .O(N__39698),
            .I(N__39681));
    Span4Mux_v I__9616 (
            .O(N__39695),
            .I(N__39678));
    Span4Mux_v I__9615 (
            .O(N__39690),
            .I(N__39673));
    Span4Mux_h I__9614 (
            .O(N__39687),
            .I(N__39673));
    InMux I__9613 (
            .O(N__39686),
            .I(N__39670));
    Span12Mux_h I__9612 (
            .O(N__39681),
            .I(N__39667));
    IoSpan4Mux I__9611 (
            .O(N__39678),
            .I(N__39664));
    Span4Mux_v I__9610 (
            .O(N__39673),
            .I(N__39661));
    LocalMux I__9609 (
            .O(N__39670),
            .I(N__39658));
    Odrv12 I__9608 (
            .O(N__39667),
            .I(port_data_in_1));
    Odrv4 I__9607 (
            .O(N__39664),
            .I(port_data_in_1));
    Odrv4 I__9606 (
            .O(N__39661),
            .I(port_data_in_1));
    Odrv12 I__9605 (
            .O(N__39658),
            .I(port_data_in_1));
    CascadeMux I__9604 (
            .O(N__39649),
            .I(M_this_map_address_qc_8_1_cascade_));
    CascadeMux I__9603 (
            .O(N__39646),
            .I(N__39643));
    CascadeBuf I__9602 (
            .O(N__39643),
            .I(N__39640));
    CascadeMux I__9601 (
            .O(N__39640),
            .I(N__39637));
    InMux I__9600 (
            .O(N__39637),
            .I(N__39634));
    LocalMux I__9599 (
            .O(N__39634),
            .I(N__39629));
    CascadeMux I__9598 (
            .O(N__39633),
            .I(N__39626));
    InMux I__9597 (
            .O(N__39632),
            .I(N__39623));
    Span4Mux_s1_v I__9596 (
            .O(N__39629),
            .I(N__39620));
    InMux I__9595 (
            .O(N__39626),
            .I(N__39617));
    LocalMux I__9594 (
            .O(N__39623),
            .I(N__39614));
    Span4Mux_v I__9593 (
            .O(N__39620),
            .I(N__39611));
    LocalMux I__9592 (
            .O(N__39617),
            .I(M_this_map_address_qZ0Z_6));
    Odrv4 I__9591 (
            .O(N__39614),
            .I(M_this_map_address_qZ0Z_6));
    Odrv4 I__9590 (
            .O(N__39611),
            .I(M_this_map_address_qZ0Z_6));
    InMux I__9589 (
            .O(N__39604),
            .I(N__39601));
    LocalMux I__9588 (
            .O(N__39601),
            .I(un1_M_this_map_address_q_cry_7_THRU_CO));
    InMux I__9587 (
            .O(N__39598),
            .I(N__39595));
    LocalMux I__9586 (
            .O(N__39595),
            .I(N__39592));
    Odrv4 I__9585 (
            .O(N__39592),
            .I(un1_M_this_map_address_q_axb_0));
    InMux I__9584 (
            .O(N__39589),
            .I(N__39586));
    LocalMux I__9583 (
            .O(N__39586),
            .I(M_this_map_address_qc_2_0));
    CascadeMux I__9582 (
            .O(N__39583),
            .I(N__39580));
    InMux I__9581 (
            .O(N__39580),
            .I(N__39577));
    LocalMux I__9580 (
            .O(N__39577),
            .I(N_1097));
    CascadeMux I__9579 (
            .O(N__39574),
            .I(N__39571));
    CascadeBuf I__9578 (
            .O(N__39571),
            .I(N__39568));
    CascadeMux I__9577 (
            .O(N__39568),
            .I(N__39565));
    InMux I__9576 (
            .O(N__39565),
            .I(N__39559));
    CascadeMux I__9575 (
            .O(N__39564),
            .I(N__39556));
    InMux I__9574 (
            .O(N__39563),
            .I(N__39551));
    InMux I__9573 (
            .O(N__39562),
            .I(N__39551));
    LocalMux I__9572 (
            .O(N__39559),
            .I(N__39548));
    InMux I__9571 (
            .O(N__39556),
            .I(N__39544));
    LocalMux I__9570 (
            .O(N__39551),
            .I(N__39541));
    Span4Mux_s1_v I__9569 (
            .O(N__39548),
            .I(N__39538));
    InMux I__9568 (
            .O(N__39547),
            .I(N__39535));
    LocalMux I__9567 (
            .O(N__39544),
            .I(N__39532));
    Span4Mux_h I__9566 (
            .O(N__39541),
            .I(N__39527));
    Span4Mux_v I__9565 (
            .O(N__39538),
            .I(N__39527));
    LocalMux I__9564 (
            .O(N__39535),
            .I(M_this_map_address_qZ0Z_0));
    Odrv4 I__9563 (
            .O(N__39532),
            .I(M_this_map_address_qZ0Z_0));
    Odrv4 I__9562 (
            .O(N__39527),
            .I(M_this_map_address_qZ0Z_0));
    InMux I__9561 (
            .O(N__39520),
            .I(N__39517));
    LocalMux I__9560 (
            .O(N__39517),
            .I(N__39514));
    Span4Mux_s2_v I__9559 (
            .O(N__39514),
            .I(N__39511));
    Odrv4 I__9558 (
            .O(N__39511),
            .I(N_921_0));
    InMux I__9557 (
            .O(N__39508),
            .I(N__39502));
    CascadeMux I__9556 (
            .O(N__39507),
            .I(N__39499));
    InMux I__9555 (
            .O(N__39506),
            .I(N__39496));
    InMux I__9554 (
            .O(N__39505),
            .I(N__39493));
    LocalMux I__9553 (
            .O(N__39502),
            .I(N__39489));
    InMux I__9552 (
            .O(N__39499),
            .I(N__39486));
    LocalMux I__9551 (
            .O(N__39496),
            .I(N__39482));
    LocalMux I__9550 (
            .O(N__39493),
            .I(N__39479));
    InMux I__9549 (
            .O(N__39492),
            .I(N__39476));
    Span4Mux_h I__9548 (
            .O(N__39489),
            .I(N__39473));
    LocalMux I__9547 (
            .O(N__39486),
            .I(N__39470));
    InMux I__9546 (
            .O(N__39485),
            .I(N__39467));
    Span4Mux_v I__9545 (
            .O(N__39482),
            .I(N__39462));
    Span4Mux_v I__9544 (
            .O(N__39479),
            .I(N__39462));
    LocalMux I__9543 (
            .O(N__39476),
            .I(N__39456));
    Span4Mux_v I__9542 (
            .O(N__39473),
            .I(N__39449));
    Span4Mux_h I__9541 (
            .O(N__39470),
            .I(N__39449));
    LocalMux I__9540 (
            .O(N__39467),
            .I(N__39449));
    Sp12to4 I__9539 (
            .O(N__39462),
            .I(N__39446));
    InMux I__9538 (
            .O(N__39461),
            .I(N__39443));
    InMux I__9537 (
            .O(N__39460),
            .I(N__39440));
    InMux I__9536 (
            .O(N__39459),
            .I(N__39437));
    Span4Mux_h I__9535 (
            .O(N__39456),
            .I(N__39434));
    Span4Mux_h I__9534 (
            .O(N__39449),
            .I(N__39431));
    Span12Mux_h I__9533 (
            .O(N__39446),
            .I(N__39422));
    LocalMux I__9532 (
            .O(N__39443),
            .I(N__39422));
    LocalMux I__9531 (
            .O(N__39440),
            .I(N__39422));
    LocalMux I__9530 (
            .O(N__39437),
            .I(N__39422));
    Odrv4 I__9529 (
            .O(N__39434),
            .I(N_842_0));
    Odrv4 I__9528 (
            .O(N__39431),
            .I(N_842_0));
    Odrv12 I__9527 (
            .O(N__39422),
            .I(N_842_0));
    InMux I__9526 (
            .O(N__39415),
            .I(N__39412));
    LocalMux I__9525 (
            .O(N__39412),
            .I(N__39409));
    Odrv12 I__9524 (
            .O(N__39409),
            .I(M_this_status_flags_qZ0Z_7));
    InMux I__9523 (
            .O(N__39406),
            .I(N__39403));
    LocalMux I__9522 (
            .O(N__39403),
            .I(N__39400));
    Span4Mux_h I__9521 (
            .O(N__39400),
            .I(N__39397));
    Odrv4 I__9520 (
            .O(N__39397),
            .I(M_this_map_address_qc_3_1));
    InMux I__9519 (
            .O(N__39394),
            .I(N__39391));
    LocalMux I__9518 (
            .O(N__39391),
            .I(un1_M_this_map_address_q_cry_0_c_RNOZ0));
    CascadeMux I__9517 (
            .O(N__39388),
            .I(N__39385));
    CascadeBuf I__9516 (
            .O(N__39385),
            .I(N__39382));
    CascadeMux I__9515 (
            .O(N__39382),
            .I(N__39378));
    InMux I__9514 (
            .O(N__39381),
            .I(N__39374));
    InMux I__9513 (
            .O(N__39378),
            .I(N__39371));
    CascadeMux I__9512 (
            .O(N__39377),
            .I(N__39368));
    LocalMux I__9511 (
            .O(N__39374),
            .I(N__39365));
    LocalMux I__9510 (
            .O(N__39371),
            .I(N__39361));
    InMux I__9509 (
            .O(N__39368),
            .I(N__39358));
    Span4Mux_h I__9508 (
            .O(N__39365),
            .I(N__39355));
    InMux I__9507 (
            .O(N__39364),
            .I(N__39352));
    Span12Mux_s10_v I__9506 (
            .O(N__39361),
            .I(N__39349));
    LocalMux I__9505 (
            .O(N__39358),
            .I(M_this_map_address_qZ0Z_1));
    Odrv4 I__9504 (
            .O(N__39355),
            .I(M_this_map_address_qZ0Z_1));
    LocalMux I__9503 (
            .O(N__39352),
            .I(M_this_map_address_qZ0Z_1));
    Odrv12 I__9502 (
            .O(N__39349),
            .I(M_this_map_address_qZ0Z_1));
    InMux I__9501 (
            .O(N__39340),
            .I(N__39337));
    LocalMux I__9500 (
            .O(N__39337),
            .I(un1_M_this_map_address_q_cry_0_THRU_CO));
    InMux I__9499 (
            .O(N__39334),
            .I(un1_M_this_map_address_q_cry_0));
    CascadeMux I__9498 (
            .O(N__39331),
            .I(N__39328));
    CascadeBuf I__9497 (
            .O(N__39328),
            .I(N__39325));
    CascadeMux I__9496 (
            .O(N__39325),
            .I(N__39322));
    InMux I__9495 (
            .O(N__39322),
            .I(N__39319));
    LocalMux I__9494 (
            .O(N__39319),
            .I(N__39314));
    InMux I__9493 (
            .O(N__39318),
            .I(N__39311));
    InMux I__9492 (
            .O(N__39317),
            .I(N__39308));
    Span12Mux_s9_h I__9491 (
            .O(N__39314),
            .I(N__39305));
    LocalMux I__9490 (
            .O(N__39311),
            .I(M_this_map_address_qZ0Z_2));
    LocalMux I__9489 (
            .O(N__39308),
            .I(M_this_map_address_qZ0Z_2));
    Odrv12 I__9488 (
            .O(N__39305),
            .I(M_this_map_address_qZ0Z_2));
    InMux I__9487 (
            .O(N__39298),
            .I(N__39295));
    LocalMux I__9486 (
            .O(N__39295),
            .I(M_this_map_address_q_RNO_1Z0Z_2));
    InMux I__9485 (
            .O(N__39292),
            .I(un1_M_this_map_address_q_cry_1));
    CascadeMux I__9484 (
            .O(N__39289),
            .I(N__39286));
    CascadeBuf I__9483 (
            .O(N__39286),
            .I(N__39283));
    CascadeMux I__9482 (
            .O(N__39283),
            .I(N__39280));
    InMux I__9481 (
            .O(N__39280),
            .I(N__39277));
    LocalMux I__9480 (
            .O(N__39277),
            .I(N__39274));
    Span4Mux_v I__9479 (
            .O(N__39274),
            .I(N__39269));
    InMux I__9478 (
            .O(N__39273),
            .I(N__39266));
    InMux I__9477 (
            .O(N__39272),
            .I(N__39263));
    Span4Mux_v I__9476 (
            .O(N__39269),
            .I(N__39260));
    LocalMux I__9475 (
            .O(N__39266),
            .I(M_this_map_address_qZ0Z_3));
    LocalMux I__9474 (
            .O(N__39263),
            .I(M_this_map_address_qZ0Z_3));
    Odrv4 I__9473 (
            .O(N__39260),
            .I(M_this_map_address_qZ0Z_3));
    InMux I__9472 (
            .O(N__39253),
            .I(N__39250));
    LocalMux I__9471 (
            .O(N__39250),
            .I(M_this_map_address_q_RNO_1Z0Z_3));
    InMux I__9470 (
            .O(N__39247),
            .I(un1_M_this_map_address_q_cry_2));
    CascadeMux I__9469 (
            .O(N__39244),
            .I(N__39241));
    CascadeBuf I__9468 (
            .O(N__39241),
            .I(N__39238));
    CascadeMux I__9467 (
            .O(N__39238),
            .I(N__39235));
    InMux I__9466 (
            .O(N__39235),
            .I(N__39232));
    LocalMux I__9465 (
            .O(N__39232),
            .I(N__39229));
    Span4Mux_v I__9464 (
            .O(N__39229),
            .I(N__39224));
    InMux I__9463 (
            .O(N__39228),
            .I(N__39221));
    InMux I__9462 (
            .O(N__39227),
            .I(N__39218));
    Span4Mux_v I__9461 (
            .O(N__39224),
            .I(N__39215));
    LocalMux I__9460 (
            .O(N__39221),
            .I(M_this_map_address_qZ0Z_4));
    LocalMux I__9459 (
            .O(N__39218),
            .I(M_this_map_address_qZ0Z_4));
    Odrv4 I__9458 (
            .O(N__39215),
            .I(M_this_map_address_qZ0Z_4));
    InMux I__9457 (
            .O(N__39208),
            .I(N__39205));
    LocalMux I__9456 (
            .O(N__39205),
            .I(M_this_map_address_q_RNO_1Z0Z_4));
    InMux I__9455 (
            .O(N__39202),
            .I(un1_M_this_map_address_q_cry_3));
    InMux I__9454 (
            .O(N__39199),
            .I(N__39195));
    InMux I__9453 (
            .O(N__39198),
            .I(N__39192));
    LocalMux I__9452 (
            .O(N__39195),
            .I(un1_M_this_state_q_7_i_0_a3_0_0));
    LocalMux I__9451 (
            .O(N__39192),
            .I(un1_M_this_state_q_7_i_0_a3_0_0));
    InMux I__9450 (
            .O(N__39187),
            .I(un1_M_this_map_address_q_cry_4));
    CEMux I__9449 (
            .O(N__39184),
            .I(N__39181));
    LocalMux I__9448 (
            .O(N__39181),
            .I(N__39177));
    CEMux I__9447 (
            .O(N__39180),
            .I(N__39174));
    Span4Mux_h I__9446 (
            .O(N__39177),
            .I(N__39169));
    LocalMux I__9445 (
            .O(N__39174),
            .I(N__39169));
    Span4Mux_v I__9444 (
            .O(N__39169),
            .I(N__39166));
    Odrv4 I__9443 (
            .O(N__39166),
            .I(\this_spr_ram.mem_WE_10 ));
    InMux I__9442 (
            .O(N__39163),
            .I(N__39160));
    LocalMux I__9441 (
            .O(N__39160),
            .I(N__39157));
    Odrv4 I__9440 (
            .O(N__39157),
            .I(\this_spr_ram.mem_out_bus4_0 ));
    InMux I__9439 (
            .O(N__39154),
            .I(N__39151));
    LocalMux I__9438 (
            .O(N__39151),
            .I(N__39148));
    Sp12to4 I__9437 (
            .O(N__39148),
            .I(N__39145));
    Span12Mux_v I__9436 (
            .O(N__39145),
            .I(N__39142));
    Odrv12 I__9435 (
            .O(N__39142),
            .I(\this_spr_ram.mem_out_bus0_0 ));
    InMux I__9434 (
            .O(N__39139),
            .I(N__39136));
    LocalMux I__9433 (
            .O(N__39136),
            .I(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0 ));
    InMux I__9432 (
            .O(N__39133),
            .I(N__39130));
    LocalMux I__9431 (
            .O(N__39130),
            .I(N__39127));
    Span4Mux_v I__9430 (
            .O(N__39127),
            .I(N__39124));
    Odrv4 I__9429 (
            .O(N__39124),
            .I(\this_spr_ram.mem_out_bus2_1 ));
    InMux I__9428 (
            .O(N__39121),
            .I(N__39118));
    LocalMux I__9427 (
            .O(N__39118),
            .I(N__39114));
    InMux I__9426 (
            .O(N__39117),
            .I(N__39101));
    Span4Mux_v I__9425 (
            .O(N__39114),
            .I(N__39094));
    InMux I__9424 (
            .O(N__39113),
            .I(N__39081));
    InMux I__9423 (
            .O(N__39112),
            .I(N__39081));
    InMux I__9422 (
            .O(N__39111),
            .I(N__39081));
    InMux I__9421 (
            .O(N__39110),
            .I(N__39081));
    InMux I__9420 (
            .O(N__39109),
            .I(N__39081));
    InMux I__9419 (
            .O(N__39108),
            .I(N__39081));
    InMux I__9418 (
            .O(N__39107),
            .I(N__39076));
    InMux I__9417 (
            .O(N__39106),
            .I(N__39076));
    InMux I__9416 (
            .O(N__39105),
            .I(N__39073));
    InMux I__9415 (
            .O(N__39104),
            .I(N__39070));
    LocalMux I__9414 (
            .O(N__39101),
            .I(N__39067));
    InMux I__9413 (
            .O(N__39100),
            .I(N__39062));
    InMux I__9412 (
            .O(N__39099),
            .I(N__39062));
    InMux I__9411 (
            .O(N__39098),
            .I(N__39059));
    InMux I__9410 (
            .O(N__39097),
            .I(N__39056));
    Span4Mux_v I__9409 (
            .O(N__39094),
            .I(N__39051));
    LocalMux I__9408 (
            .O(N__39081),
            .I(N__39051));
    LocalMux I__9407 (
            .O(N__39076),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    LocalMux I__9406 (
            .O(N__39073),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    LocalMux I__9405 (
            .O(N__39070),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    Odrv4 I__9404 (
            .O(N__39067),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    LocalMux I__9403 (
            .O(N__39062),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    LocalMux I__9402 (
            .O(N__39059),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    LocalMux I__9401 (
            .O(N__39056),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    Odrv4 I__9400 (
            .O(N__39051),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    InMux I__9399 (
            .O(N__39034),
            .I(N__39031));
    LocalMux I__9398 (
            .O(N__39031),
            .I(N__39028));
    Span4Mux_v I__9397 (
            .O(N__39028),
            .I(N__39025));
    Span4Mux_v I__9396 (
            .O(N__39025),
            .I(N__39022));
    Odrv4 I__9395 (
            .O(N__39022),
            .I(\this_spr_ram.mem_out_bus6_1 ));
    InMux I__9394 (
            .O(N__39019),
            .I(N__39016));
    LocalMux I__9393 (
            .O(N__39016),
            .I(N__39013));
    Odrv4 I__9392 (
            .O(N__39013),
            .I(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0 ));
    InMux I__9391 (
            .O(N__39010),
            .I(N__39007));
    LocalMux I__9390 (
            .O(N__39007),
            .I(N__39003));
    InMux I__9389 (
            .O(N__39006),
            .I(N__39000));
    Span4Mux_v I__9388 (
            .O(N__39003),
            .I(N__38995));
    LocalMux I__9387 (
            .O(N__39000),
            .I(N__38995));
    Span4Mux_h I__9386 (
            .O(N__38995),
            .I(N__38992));
    Sp12to4 I__9385 (
            .O(N__38992),
            .I(N__38989));
    Span12Mux_v I__9384 (
            .O(N__38989),
            .I(N__38986));
    Odrv12 I__9383 (
            .O(N__38986),
            .I(M_this_map_ram_read_data_7));
    IoInMux I__9382 (
            .O(N__38983),
            .I(N__38980));
    LocalMux I__9381 (
            .O(N__38980),
            .I(N__38977));
    IoSpan4Mux I__9380 (
            .O(N__38977),
            .I(N__38974));
    IoSpan4Mux I__9379 (
            .O(N__38974),
            .I(N__38971));
    Span4Mux_s3_h I__9378 (
            .O(N__38971),
            .I(N__38968));
    Span4Mux_h I__9377 (
            .O(N__38968),
            .I(N__38965));
    Odrv4 I__9376 (
            .O(N__38965),
            .I(IO_port_data_write_i_m2_i_m2_7));
    CEMux I__9375 (
            .O(N__38962),
            .I(N__38958));
    CEMux I__9374 (
            .O(N__38961),
            .I(N__38955));
    LocalMux I__9373 (
            .O(N__38958),
            .I(N__38950));
    LocalMux I__9372 (
            .O(N__38955),
            .I(N__38950));
    Span4Mux_v I__9371 (
            .O(N__38950),
            .I(N__38947));
    Odrv4 I__9370 (
            .O(N__38947),
            .I(\this_spr_ram.mem_WE_6 ));
    CEMux I__9369 (
            .O(N__38944),
            .I(N__38940));
    CEMux I__9368 (
            .O(N__38943),
            .I(N__38937));
    LocalMux I__9367 (
            .O(N__38940),
            .I(N__38932));
    LocalMux I__9366 (
            .O(N__38937),
            .I(N__38932));
    Span4Mux_v I__9365 (
            .O(N__38932),
            .I(N__38929));
    Odrv4 I__9364 (
            .O(N__38929),
            .I(\this_spr_ram.mem_WE_4 ));
    InMux I__9363 (
            .O(N__38926),
            .I(N__38914));
    InMux I__9362 (
            .O(N__38925),
            .I(N__38914));
    InMux I__9361 (
            .O(N__38924),
            .I(N__38914));
    InMux I__9360 (
            .O(N__38923),
            .I(N__38911));
    InMux I__9359 (
            .O(N__38922),
            .I(N__38908));
    InMux I__9358 (
            .O(N__38921),
            .I(N__38905));
    LocalMux I__9357 (
            .O(N__38914),
            .I(N__38895));
    LocalMux I__9356 (
            .O(N__38911),
            .I(N__38895));
    LocalMux I__9355 (
            .O(N__38908),
            .I(N__38895));
    LocalMux I__9354 (
            .O(N__38905),
            .I(N__38892));
    InMux I__9353 (
            .O(N__38904),
            .I(N__38887));
    InMux I__9352 (
            .O(N__38903),
            .I(N__38887));
    InMux I__9351 (
            .O(N__38902),
            .I(N__38884));
    Span4Mux_v I__9350 (
            .O(N__38895),
            .I(N__38881));
    Span4Mux_h I__9349 (
            .O(N__38892),
            .I(N__38878));
    LocalMux I__9348 (
            .O(N__38887),
            .I(N__38875));
    LocalMux I__9347 (
            .O(N__38884),
            .I(M_this_spr_address_qZ0Z_12));
    Odrv4 I__9346 (
            .O(N__38881),
            .I(M_this_spr_address_qZ0Z_12));
    Odrv4 I__9345 (
            .O(N__38878),
            .I(M_this_spr_address_qZ0Z_12));
    Odrv12 I__9344 (
            .O(N__38875),
            .I(M_this_spr_address_qZ0Z_12));
    CascadeMux I__9343 (
            .O(N__38866),
            .I(N__38862));
    InMux I__9342 (
            .O(N__38865),
            .I(N__38855));
    InMux I__9341 (
            .O(N__38862),
            .I(N__38848));
    InMux I__9340 (
            .O(N__38861),
            .I(N__38848));
    InMux I__9339 (
            .O(N__38860),
            .I(N__38848));
    InMux I__9338 (
            .O(N__38859),
            .I(N__38843));
    CascadeMux I__9337 (
            .O(N__38858),
            .I(N__38840));
    LocalMux I__9336 (
            .O(N__38855),
            .I(N__38836));
    LocalMux I__9335 (
            .O(N__38848),
            .I(N__38833));
    InMux I__9334 (
            .O(N__38847),
            .I(N__38830));
    InMux I__9333 (
            .O(N__38846),
            .I(N__38827));
    LocalMux I__9332 (
            .O(N__38843),
            .I(N__38824));
    InMux I__9331 (
            .O(N__38840),
            .I(N__38819));
    InMux I__9330 (
            .O(N__38839),
            .I(N__38819));
    Span4Mux_v I__9329 (
            .O(N__38836),
            .I(N__38814));
    Span4Mux_v I__9328 (
            .O(N__38833),
            .I(N__38814));
    LocalMux I__9327 (
            .O(N__38830),
            .I(N__38811));
    LocalMux I__9326 (
            .O(N__38827),
            .I(N__38802));
    Span4Mux_v I__9325 (
            .O(N__38824),
            .I(N__38802));
    LocalMux I__9324 (
            .O(N__38819),
            .I(N__38802));
    Span4Mux_h I__9323 (
            .O(N__38814),
            .I(N__38802));
    Odrv4 I__9322 (
            .O(N__38811),
            .I(M_this_spr_address_qZ0Z_11));
    Odrv4 I__9321 (
            .O(N__38802),
            .I(M_this_spr_address_qZ0Z_11));
    CascadeMux I__9320 (
            .O(N__38797),
            .I(N__38790));
    CascadeMux I__9319 (
            .O(N__38796),
            .I(N__38786));
    CascadeMux I__9318 (
            .O(N__38795),
            .I(N__38783));
    CascadeMux I__9317 (
            .O(N__38794),
            .I(N__38780));
    CascadeMux I__9316 (
            .O(N__38793),
            .I(N__38777));
    InMux I__9315 (
            .O(N__38790),
            .I(N__38769));
    InMux I__9314 (
            .O(N__38789),
            .I(N__38769));
    InMux I__9313 (
            .O(N__38786),
            .I(N__38769));
    InMux I__9312 (
            .O(N__38783),
            .I(N__38766));
    InMux I__9311 (
            .O(N__38780),
            .I(N__38763));
    InMux I__9310 (
            .O(N__38777),
            .I(N__38760));
    CascadeMux I__9309 (
            .O(N__38776),
            .I(N__38756));
    LocalMux I__9308 (
            .O(N__38769),
            .I(N__38748));
    LocalMux I__9307 (
            .O(N__38766),
            .I(N__38748));
    LocalMux I__9306 (
            .O(N__38763),
            .I(N__38748));
    LocalMux I__9305 (
            .O(N__38760),
            .I(N__38745));
    InMux I__9304 (
            .O(N__38759),
            .I(N__38740));
    InMux I__9303 (
            .O(N__38756),
            .I(N__38740));
    InMux I__9302 (
            .O(N__38755),
            .I(N__38737));
    Span4Mux_v I__9301 (
            .O(N__38748),
            .I(N__38734));
    Span4Mux_h I__9300 (
            .O(N__38745),
            .I(N__38731));
    LocalMux I__9299 (
            .O(N__38740),
            .I(N__38728));
    LocalMux I__9298 (
            .O(N__38737),
            .I(M_this_spr_address_qZ0Z_13));
    Odrv4 I__9297 (
            .O(N__38734),
            .I(M_this_spr_address_qZ0Z_13));
    Odrv4 I__9296 (
            .O(N__38731),
            .I(M_this_spr_address_qZ0Z_13));
    Odrv4 I__9295 (
            .O(N__38728),
            .I(M_this_spr_address_qZ0Z_13));
    InMux I__9294 (
            .O(N__38719),
            .I(N__38713));
    InMux I__9293 (
            .O(N__38718),
            .I(N__38710));
    InMux I__9292 (
            .O(N__38717),
            .I(N__38704));
    InMux I__9291 (
            .O(N__38716),
            .I(N__38704));
    LocalMux I__9290 (
            .O(N__38713),
            .I(N__38698));
    LocalMux I__9289 (
            .O(N__38710),
            .I(N__38695));
    InMux I__9288 (
            .O(N__38709),
            .I(N__38692));
    LocalMux I__9287 (
            .O(N__38704),
            .I(N__38689));
    InMux I__9286 (
            .O(N__38703),
            .I(N__38682));
    InMux I__9285 (
            .O(N__38702),
            .I(N__38682));
    InMux I__9284 (
            .O(N__38701),
            .I(N__38682));
    Span4Mux_h I__9283 (
            .O(N__38698),
            .I(N__38679));
    Span4Mux_h I__9282 (
            .O(N__38695),
            .I(N__38674));
    LocalMux I__9281 (
            .O(N__38692),
            .I(N__38674));
    Span4Mux_h I__9280 (
            .O(N__38689),
            .I(N__38671));
    LocalMux I__9279 (
            .O(N__38682),
            .I(N__38668));
    Span4Mux_v I__9278 (
            .O(N__38679),
            .I(N__38665));
    Span4Mux_v I__9277 (
            .O(N__38674),
            .I(N__38662));
    Span4Mux_v I__9276 (
            .O(N__38671),
            .I(N__38657));
    Span4Mux_h I__9275 (
            .O(N__38668),
            .I(N__38657));
    Odrv4 I__9274 (
            .O(N__38665),
            .I(M_this_spr_ram_write_en_0_i_1_0_0));
    Odrv4 I__9273 (
            .O(N__38662),
            .I(M_this_spr_ram_write_en_0_i_1_0_0));
    Odrv4 I__9272 (
            .O(N__38657),
            .I(M_this_spr_ram_write_en_0_i_1_0_0));
    CEMux I__9271 (
            .O(N__38650),
            .I(N__38647));
    LocalMux I__9270 (
            .O(N__38647),
            .I(N__38643));
    CEMux I__9269 (
            .O(N__38646),
            .I(N__38640));
    Sp12to4 I__9268 (
            .O(N__38643),
            .I(N__38637));
    LocalMux I__9267 (
            .O(N__38640),
            .I(N__38634));
    Span12Mux_v I__9266 (
            .O(N__38637),
            .I(N__38631));
    Span4Mux_v I__9265 (
            .O(N__38634),
            .I(N__38628));
    Span12Mux_h I__9264 (
            .O(N__38631),
            .I(N__38625));
    Span4Mux_v I__9263 (
            .O(N__38628),
            .I(N__38622));
    Odrv12 I__9262 (
            .O(N__38625),
            .I(\this_spr_ram.mem_WE_2 ));
    Odrv4 I__9261 (
            .O(N__38622),
            .I(\this_spr_ram.mem_WE_2 ));
    InMux I__9260 (
            .O(N__38617),
            .I(N__38614));
    LocalMux I__9259 (
            .O(N__38614),
            .I(N_1066));
    CascadeMux I__9258 (
            .O(N__38611),
            .I(M_this_map_address_qc_6_0_cascade_));
    InMux I__9257 (
            .O(N__38608),
            .I(N__38602));
    InMux I__9256 (
            .O(N__38607),
            .I(N__38599));
    InMux I__9255 (
            .O(N__38606),
            .I(N__38592));
    InMux I__9254 (
            .O(N__38605),
            .I(N__38589));
    LocalMux I__9253 (
            .O(N__38602),
            .I(N__38581));
    LocalMux I__9252 (
            .O(N__38599),
            .I(N__38581));
    InMux I__9251 (
            .O(N__38598),
            .I(N__38578));
    InMux I__9250 (
            .O(N__38597),
            .I(N__38571));
    InMux I__9249 (
            .O(N__38596),
            .I(N__38571));
    InMux I__9248 (
            .O(N__38595),
            .I(N__38571));
    LocalMux I__9247 (
            .O(N__38592),
            .I(N__38566));
    LocalMux I__9246 (
            .O(N__38589),
            .I(N__38566));
    InMux I__9245 (
            .O(N__38588),
            .I(N__38563));
    InMux I__9244 (
            .O(N__38587),
            .I(N__38560));
    InMux I__9243 (
            .O(N__38586),
            .I(N__38557));
    Span4Mux_v I__9242 (
            .O(N__38581),
            .I(N__38550));
    LocalMux I__9241 (
            .O(N__38578),
            .I(N__38550));
    LocalMux I__9240 (
            .O(N__38571),
            .I(N__38550));
    Span4Mux_v I__9239 (
            .O(N__38566),
            .I(N__38545));
    LocalMux I__9238 (
            .O(N__38563),
            .I(N__38545));
    LocalMux I__9237 (
            .O(N__38560),
            .I(M_this_state_qZ0Z_4));
    LocalMux I__9236 (
            .O(N__38557),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__9235 (
            .O(N__38550),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__9234 (
            .O(N__38545),
            .I(M_this_state_qZ0Z_4));
    InMux I__9233 (
            .O(N__38536),
            .I(N__38527));
    InMux I__9232 (
            .O(N__38535),
            .I(N__38527));
    InMux I__9231 (
            .O(N__38534),
            .I(N__38524));
    InMux I__9230 (
            .O(N__38533),
            .I(N__38519));
    InMux I__9229 (
            .O(N__38532),
            .I(N__38519));
    LocalMux I__9228 (
            .O(N__38527),
            .I(N__38514));
    LocalMux I__9227 (
            .O(N__38524),
            .I(N__38514));
    LocalMux I__9226 (
            .O(N__38519),
            .I(N__38511));
    Span4Mux_h I__9225 (
            .O(N__38514),
            .I(N__38508));
    Odrv12 I__9224 (
            .O(N__38511),
            .I(N_794_0));
    Odrv4 I__9223 (
            .O(N__38508),
            .I(N_794_0));
    InMux I__9222 (
            .O(N__38503),
            .I(N__38500));
    LocalMux I__9221 (
            .O(N__38500),
            .I(N__38497));
    Odrv4 I__9220 (
            .O(N__38497),
            .I(M_this_map_address_qc_4_0));
    InMux I__9219 (
            .O(N__38494),
            .I(N__38491));
    LocalMux I__9218 (
            .O(N__38491),
            .I(N__38488));
    Span4Mux_h I__9217 (
            .O(N__38488),
            .I(N__38485));
    Odrv4 I__9216 (
            .O(N__38485),
            .I(N_918_0));
    InMux I__9215 (
            .O(N__38482),
            .I(N__38479));
    LocalMux I__9214 (
            .O(N__38479),
            .I(N__38475));
    InMux I__9213 (
            .O(N__38478),
            .I(N__38472));
    Span12Mux_v I__9212 (
            .O(N__38475),
            .I(N__38469));
    LocalMux I__9211 (
            .O(N__38472),
            .I(N__38466));
    Odrv12 I__9210 (
            .O(N__38469),
            .I(m5_i_a2_i_o3_i_a3));
    Odrv12 I__9209 (
            .O(N__38466),
            .I(m5_i_a2_i_o3_i_a3));
    IoInMux I__9208 (
            .O(N__38461),
            .I(N__38458));
    LocalMux I__9207 (
            .O(N__38458),
            .I(N__38454));
    IoInMux I__9206 (
            .O(N__38457),
            .I(N__38451));
    IoSpan4Mux I__9205 (
            .O(N__38454),
            .I(N__38446));
    LocalMux I__9204 (
            .O(N__38451),
            .I(N__38446));
    IoSpan4Mux I__9203 (
            .O(N__38446),
            .I(N__38442));
    IoInMux I__9202 (
            .O(N__38445),
            .I(N__38439));
    IoSpan4Mux I__9201 (
            .O(N__38442),
            .I(N__38432));
    LocalMux I__9200 (
            .O(N__38439),
            .I(N__38432));
    IoInMux I__9199 (
            .O(N__38438),
            .I(N__38428));
    IoInMux I__9198 (
            .O(N__38437),
            .I(N__38425));
    IoSpan4Mux I__9197 (
            .O(N__38432),
            .I(N__38422));
    IoInMux I__9196 (
            .O(N__38431),
            .I(N__38419));
    LocalMux I__9195 (
            .O(N__38428),
            .I(N__38414));
    LocalMux I__9194 (
            .O(N__38425),
            .I(N__38414));
    IoSpan4Mux I__9193 (
            .O(N__38422),
            .I(N__38408));
    LocalMux I__9192 (
            .O(N__38419),
            .I(N__38408));
    IoSpan4Mux I__9191 (
            .O(N__38414),
            .I(N__38405));
    IoInMux I__9190 (
            .O(N__38413),
            .I(N__38402));
    IoSpan4Mux I__9189 (
            .O(N__38408),
            .I(N__38398));
    IoSpan4Mux I__9188 (
            .O(N__38405),
            .I(N__38395));
    LocalMux I__9187 (
            .O(N__38402),
            .I(N__38392));
    IoInMux I__9186 (
            .O(N__38401),
            .I(N__38389));
    Span4Mux_s1_h I__9185 (
            .O(N__38398),
            .I(N__38386));
    IoSpan4Mux I__9184 (
            .O(N__38395),
            .I(N__38383));
    IoSpan4Mux I__9183 (
            .O(N__38392),
            .I(N__38380));
    LocalMux I__9182 (
            .O(N__38389),
            .I(N__38377));
    Span4Mux_h I__9181 (
            .O(N__38386),
            .I(N__38368));
    Span4Mux_s2_v I__9180 (
            .O(N__38383),
            .I(N__38368));
    Span4Mux_s2_v I__9179 (
            .O(N__38380),
            .I(N__38368));
    Span4Mux_s2_v I__9178 (
            .O(N__38377),
            .I(N__38368));
    Odrv4 I__9177 (
            .O(N__38368),
            .I(N_1048_i_0));
    CEMux I__9176 (
            .O(N__38365),
            .I(N__38361));
    CEMux I__9175 (
            .O(N__38364),
            .I(N__38358));
    LocalMux I__9174 (
            .O(N__38361),
            .I(N__38353));
    LocalMux I__9173 (
            .O(N__38358),
            .I(N__38353));
    Span4Mux_v I__9172 (
            .O(N__38353),
            .I(N__38350));
    Odrv4 I__9171 (
            .O(N__38350),
            .I(\this_spr_ram.mem_WE_12 ));
    CEMux I__9170 (
            .O(N__38347),
            .I(N__38343));
    CEMux I__9169 (
            .O(N__38346),
            .I(N__38340));
    LocalMux I__9168 (
            .O(N__38343),
            .I(N__38337));
    LocalMux I__9167 (
            .O(N__38340),
            .I(N__38334));
    Span4Mux_v I__9166 (
            .O(N__38337),
            .I(N__38331));
    Span4Mux_h I__9165 (
            .O(N__38334),
            .I(N__38328));
    Odrv4 I__9164 (
            .O(N__38331),
            .I(\this_spr_ram.mem_WE_8 ));
    Odrv4 I__9163 (
            .O(N__38328),
            .I(\this_spr_ram.mem_WE_8 ));
    CEMux I__9162 (
            .O(N__38323),
            .I(N__38319));
    CEMux I__9161 (
            .O(N__38322),
            .I(N__38316));
    LocalMux I__9160 (
            .O(N__38319),
            .I(N__38313));
    LocalMux I__9159 (
            .O(N__38316),
            .I(N__38310));
    Span4Mux_h I__9158 (
            .O(N__38313),
            .I(N__38307));
    Span4Mux_h I__9157 (
            .O(N__38310),
            .I(N__38304));
    Span4Mux_v I__9156 (
            .O(N__38307),
            .I(N__38301));
    Span4Mux_v I__9155 (
            .O(N__38304),
            .I(N__38298));
    Span4Mux_v I__9154 (
            .O(N__38301),
            .I(N__38295));
    Span4Mux_v I__9153 (
            .O(N__38298),
            .I(N__38292));
    Odrv4 I__9152 (
            .O(N__38295),
            .I(\this_spr_ram.mem_WE_14 ));
    Odrv4 I__9151 (
            .O(N__38292),
            .I(\this_spr_ram.mem_WE_14 ));
    InMux I__9150 (
            .O(N__38287),
            .I(N__38282));
    InMux I__9149 (
            .O(N__38286),
            .I(N__38277));
    InMux I__9148 (
            .O(N__38285),
            .I(N__38277));
    LocalMux I__9147 (
            .O(N__38282),
            .I(N__38270));
    LocalMux I__9146 (
            .O(N__38277),
            .I(N__38270));
    InMux I__9145 (
            .O(N__38276),
            .I(N__38265));
    InMux I__9144 (
            .O(N__38275),
            .I(N__38265));
    Odrv4 I__9143 (
            .O(N__38270),
            .I(M_this_state_qZ0Z_6));
    LocalMux I__9142 (
            .O(N__38265),
            .I(M_this_state_qZ0Z_6));
    InMux I__9141 (
            .O(N__38260),
            .I(N__38257));
    LocalMux I__9140 (
            .O(N__38257),
            .I(this_ppu_un1_M_this_state_q_7_i_0_0_0));
    CascadeMux I__9139 (
            .O(N__38254),
            .I(un1_M_this_state_q_7_i_0_a3_0_0_cascade_));
    InMux I__9138 (
            .O(N__38251),
            .I(N__38248));
    LocalMux I__9137 (
            .O(N__38248),
            .I(N__38245));
    Span4Mux_h I__9136 (
            .O(N__38245),
            .I(N__38242));
    Span4Mux_h I__9135 (
            .O(N__38242),
            .I(N__38239));
    Span4Mux_h I__9134 (
            .O(N__38239),
            .I(N__38236));
    Odrv4 I__9133 (
            .O(N__38236),
            .I(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0 ));
    InMux I__9132 (
            .O(N__38233),
            .I(N__38230));
    LocalMux I__9131 (
            .O(N__38230),
            .I(N__38227));
    Span4Mux_v I__9130 (
            .O(N__38227),
            .I(N__38223));
    InMux I__9129 (
            .O(N__38226),
            .I(N__38220));
    Sp12to4 I__9128 (
            .O(N__38223),
            .I(N__38217));
    LocalMux I__9127 (
            .O(N__38220),
            .I(N__38214));
    Span12Mux_h I__9126 (
            .O(N__38217),
            .I(N__38209));
    Span12Mux_v I__9125 (
            .O(N__38214),
            .I(N__38209));
    Odrv12 I__9124 (
            .O(N__38209),
            .I(M_this_map_ram_read_data_0));
    InMux I__9123 (
            .O(N__38206),
            .I(N__38199));
    InMux I__9122 (
            .O(N__38205),
            .I(N__38199));
    InMux I__9121 (
            .O(N__38204),
            .I(N__38195));
    LocalMux I__9120 (
            .O(N__38199),
            .I(N__38192));
    InMux I__9119 (
            .O(N__38198),
            .I(N__38189));
    LocalMux I__9118 (
            .O(N__38195),
            .I(N__38184));
    Span4Mux_v I__9117 (
            .O(N__38192),
            .I(N__38179));
    LocalMux I__9116 (
            .O(N__38189),
            .I(N__38179));
    InMux I__9115 (
            .O(N__38188),
            .I(N__38169));
    InMux I__9114 (
            .O(N__38187),
            .I(N__38169));
    Span4Mux_v I__9113 (
            .O(N__38184),
            .I(N__38164));
    Span4Mux_v I__9112 (
            .O(N__38179),
            .I(N__38164));
    InMux I__9111 (
            .O(N__38178),
            .I(N__38152));
    InMux I__9110 (
            .O(N__38177),
            .I(N__38152));
    InMux I__9109 (
            .O(N__38176),
            .I(N__38152));
    InMux I__9108 (
            .O(N__38175),
            .I(N__38152));
    InMux I__9107 (
            .O(N__38174),
            .I(N__38152));
    LocalMux I__9106 (
            .O(N__38169),
            .I(N__38147));
    Span4Mux_h I__9105 (
            .O(N__38164),
            .I(N__38144));
    InMux I__9104 (
            .O(N__38163),
            .I(N__38141));
    LocalMux I__9103 (
            .O(N__38152),
            .I(N__38138));
    InMux I__9102 (
            .O(N__38151),
            .I(N__38135));
    InMux I__9101 (
            .O(N__38150),
            .I(N__38132));
    Span4Mux_h I__9100 (
            .O(N__38147),
            .I(N__38129));
    Span4Mux_h I__9099 (
            .O(N__38144),
            .I(N__38126));
    LocalMux I__9098 (
            .O(N__38141),
            .I(N__38121));
    Span4Mux_v I__9097 (
            .O(N__38138),
            .I(N__38121));
    LocalMux I__9096 (
            .O(N__38135),
            .I(N__38114));
    LocalMux I__9095 (
            .O(N__38132),
            .I(N__38114));
    Span4Mux_h I__9094 (
            .O(N__38129),
            .I(N__38114));
    Odrv4 I__9093 (
            .O(N__38126),
            .I(\this_ppu.N_785_0 ));
    Odrv4 I__9092 (
            .O(N__38121),
            .I(\this_ppu.N_785_0 ));
    Odrv4 I__9091 (
            .O(N__38114),
            .I(\this_ppu.N_785_0 ));
    CascadeMux I__9090 (
            .O(N__38107),
            .I(N__38101));
    CascadeMux I__9089 (
            .O(N__38106),
            .I(N__38098));
    CascadeMux I__9088 (
            .O(N__38105),
            .I(N__38094));
    CascadeMux I__9087 (
            .O(N__38104),
            .I(N__38091));
    InMux I__9086 (
            .O(N__38101),
            .I(N__38087));
    InMux I__9085 (
            .O(N__38098),
            .I(N__38084));
    CascadeMux I__9084 (
            .O(N__38097),
            .I(N__38081));
    InMux I__9083 (
            .O(N__38094),
            .I(N__38076));
    InMux I__9082 (
            .O(N__38091),
            .I(N__38073));
    CascadeMux I__9081 (
            .O(N__38090),
            .I(N__38070));
    LocalMux I__9080 (
            .O(N__38087),
            .I(N__38063));
    LocalMux I__9079 (
            .O(N__38084),
            .I(N__38063));
    InMux I__9078 (
            .O(N__38081),
            .I(N__38060));
    CascadeMux I__9077 (
            .O(N__38080),
            .I(N__38057));
    CascadeMux I__9076 (
            .O(N__38079),
            .I(N__38054));
    LocalMux I__9075 (
            .O(N__38076),
            .I(N__38050));
    LocalMux I__9074 (
            .O(N__38073),
            .I(N__38047));
    InMux I__9073 (
            .O(N__38070),
            .I(N__38044));
    CascadeMux I__9072 (
            .O(N__38069),
            .I(N__38041));
    CascadeMux I__9071 (
            .O(N__38068),
            .I(N__38034));
    Span4Mux_v I__9070 (
            .O(N__38063),
            .I(N__38029));
    LocalMux I__9069 (
            .O(N__38060),
            .I(N__38029));
    InMux I__9068 (
            .O(N__38057),
            .I(N__38026));
    InMux I__9067 (
            .O(N__38054),
            .I(N__38023));
    CascadeMux I__9066 (
            .O(N__38053),
            .I(N__38020));
    Span4Mux_v I__9065 (
            .O(N__38050),
            .I(N__38013));
    Span4Mux_h I__9064 (
            .O(N__38047),
            .I(N__38013));
    LocalMux I__9063 (
            .O(N__38044),
            .I(N__38013));
    InMux I__9062 (
            .O(N__38041),
            .I(N__38010));
    CascadeMux I__9061 (
            .O(N__38040),
            .I(N__38007));
    CascadeMux I__9060 (
            .O(N__38039),
            .I(N__38004));
    CascadeMux I__9059 (
            .O(N__38038),
            .I(N__38001));
    CascadeMux I__9058 (
            .O(N__38037),
            .I(N__37998));
    InMux I__9057 (
            .O(N__38034),
            .I(N__37994));
    Span4Mux_h I__9056 (
            .O(N__38029),
            .I(N__37991));
    LocalMux I__9055 (
            .O(N__38026),
            .I(N__37986));
    LocalMux I__9054 (
            .O(N__38023),
            .I(N__37986));
    InMux I__9053 (
            .O(N__38020),
            .I(N__37983));
    Span4Mux_v I__9052 (
            .O(N__38013),
            .I(N__37978));
    LocalMux I__9051 (
            .O(N__38010),
            .I(N__37978));
    InMux I__9050 (
            .O(N__38007),
            .I(N__37975));
    InMux I__9049 (
            .O(N__38004),
            .I(N__37972));
    InMux I__9048 (
            .O(N__38001),
            .I(N__37969));
    InMux I__9047 (
            .O(N__37998),
            .I(N__37966));
    CascadeMux I__9046 (
            .O(N__37997),
            .I(N__37963));
    LocalMux I__9045 (
            .O(N__37994),
            .I(N__37960));
    Span4Mux_v I__9044 (
            .O(N__37991),
            .I(N__37957));
    Span12Mux_s10_v I__9043 (
            .O(N__37986),
            .I(N__37946));
    LocalMux I__9042 (
            .O(N__37983),
            .I(N__37946));
    Sp12to4 I__9041 (
            .O(N__37978),
            .I(N__37946));
    LocalMux I__9040 (
            .O(N__37975),
            .I(N__37946));
    LocalMux I__9039 (
            .O(N__37972),
            .I(N__37946));
    LocalMux I__9038 (
            .O(N__37969),
            .I(N__37943));
    LocalMux I__9037 (
            .O(N__37966),
            .I(N__37940));
    InMux I__9036 (
            .O(N__37963),
            .I(N__37937));
    Span4Mux_v I__9035 (
            .O(N__37960),
            .I(N__37934));
    Sp12to4 I__9034 (
            .O(N__37957),
            .I(N__37929));
    Span12Mux_v I__9033 (
            .O(N__37946),
            .I(N__37929));
    Span4Mux_h I__9032 (
            .O(N__37943),
            .I(N__37924));
    Span4Mux_h I__9031 (
            .O(N__37940),
            .I(N__37924));
    LocalMux I__9030 (
            .O(N__37937),
            .I(N__37921));
    Odrv4 I__9029 (
            .O(N__37934),
            .I(read_data_RNI4PFJ1_0));
    Odrv12 I__9028 (
            .O(N__37929),
            .I(read_data_RNI4PFJ1_0));
    Odrv4 I__9027 (
            .O(N__37924),
            .I(read_data_RNI4PFJ1_0));
    Odrv12 I__9026 (
            .O(N__37921),
            .I(read_data_RNI4PFJ1_0));
    CascadeMux I__9025 (
            .O(N__37912),
            .I(N__37909));
    InMux I__9024 (
            .O(N__37909),
            .I(N__37906));
    LocalMux I__9023 (
            .O(N__37906),
            .I(N__37903));
    Odrv4 I__9022 (
            .O(N__37903),
            .I(N_1058));
    CascadeMux I__9021 (
            .O(N__37900),
            .I(N_1062_cascade_));
    InMux I__9020 (
            .O(N__37897),
            .I(N__37894));
    LocalMux I__9019 (
            .O(N__37894),
            .I(M_this_map_address_qc_5_0));
    InMux I__9018 (
            .O(N__37891),
            .I(N__37888));
    LocalMux I__9017 (
            .O(N__37888),
            .I(N__37885));
    Sp12to4 I__9016 (
            .O(N__37885),
            .I(N__37882));
    Span12Mux_v I__9015 (
            .O(N__37882),
            .I(N__37879));
    Span12Mux_h I__9014 (
            .O(N__37879),
            .I(N__37876));
    Odrv12 I__9013 (
            .O(N__37876),
            .I(\this_spr_ram.mem_out_bus7_2 ));
    InMux I__9012 (
            .O(N__37873),
            .I(N__37870));
    LocalMux I__9011 (
            .O(N__37870),
            .I(N__37867));
    Span4Mux_v I__9010 (
            .O(N__37867),
            .I(N__37864));
    Odrv4 I__9009 (
            .O(N__37864),
            .I(\this_spr_ram.mem_out_bus3_2 ));
    InMux I__9008 (
            .O(N__37861),
            .I(N__37858));
    LocalMux I__9007 (
            .O(N__37858),
            .I(N__37855));
    Span4Mux_h I__9006 (
            .O(N__37855),
            .I(N__37852));
    Odrv4 I__9005 (
            .O(N__37852),
            .I(\this_spr_ram.mem_mem_3_1_RNISI5GZ0 ));
    CascadeMux I__9004 (
            .O(N__37849),
            .I(N__37846));
    InMux I__9003 (
            .O(N__37846),
            .I(N__37843));
    LocalMux I__9002 (
            .O(N__37843),
            .I(N__37840));
    Span12Mux_h I__9001 (
            .O(N__37840),
            .I(N__37837));
    Span12Mux_v I__9000 (
            .O(N__37837),
            .I(N__37834));
    Odrv12 I__8999 (
            .O(N__37834),
            .I(\this_spr_ram.mem_out_bus7_3 ));
    InMux I__8998 (
            .O(N__37831),
            .I(N__37828));
    LocalMux I__8997 (
            .O(N__37828),
            .I(N__37825));
    Span4Mux_h I__8996 (
            .O(N__37825),
            .I(N__37822));
    Odrv4 I__8995 (
            .O(N__37822),
            .I(\this_spr_ram.mem_out_bus3_3 ));
    InMux I__8994 (
            .O(N__37819),
            .I(N__37816));
    LocalMux I__8993 (
            .O(N__37816),
            .I(\this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0 ));
    InMux I__8992 (
            .O(N__37813),
            .I(N__37810));
    LocalMux I__8991 (
            .O(N__37810),
            .I(N__37807));
    Span4Mux_v I__8990 (
            .O(N__37807),
            .I(N__37804));
    Sp12to4 I__8989 (
            .O(N__37804),
            .I(N__37801));
    Span12Mux_h I__8988 (
            .O(N__37801),
            .I(N__37797));
    InMux I__8987 (
            .O(N__37800),
            .I(N__37794));
    Odrv12 I__8986 (
            .O(N__37797),
            .I(M_this_ctrl_flags_qZ0Z_7));
    LocalMux I__8985 (
            .O(N__37794),
            .I(M_this_ctrl_flags_qZ0Z_7));
    InMux I__8984 (
            .O(N__37789),
            .I(N__37786));
    LocalMux I__8983 (
            .O(N__37786),
            .I(N__37782));
    InMux I__8982 (
            .O(N__37785),
            .I(N__37778));
    Span4Mux_v I__8981 (
            .O(N__37782),
            .I(N__37775));
    InMux I__8980 (
            .O(N__37781),
            .I(N__37772));
    LocalMux I__8979 (
            .O(N__37778),
            .I(N__37769));
    Odrv4 I__8978 (
            .O(N__37775),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__8977 (
            .O(N__37772),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__8976 (
            .O(N__37769),
            .I(M_this_state_qZ0Z_2));
    IoInMux I__8975 (
            .O(N__37762),
            .I(N__37759));
    LocalMux I__8974 (
            .O(N__37759),
            .I(N__37756));
    Span4Mux_s2_h I__8973 (
            .O(N__37756),
            .I(N__37752));
    InMux I__8972 (
            .O(N__37755),
            .I(N__37749));
    Sp12to4 I__8971 (
            .O(N__37752),
            .I(N__37744));
    LocalMux I__8970 (
            .O(N__37749),
            .I(N__37741));
    InMux I__8969 (
            .O(N__37748),
            .I(N__37737));
    InMux I__8968 (
            .O(N__37747),
            .I(N__37731));
    Span12Mux_s10_v I__8967 (
            .O(N__37744),
            .I(N__37727));
    Span4Mux_v I__8966 (
            .O(N__37741),
            .I(N__37724));
    InMux I__8965 (
            .O(N__37740),
            .I(N__37721));
    LocalMux I__8964 (
            .O(N__37737),
            .I(N__37718));
    InMux I__8963 (
            .O(N__37736),
            .I(N__37715));
    InMux I__8962 (
            .O(N__37735),
            .I(N__37712));
    InMux I__8961 (
            .O(N__37734),
            .I(N__37709));
    LocalMux I__8960 (
            .O(N__37731),
            .I(N__37706));
    InMux I__8959 (
            .O(N__37730),
            .I(N__37703));
    Span12Mux_h I__8958 (
            .O(N__37727),
            .I(N__37700));
    Sp12to4 I__8957 (
            .O(N__37724),
            .I(N__37697));
    LocalMux I__8956 (
            .O(N__37721),
            .I(N__37693));
    Span4Mux_v I__8955 (
            .O(N__37718),
            .I(N__37688));
    LocalMux I__8954 (
            .O(N__37715),
            .I(N__37688));
    LocalMux I__8953 (
            .O(N__37712),
            .I(N__37685));
    LocalMux I__8952 (
            .O(N__37709),
            .I(N__37682));
    Span4Mux_v I__8951 (
            .O(N__37706),
            .I(N__37677));
    LocalMux I__8950 (
            .O(N__37703),
            .I(N__37677));
    Span12Mux_v I__8949 (
            .O(N__37700),
            .I(N__37674));
    Span12Mux_s6_h I__8948 (
            .O(N__37697),
            .I(N__37671));
    InMux I__8947 (
            .O(N__37696),
            .I(N__37668));
    Span4Mux_v I__8946 (
            .O(N__37693),
            .I(N__37665));
    Span4Mux_h I__8945 (
            .O(N__37688),
            .I(N__37662));
    Span12Mux_h I__8944 (
            .O(N__37685),
            .I(N__37657));
    Span12Mux_h I__8943 (
            .O(N__37682),
            .I(N__37657));
    Span4Mux_h I__8942 (
            .O(N__37677),
            .I(N__37654));
    Odrv12 I__8941 (
            .O(N__37674),
            .I(N_38_i_0));
    Odrv12 I__8940 (
            .O(N__37671),
            .I(N_38_i_0));
    LocalMux I__8939 (
            .O(N__37668),
            .I(N_38_i_0));
    Odrv4 I__8938 (
            .O(N__37665),
            .I(N_38_i_0));
    Odrv4 I__8937 (
            .O(N__37662),
            .I(N_38_i_0));
    Odrv12 I__8936 (
            .O(N__37657),
            .I(N_38_i_0));
    Odrv4 I__8935 (
            .O(N__37654),
            .I(N_38_i_0));
    IoInMux I__8934 (
            .O(N__37639),
            .I(N__37636));
    LocalMux I__8933 (
            .O(N__37636),
            .I(N__37632));
    IoInMux I__8932 (
            .O(N__37635),
            .I(N__37629));
    IoSpan4Mux I__8931 (
            .O(N__37632),
            .I(N__37624));
    LocalMux I__8930 (
            .O(N__37629),
            .I(N__37624));
    IoSpan4Mux I__8929 (
            .O(N__37624),
            .I(N__37619));
    IoInMux I__8928 (
            .O(N__37623),
            .I(N__37616));
    IoInMux I__8927 (
            .O(N__37622),
            .I(N__37613));
    IoSpan4Mux I__8926 (
            .O(N__37619),
            .I(N__37601));
    LocalMux I__8925 (
            .O(N__37616),
            .I(N__37601));
    LocalMux I__8924 (
            .O(N__37613),
            .I(N__37598));
    IoInMux I__8923 (
            .O(N__37612),
            .I(N__37595));
    IoInMux I__8922 (
            .O(N__37611),
            .I(N__37592));
    IoInMux I__8921 (
            .O(N__37610),
            .I(N__37589));
    IoInMux I__8920 (
            .O(N__37609),
            .I(N__37586));
    IoInMux I__8919 (
            .O(N__37608),
            .I(N__37581));
    IoInMux I__8918 (
            .O(N__37607),
            .I(N__37578));
    IoInMux I__8917 (
            .O(N__37606),
            .I(N__37573));
    IoSpan4Mux I__8916 (
            .O(N__37601),
            .I(N__37570));
    IoSpan4Mux I__8915 (
            .O(N__37598),
            .I(N__37563));
    LocalMux I__8914 (
            .O(N__37595),
            .I(N__37563));
    LocalMux I__8913 (
            .O(N__37592),
            .I(N__37563));
    LocalMux I__8912 (
            .O(N__37589),
            .I(N__37558));
    LocalMux I__8911 (
            .O(N__37586),
            .I(N__37555));
    IoInMux I__8910 (
            .O(N__37585),
            .I(N__37552));
    IoInMux I__8909 (
            .O(N__37584),
            .I(N__37549));
    LocalMux I__8908 (
            .O(N__37581),
            .I(N__37544));
    LocalMux I__8907 (
            .O(N__37578),
            .I(N__37544));
    IoInMux I__8906 (
            .O(N__37577),
            .I(N__37541));
    IoInMux I__8905 (
            .O(N__37576),
            .I(N__37538));
    LocalMux I__8904 (
            .O(N__37573),
            .I(N__37535));
    IoSpan4Mux I__8903 (
            .O(N__37570),
            .I(N__37530));
    IoSpan4Mux I__8902 (
            .O(N__37563),
            .I(N__37530));
    IoInMux I__8901 (
            .O(N__37562),
            .I(N__37527));
    IoInMux I__8900 (
            .O(N__37561),
            .I(N__37524));
    IoSpan4Mux I__8899 (
            .O(N__37558),
            .I(N__37521));
    IoSpan4Mux I__8898 (
            .O(N__37555),
            .I(N__37514));
    LocalMux I__8897 (
            .O(N__37552),
            .I(N__37514));
    LocalMux I__8896 (
            .O(N__37549),
            .I(N__37514));
    IoSpan4Mux I__8895 (
            .O(N__37544),
            .I(N__37507));
    LocalMux I__8894 (
            .O(N__37541),
            .I(N__37507));
    LocalMux I__8893 (
            .O(N__37538),
            .I(N__37507));
    Span4Mux_s1_h I__8892 (
            .O(N__37535),
            .I(N__37504));
    Span4Mux_s1_h I__8891 (
            .O(N__37530),
            .I(N__37501));
    LocalMux I__8890 (
            .O(N__37527),
            .I(N__37496));
    LocalMux I__8889 (
            .O(N__37524),
            .I(N__37496));
    Span4Mux_s3_h I__8888 (
            .O(N__37521),
            .I(N__37493));
    IoSpan4Mux I__8887 (
            .O(N__37514),
            .I(N__37488));
    IoSpan4Mux I__8886 (
            .O(N__37507),
            .I(N__37488));
    Span4Mux_v I__8885 (
            .O(N__37504),
            .I(N__37481));
    Span4Mux_v I__8884 (
            .O(N__37501),
            .I(N__37481));
    Span4Mux_s1_h I__8883 (
            .O(N__37496),
            .I(N__37481));
    Sp12to4 I__8882 (
            .O(N__37493),
            .I(N__37478));
    Span4Mux_s3_v I__8881 (
            .O(N__37488),
            .I(N__37475));
    Span4Mux_h I__8880 (
            .O(N__37481),
            .I(N__37472));
    Span12Mux_s11_h I__8879 (
            .O(N__37478),
            .I(N__37469));
    Span4Mux_v I__8878 (
            .O(N__37475),
            .I(N__37464));
    Span4Mux_h I__8877 (
            .O(N__37472),
            .I(N__37464));
    Odrv12 I__8876 (
            .O(N__37469),
            .I(N_38_i_0_i));
    Odrv4 I__8875 (
            .O(N__37464),
            .I(N_38_i_0_i));
    InMux I__8874 (
            .O(N__37459),
            .I(N__37456));
    LocalMux I__8873 (
            .O(N__37456),
            .I(N__37452));
    InMux I__8872 (
            .O(N__37455),
            .I(N__37449));
    Span4Mux_h I__8871 (
            .O(N__37452),
            .I(N__37446));
    LocalMux I__8870 (
            .O(N__37449),
            .I(\this_ppu.N_856_0 ));
    Odrv4 I__8869 (
            .O(N__37446),
            .I(\this_ppu.N_856_0 ));
    CascadeMux I__8868 (
            .O(N__37441),
            .I(this_ppu_un1_M_this_state_q_7_i_0_0_0_cascade_));
    InMux I__8867 (
            .O(N__37438),
            .I(N__37434));
    InMux I__8866 (
            .O(N__37437),
            .I(N__37431));
    LocalMux I__8865 (
            .O(N__37434),
            .I(N__37428));
    LocalMux I__8864 (
            .O(N__37431),
            .I(N__37423));
    Span4Mux_h I__8863 (
            .O(N__37428),
            .I(N__37420));
    InMux I__8862 (
            .O(N__37427),
            .I(N__37417));
    InMux I__8861 (
            .O(N__37426),
            .I(N__37414));
    Odrv12 I__8860 (
            .O(N__37423),
            .I(N_816_0));
    Odrv4 I__8859 (
            .O(N__37420),
            .I(N_816_0));
    LocalMux I__8858 (
            .O(N__37417),
            .I(N_816_0));
    LocalMux I__8857 (
            .O(N__37414),
            .I(N_816_0));
    InMux I__8856 (
            .O(N__37405),
            .I(N__37402));
    LocalMux I__8855 (
            .O(N__37402),
            .I(N_1416));
    InMux I__8854 (
            .O(N__37399),
            .I(N__37396));
    LocalMux I__8853 (
            .O(N__37396),
            .I(N__37391));
    InMux I__8852 (
            .O(N__37395),
            .I(N__37388));
    InMux I__8851 (
            .O(N__37394),
            .I(N__37383));
    Span4Mux_v I__8850 (
            .O(N__37391),
            .I(N__37378));
    LocalMux I__8849 (
            .O(N__37388),
            .I(N__37378));
    InMux I__8848 (
            .O(N__37387),
            .I(N__37375));
    InMux I__8847 (
            .O(N__37386),
            .I(N__37372));
    LocalMux I__8846 (
            .O(N__37383),
            .I(N__37369));
    Odrv4 I__8845 (
            .O(N__37378),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__8844 (
            .O(N__37375),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__8843 (
            .O(N__37372),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__8842 (
            .O(N__37369),
            .I(M_this_state_qZ0Z_5));
    IoInMux I__8841 (
            .O(N__37360),
            .I(N__37357));
    LocalMux I__8840 (
            .O(N__37357),
            .I(N__37354));
    Span12Mux_s9_h I__8839 (
            .O(N__37354),
            .I(N__37351));
    Span12Mux_v I__8838 (
            .O(N__37351),
            .I(N__37348));
    Odrv12 I__8837 (
            .O(N__37348),
            .I(led_c_6));
    CascadeMux I__8836 (
            .O(N__37345),
            .I(N__37340));
    InMux I__8835 (
            .O(N__37344),
            .I(N__37337));
    InMux I__8834 (
            .O(N__37343),
            .I(N__37334));
    InMux I__8833 (
            .O(N__37340),
            .I(N__37331));
    LocalMux I__8832 (
            .O(N__37337),
            .I(N__37322));
    LocalMux I__8831 (
            .O(N__37334),
            .I(N__37322));
    LocalMux I__8830 (
            .O(N__37331),
            .I(N__37322));
    InMux I__8829 (
            .O(N__37330),
            .I(N__37319));
    InMux I__8828 (
            .O(N__37329),
            .I(N__37315));
    Span4Mux_h I__8827 (
            .O(N__37322),
            .I(N__37312));
    LocalMux I__8826 (
            .O(N__37319),
            .I(N__37309));
    InMux I__8825 (
            .O(N__37318),
            .I(N__37306));
    LocalMux I__8824 (
            .O(N__37315),
            .I(N__37303));
    Span4Mux_h I__8823 (
            .O(N__37312),
            .I(N__37298));
    Span4Mux_v I__8822 (
            .O(N__37309),
            .I(N__37298));
    LocalMux I__8821 (
            .O(N__37306),
            .I(\this_ppu.M_screen_y_qZ0Z_4 ));
    Odrv4 I__8820 (
            .O(N__37303),
            .I(\this_ppu.M_screen_y_qZ0Z_4 ));
    Odrv4 I__8819 (
            .O(N__37298),
            .I(\this_ppu.M_screen_y_qZ0Z_4 ));
    InMux I__8818 (
            .O(N__37291),
            .I(N__37286));
    InMux I__8817 (
            .O(N__37290),
            .I(N__37283));
    InMux I__8816 (
            .O(N__37289),
            .I(N__37280));
    LocalMux I__8815 (
            .O(N__37286),
            .I(N__37275));
    LocalMux I__8814 (
            .O(N__37283),
            .I(N__37275));
    LocalMux I__8813 (
            .O(N__37280),
            .I(N__37272));
    Span12Mux_h I__8812 (
            .O(N__37275),
            .I(N__37269));
    Odrv4 I__8811 (
            .O(N__37272),
            .I(\this_ppu.un3_M_screen_y_d_0_c4 ));
    Odrv12 I__8810 (
            .O(N__37269),
            .I(\this_ppu.un3_M_screen_y_d_0_c4 ));
    InMux I__8809 (
            .O(N__37264),
            .I(N__37261));
    LocalMux I__8808 (
            .O(N__37261),
            .I(N__37256));
    InMux I__8807 (
            .O(N__37260),
            .I(N__37245));
    InMux I__8806 (
            .O(N__37259),
            .I(N__37245));
    Span4Mux_h I__8805 (
            .O(N__37256),
            .I(N__37242));
    CascadeMux I__8804 (
            .O(N__37255),
            .I(N__37239));
    InMux I__8803 (
            .O(N__37254),
            .I(N__37222));
    InMux I__8802 (
            .O(N__37253),
            .I(N__37222));
    InMux I__8801 (
            .O(N__37252),
            .I(N__37222));
    InMux I__8800 (
            .O(N__37251),
            .I(N__37222));
    InMux I__8799 (
            .O(N__37250),
            .I(N__37222));
    LocalMux I__8798 (
            .O(N__37245),
            .I(N__37219));
    Span4Mux_h I__8797 (
            .O(N__37242),
            .I(N__37216));
    InMux I__8796 (
            .O(N__37239),
            .I(N__37213));
    InMux I__8795 (
            .O(N__37238),
            .I(N__37210));
    InMux I__8794 (
            .O(N__37237),
            .I(N__37207));
    InMux I__8793 (
            .O(N__37236),
            .I(N__37200));
    InMux I__8792 (
            .O(N__37235),
            .I(N__37200));
    InMux I__8791 (
            .O(N__37234),
            .I(N__37200));
    InMux I__8790 (
            .O(N__37233),
            .I(N__37197));
    LocalMux I__8789 (
            .O(N__37222),
            .I(N__37194));
    Odrv4 I__8788 (
            .O(N__37219),
            .I(N_861_0));
    Odrv4 I__8787 (
            .O(N__37216),
            .I(N_861_0));
    LocalMux I__8786 (
            .O(N__37213),
            .I(N_861_0));
    LocalMux I__8785 (
            .O(N__37210),
            .I(N_861_0));
    LocalMux I__8784 (
            .O(N__37207),
            .I(N_861_0));
    LocalMux I__8783 (
            .O(N__37200),
            .I(N_861_0));
    LocalMux I__8782 (
            .O(N__37197),
            .I(N_861_0));
    Odrv4 I__8781 (
            .O(N__37194),
            .I(N_861_0));
    CEMux I__8780 (
            .O(N__37177),
            .I(N__37173));
    CEMux I__8779 (
            .O(N__37176),
            .I(N__37170));
    LocalMux I__8778 (
            .O(N__37173),
            .I(N__37166));
    LocalMux I__8777 (
            .O(N__37170),
            .I(N__37162));
    CEMux I__8776 (
            .O(N__37169),
            .I(N__37159));
    Span4Mux_v I__8775 (
            .O(N__37166),
            .I(N__37156));
    CEMux I__8774 (
            .O(N__37165),
            .I(N__37153));
    Span4Mux_h I__8773 (
            .O(N__37162),
            .I(N__37150));
    LocalMux I__8772 (
            .O(N__37159),
            .I(N__37147));
    Sp12to4 I__8771 (
            .O(N__37156),
            .I(N__37142));
    LocalMux I__8770 (
            .O(N__37153),
            .I(N__37142));
    Odrv4 I__8769 (
            .O(N__37150),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_0 ));
    Odrv4 I__8768 (
            .O(N__37147),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_0 ));
    Odrv12 I__8767 (
            .O(N__37142),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_0 ));
    InMux I__8766 (
            .O(N__37135),
            .I(N__37130));
    CascadeMux I__8765 (
            .O(N__37134),
            .I(N__37127));
    CascadeMux I__8764 (
            .O(N__37133),
            .I(N__37124));
    LocalMux I__8763 (
            .O(N__37130),
            .I(N__37119));
    InMux I__8762 (
            .O(N__37127),
            .I(N__37116));
    InMux I__8761 (
            .O(N__37124),
            .I(N__37111));
    InMux I__8760 (
            .O(N__37123),
            .I(N__37111));
    InMux I__8759 (
            .O(N__37122),
            .I(N__37108));
    Span12Mux_h I__8758 (
            .O(N__37119),
            .I(N__37105));
    LocalMux I__8757 (
            .O(N__37116),
            .I(N__37100));
    LocalMux I__8756 (
            .O(N__37111),
            .I(N__37100));
    LocalMux I__8755 (
            .O(N__37108),
            .I(\this_ppu.M_screen_y_qZ0Z_5 ));
    Odrv12 I__8754 (
            .O(N__37105),
            .I(\this_ppu.M_screen_y_qZ0Z_5 ));
    Odrv4 I__8753 (
            .O(N__37100),
            .I(\this_ppu.M_screen_y_qZ0Z_5 ));
    CascadeMux I__8752 (
            .O(N__37093),
            .I(N__37090));
    InMux I__8751 (
            .O(N__37090),
            .I(N__37087));
    LocalMux I__8750 (
            .O(N__37087),
            .I(N__37083));
    CascadeMux I__8749 (
            .O(N__37086),
            .I(N__37080));
    Span4Mux_v I__8748 (
            .O(N__37083),
            .I(N__37077));
    InMux I__8747 (
            .O(N__37080),
            .I(N__37074));
    Span4Mux_h I__8746 (
            .O(N__37077),
            .I(N__37071));
    LocalMux I__8745 (
            .O(N__37074),
            .I(N__37068));
    Span4Mux_h I__8744 (
            .O(N__37071),
            .I(N__37063));
    Span4Mux_h I__8743 (
            .O(N__37068),
            .I(N__37063));
    Odrv4 I__8742 (
            .O(N__37063),
            .I(M_this_scroll_qZ0Z_5));
    InMux I__8741 (
            .O(N__37060),
            .I(N__37057));
    LocalMux I__8740 (
            .O(N__37057),
            .I(N__37054));
    Span4Mux_h I__8739 (
            .O(N__37054),
            .I(N__37051));
    Span4Mux_h I__8738 (
            .O(N__37051),
            .I(N__37048));
    Span4Mux_h I__8737 (
            .O(N__37048),
            .I(N__37045));
    Odrv4 I__8736 (
            .O(N__37045),
            .I(\this_ppu.M_screen_y_q_esr_RNIJB7F7Z0Z_5 ));
    CascadeMux I__8735 (
            .O(N__37042),
            .I(N__37039));
    InMux I__8734 (
            .O(N__37039),
            .I(N__37034));
    InMux I__8733 (
            .O(N__37038),
            .I(N__37031));
    InMux I__8732 (
            .O(N__37037),
            .I(N__37028));
    LocalMux I__8731 (
            .O(N__37034),
            .I(N__37020));
    LocalMux I__8730 (
            .O(N__37031),
            .I(N__37020));
    LocalMux I__8729 (
            .O(N__37028),
            .I(N__37020));
    InMux I__8728 (
            .O(N__37027),
            .I(N__37017));
    Span4Mux_v I__8727 (
            .O(N__37020),
            .I(N__37014));
    LocalMux I__8726 (
            .O(N__37017),
            .I(\this_spr_ram.mem_radregZ0Z_12 ));
    Odrv4 I__8725 (
            .O(N__37014),
            .I(\this_spr_ram.mem_radregZ0Z_12 ));
    InMux I__8724 (
            .O(N__37009),
            .I(N__37006));
    LocalMux I__8723 (
            .O(N__37006),
            .I(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0 ));
    CascadeMux I__8722 (
            .O(N__37003),
            .I(N__36996));
    InMux I__8721 (
            .O(N__37002),
            .I(N__36992));
    InMux I__8720 (
            .O(N__37001),
            .I(N__36987));
    InMux I__8719 (
            .O(N__37000),
            .I(N__36987));
    InMux I__8718 (
            .O(N__36999),
            .I(N__36980));
    InMux I__8717 (
            .O(N__36996),
            .I(N__36980));
    InMux I__8716 (
            .O(N__36995),
            .I(N__36980));
    LocalMux I__8715 (
            .O(N__36992),
            .I(N__36975));
    LocalMux I__8714 (
            .O(N__36987),
            .I(N__36972));
    LocalMux I__8713 (
            .O(N__36980),
            .I(N__36969));
    InMux I__8712 (
            .O(N__36979),
            .I(N__36964));
    InMux I__8711 (
            .O(N__36978),
            .I(N__36964));
    Span4Mux_h I__8710 (
            .O(N__36975),
            .I(N__36961));
    Odrv4 I__8709 (
            .O(N__36972),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    Odrv4 I__8708 (
            .O(N__36969),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    LocalMux I__8707 (
            .O(N__36964),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    Odrv4 I__8706 (
            .O(N__36961),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    CascadeMux I__8705 (
            .O(N__36952),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ));
    InMux I__8704 (
            .O(N__36949),
            .I(N__36946));
    LocalMux I__8703 (
            .O(N__36946),
            .I(N__36942));
    InMux I__8702 (
            .O(N__36945),
            .I(N__36939));
    Odrv4 I__8701 (
            .O(N__36942),
            .I(M_this_spr_ram_read_data_3));
    LocalMux I__8700 (
            .O(N__36939),
            .I(M_this_spr_ram_read_data_3));
    InMux I__8699 (
            .O(N__36934),
            .I(N__36931));
    LocalMux I__8698 (
            .O(N__36931),
            .I(N__36928));
    Span4Mux_h I__8697 (
            .O(N__36928),
            .I(N__36925));
    Span4Mux_v I__8696 (
            .O(N__36925),
            .I(N__36922));
    Odrv4 I__8695 (
            .O(N__36922),
            .I(\this_spr_ram.mem_out_bus5_3 ));
    InMux I__8694 (
            .O(N__36919),
            .I(N__36916));
    LocalMux I__8693 (
            .O(N__36916),
            .I(N__36913));
    Span4Mux_h I__8692 (
            .O(N__36913),
            .I(N__36910));
    Span4Mux_v I__8691 (
            .O(N__36910),
            .I(N__36907));
    Span4Mux_v I__8690 (
            .O(N__36907),
            .I(N__36904));
    Odrv4 I__8689 (
            .O(N__36904),
            .I(\this_spr_ram.mem_out_bus1_3 ));
    InMux I__8688 (
            .O(N__36901),
            .I(N__36898));
    LocalMux I__8687 (
            .O(N__36898),
            .I(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0 ));
    InMux I__8686 (
            .O(N__36895),
            .I(N__36892));
    LocalMux I__8685 (
            .O(N__36892),
            .I(N__36889));
    Span12Mux_h I__8684 (
            .O(N__36889),
            .I(N__36886));
    Span12Mux_h I__8683 (
            .O(N__36886),
            .I(N__36883));
    Odrv12 I__8682 (
            .O(N__36883),
            .I(\this_spr_ram.mem_out_bus6_3 ));
    InMux I__8681 (
            .O(N__36880),
            .I(N__36877));
    LocalMux I__8680 (
            .O(N__36877),
            .I(N__36874));
    Span4Mux_h I__8679 (
            .O(N__36874),
            .I(N__36871));
    Span4Mux_v I__8678 (
            .O(N__36871),
            .I(N__36868));
    Odrv4 I__8677 (
            .O(N__36868),
            .I(\this_spr_ram.mem_out_bus2_3 ));
    InMux I__8676 (
            .O(N__36865),
            .I(N__36862));
    LocalMux I__8675 (
            .O(N__36862),
            .I(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0 ));
    InMux I__8674 (
            .O(N__36859),
            .I(N__36856));
    LocalMux I__8673 (
            .O(N__36856),
            .I(N__36853));
    Span4Mux_v I__8672 (
            .O(N__36853),
            .I(N__36850));
    Span4Mux_h I__8671 (
            .O(N__36850),
            .I(N__36847));
    Sp12to4 I__8670 (
            .O(N__36847),
            .I(N__36844));
    Span12Mux_h I__8669 (
            .O(N__36844),
            .I(N__36841));
    Odrv12 I__8668 (
            .O(N__36841),
            .I(\this_spr_ram.mem_out_bus7_0 ));
    InMux I__8667 (
            .O(N__36838),
            .I(N__36835));
    LocalMux I__8666 (
            .O(N__36835),
            .I(N__36832));
    Span4Mux_h I__8665 (
            .O(N__36832),
            .I(N__36829));
    Odrv4 I__8664 (
            .O(N__36829),
            .I(\this_spr_ram.mem_out_bus3_0 ));
    InMux I__8663 (
            .O(N__36826),
            .I(N__36823));
    LocalMux I__8662 (
            .O(N__36823),
            .I(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0 ));
    InMux I__8661 (
            .O(N__36820),
            .I(N__36817));
    LocalMux I__8660 (
            .O(N__36817),
            .I(N__36814));
    Sp12to4 I__8659 (
            .O(N__36814),
            .I(N__36811));
    Span12Mux_v I__8658 (
            .O(N__36811),
            .I(N__36808));
    Span12Mux_h I__8657 (
            .O(N__36808),
            .I(N__36805));
    Odrv12 I__8656 (
            .O(N__36805),
            .I(\this_spr_ram.mem_out_bus7_1 ));
    InMux I__8655 (
            .O(N__36802),
            .I(N__36799));
    LocalMux I__8654 (
            .O(N__36799),
            .I(N__36796));
    Span4Mux_v I__8653 (
            .O(N__36796),
            .I(N__36793));
    Odrv4 I__8652 (
            .O(N__36793),
            .I(\this_spr_ram.mem_out_bus3_1 ));
    InMux I__8651 (
            .O(N__36790),
            .I(N__36787));
    LocalMux I__8650 (
            .O(N__36787),
            .I(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0 ));
    InMux I__8649 (
            .O(N__36784),
            .I(N__36781));
    LocalMux I__8648 (
            .O(N__36781),
            .I(N__36778));
    Span4Mux_h I__8647 (
            .O(N__36778),
            .I(N__36775));
    Sp12to4 I__8646 (
            .O(N__36775),
            .I(N__36772));
    Odrv12 I__8645 (
            .O(N__36772),
            .I(\this_spr_ram.mem_out_bus5_2 ));
    InMux I__8644 (
            .O(N__36769),
            .I(N__36766));
    LocalMux I__8643 (
            .O(N__36766),
            .I(N__36763));
    Span4Mux_h I__8642 (
            .O(N__36763),
            .I(N__36760));
    Span4Mux_v I__8641 (
            .O(N__36760),
            .I(N__36757));
    Odrv4 I__8640 (
            .O(N__36757),
            .I(\this_spr_ram.mem_out_bus1_2 ));
    InMux I__8639 (
            .O(N__36754),
            .I(N__36751));
    LocalMux I__8638 (
            .O(N__36751),
            .I(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0 ));
    InMux I__8637 (
            .O(N__36748),
            .I(N__36745));
    LocalMux I__8636 (
            .O(N__36745),
            .I(N__36742));
    Span4Mux_v I__8635 (
            .O(N__36742),
            .I(N__36739));
    Span4Mux_v I__8634 (
            .O(N__36739),
            .I(N__36736));
    Span4Mux_v I__8633 (
            .O(N__36736),
            .I(N__36733));
    Odrv4 I__8632 (
            .O(N__36733),
            .I(\this_spr_ram.mem_out_bus6_0 ));
    InMux I__8631 (
            .O(N__36730),
            .I(N__36727));
    LocalMux I__8630 (
            .O(N__36727),
            .I(N__36724));
    Span4Mux_v I__8629 (
            .O(N__36724),
            .I(N__36721));
    Span4Mux_v I__8628 (
            .O(N__36721),
            .I(N__36718));
    Odrv4 I__8627 (
            .O(N__36718),
            .I(\this_spr_ram.mem_out_bus2_0 ));
    CascadeMux I__8626 (
            .O(N__36715),
            .I(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_ ));
    InMux I__8625 (
            .O(N__36712),
            .I(N__36709));
    LocalMux I__8624 (
            .O(N__36709),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_0 ));
    CEMux I__8623 (
            .O(N__36706),
            .I(N__36703));
    LocalMux I__8622 (
            .O(N__36703),
            .I(N__36699));
    CEMux I__8621 (
            .O(N__36702),
            .I(N__36696));
    Span4Mux_s2_v I__8620 (
            .O(N__36699),
            .I(N__36691));
    LocalMux I__8619 (
            .O(N__36696),
            .I(N__36691));
    Span4Mux_h I__8618 (
            .O(N__36691),
            .I(N__36688));
    Span4Mux_h I__8617 (
            .O(N__36688),
            .I(N__36685));
    Sp12to4 I__8616 (
            .O(N__36685),
            .I(N__36682));
    Span12Mux_v I__8615 (
            .O(N__36682),
            .I(N__36679));
    Odrv12 I__8614 (
            .O(N__36679),
            .I(\this_spr_ram.mem_WE_0 ));
    InMux I__8613 (
            .O(N__36676),
            .I(N__36673));
    LocalMux I__8612 (
            .O(N__36673),
            .I(N__36670));
    Sp12to4 I__8611 (
            .O(N__36670),
            .I(N__36667));
    Span12Mux_h I__8610 (
            .O(N__36667),
            .I(N__36664));
    Odrv12 I__8609 (
            .O(N__36664),
            .I(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7 ));
    InMux I__8608 (
            .O(N__36661),
            .I(N__36658));
    LocalMux I__8607 (
            .O(N__36658),
            .I(N__36655));
    Span4Mux_v I__8606 (
            .O(N__36655),
            .I(N__36652));
    Span4Mux_h I__8605 (
            .O(N__36652),
            .I(N__36649));
    Sp12to4 I__8604 (
            .O(N__36649),
            .I(N__36646));
    Span12Mux_h I__8603 (
            .O(N__36646),
            .I(N__36643));
    Odrv12 I__8602 (
            .O(N__36643),
            .I(\this_spr_ram.mem_out_bus6_2 ));
    InMux I__8601 (
            .O(N__36640),
            .I(N__36637));
    LocalMux I__8600 (
            .O(N__36637),
            .I(N__36634));
    Span4Mux_h I__8599 (
            .O(N__36634),
            .I(N__36631));
    Odrv4 I__8598 (
            .O(N__36631),
            .I(\this_spr_ram.mem_out_bus2_2 ));
    InMux I__8597 (
            .O(N__36628),
            .I(N__36625));
    LocalMux I__8596 (
            .O(N__36625),
            .I(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0 ));
    InMux I__8595 (
            .O(N__36622),
            .I(N__36619));
    LocalMux I__8594 (
            .O(N__36619),
            .I(N__36616));
    Span4Mux_h I__8593 (
            .O(N__36616),
            .I(N__36613));
    Odrv4 I__8592 (
            .O(N__36613),
            .I(\this_spr_ram.mem_out_bus4_3 ));
    InMux I__8591 (
            .O(N__36610),
            .I(N__36607));
    LocalMux I__8590 (
            .O(N__36607),
            .I(N__36604));
    Span12Mux_h I__8589 (
            .O(N__36604),
            .I(N__36601));
    Span12Mux_v I__8588 (
            .O(N__36601),
            .I(N__36598));
    Odrv12 I__8587 (
            .O(N__36598),
            .I(\this_spr_ram.mem_out_bus0_3 ));
    InMux I__8586 (
            .O(N__36595),
            .I(N__36591));
    InMux I__8585 (
            .O(N__36594),
            .I(N__36588));
    LocalMux I__8584 (
            .O(N__36591),
            .I(N__36585));
    LocalMux I__8583 (
            .O(N__36588),
            .I(N__36582));
    Span12Mux_h I__8582 (
            .O(N__36585),
            .I(N__36579));
    Span4Mux_h I__8581 (
            .O(N__36582),
            .I(N__36576));
    Odrv12 I__8580 (
            .O(N__36579),
            .I(\this_ppu.N_753_0 ));
    Odrv4 I__8579 (
            .O(N__36576),
            .I(\this_ppu.N_753_0 ));
    CascadeMux I__8578 (
            .O(N__36571),
            .I(N__36568));
    InMux I__8577 (
            .O(N__36568),
            .I(N__36564));
    CascadeMux I__8576 (
            .O(N__36567),
            .I(N__36561));
    LocalMux I__8575 (
            .O(N__36564),
            .I(N__36557));
    InMux I__8574 (
            .O(N__36561),
            .I(N__36554));
    InMux I__8573 (
            .O(N__36560),
            .I(N__36551));
    Span4Mux_v I__8572 (
            .O(N__36557),
            .I(N__36548));
    LocalMux I__8571 (
            .O(N__36554),
            .I(N__36543));
    LocalMux I__8570 (
            .O(N__36551),
            .I(N__36543));
    Span4Mux_h I__8569 (
            .O(N__36548),
            .I(N__36538));
    Span4Mux_v I__8568 (
            .O(N__36543),
            .I(N__36538));
    Odrv4 I__8567 (
            .O(N__36538),
            .I(\this_ppu.M_screen_y_qZ0Z_6 ));
    InMux I__8566 (
            .O(N__36535),
            .I(N__36528));
    InMux I__8565 (
            .O(N__36534),
            .I(N__36525));
    InMux I__8564 (
            .O(N__36533),
            .I(N__36522));
    CascadeMux I__8563 (
            .O(N__36532),
            .I(N__36519));
    InMux I__8562 (
            .O(N__36531),
            .I(N__36515));
    LocalMux I__8561 (
            .O(N__36528),
            .I(N__36506));
    LocalMux I__8560 (
            .O(N__36525),
            .I(N__36506));
    LocalMux I__8559 (
            .O(N__36522),
            .I(N__36506));
    InMux I__8558 (
            .O(N__36519),
            .I(N__36503));
    InMux I__8557 (
            .O(N__36518),
            .I(N__36500));
    LocalMux I__8556 (
            .O(N__36515),
            .I(N__36497));
    InMux I__8555 (
            .O(N__36514),
            .I(N__36492));
    InMux I__8554 (
            .O(N__36513),
            .I(N__36492));
    Span4Mux_v I__8553 (
            .O(N__36506),
            .I(N__36485));
    LocalMux I__8552 (
            .O(N__36503),
            .I(N__36485));
    LocalMux I__8551 (
            .O(N__36500),
            .I(N__36485));
    Span4Mux_h I__8550 (
            .O(N__36497),
            .I(N__36479));
    LocalMux I__8549 (
            .O(N__36492),
            .I(N__36479));
    Span4Mux_h I__8548 (
            .O(N__36485),
            .I(N__36473));
    InMux I__8547 (
            .O(N__36484),
            .I(N__36470));
    Span4Mux_v I__8546 (
            .O(N__36479),
            .I(N__36467));
    InMux I__8545 (
            .O(N__36478),
            .I(N__36462));
    InMux I__8544 (
            .O(N__36477),
            .I(N__36462));
    InMux I__8543 (
            .O(N__36476),
            .I(N__36459));
    Span4Mux_h I__8542 (
            .O(N__36473),
            .I(N__36456));
    LocalMux I__8541 (
            .O(N__36470),
            .I(M_this_state_qZ0Z_14));
    Odrv4 I__8540 (
            .O(N__36467),
            .I(M_this_state_qZ0Z_14));
    LocalMux I__8539 (
            .O(N__36462),
            .I(M_this_state_qZ0Z_14));
    LocalMux I__8538 (
            .O(N__36459),
            .I(M_this_state_qZ0Z_14));
    Odrv4 I__8537 (
            .O(N__36456),
            .I(M_this_state_qZ0Z_14));
    InMux I__8536 (
            .O(N__36445),
            .I(N__36439));
    InMux I__8535 (
            .O(N__36444),
            .I(N__36434));
    CascadeMux I__8534 (
            .O(N__36443),
            .I(N__36431));
    CascadeMux I__8533 (
            .O(N__36442),
            .I(N__36427));
    LocalMux I__8532 (
            .O(N__36439),
            .I(N__36424));
    InMux I__8531 (
            .O(N__36438),
            .I(N__36421));
    InMux I__8530 (
            .O(N__36437),
            .I(N__36418));
    LocalMux I__8529 (
            .O(N__36434),
            .I(N__36415));
    InMux I__8528 (
            .O(N__36431),
            .I(N__36412));
    InMux I__8527 (
            .O(N__36430),
            .I(N__36409));
    InMux I__8526 (
            .O(N__36427),
            .I(N__36406));
    Span4Mux_h I__8525 (
            .O(N__36424),
            .I(N__36403));
    LocalMux I__8524 (
            .O(N__36421),
            .I(N__36398));
    LocalMux I__8523 (
            .O(N__36418),
            .I(N__36398));
    Span4Mux_v I__8522 (
            .O(N__36415),
            .I(N__36395));
    LocalMux I__8521 (
            .O(N__36412),
            .I(N__36392));
    LocalMux I__8520 (
            .O(N__36409),
            .I(M_this_state_qZ0Z_13));
    LocalMux I__8519 (
            .O(N__36406),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__8518 (
            .O(N__36403),
            .I(M_this_state_qZ0Z_13));
    Odrv12 I__8517 (
            .O(N__36398),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__8516 (
            .O(N__36395),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__8515 (
            .O(N__36392),
            .I(M_this_state_qZ0Z_13));
    CascadeMux I__8514 (
            .O(N__36379),
            .I(N__36375));
    InMux I__8513 (
            .O(N__36378),
            .I(N__36372));
    InMux I__8512 (
            .O(N__36375),
            .I(N__36369));
    LocalMux I__8511 (
            .O(N__36372),
            .I(N__36364));
    LocalMux I__8510 (
            .O(N__36369),
            .I(N__36364));
    Span12Mux_v I__8509 (
            .O(N__36364),
            .I(N__36361));
    Odrv12 I__8508 (
            .O(N__36361),
            .I(M_this_spr_ram_write_en_0_i_1_0));
    CascadeMux I__8507 (
            .O(N__36358),
            .I(N__36355));
    InMux I__8506 (
            .O(N__36355),
            .I(N__36351));
    InMux I__8505 (
            .O(N__36354),
            .I(N__36347));
    LocalMux I__8504 (
            .O(N__36351),
            .I(N__36344));
    InMux I__8503 (
            .O(N__36350),
            .I(N__36340));
    LocalMux I__8502 (
            .O(N__36347),
            .I(N__36337));
    Span12Mux_h I__8501 (
            .O(N__36344),
            .I(N__36332));
    InMux I__8500 (
            .O(N__36343),
            .I(N__36329));
    LocalMux I__8499 (
            .O(N__36340),
            .I(N__36326));
    Span4Mux_v I__8498 (
            .O(N__36337),
            .I(N__36323));
    InMux I__8497 (
            .O(N__36336),
            .I(N__36318));
    InMux I__8496 (
            .O(N__36335),
            .I(N__36318));
    Odrv12 I__8495 (
            .O(N__36332),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__8494 (
            .O(N__36329),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__8493 (
            .O(N__36326),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__8492 (
            .O(N__36323),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__8491 (
            .O(N__36318),
            .I(M_this_state_qZ0Z_3));
    InMux I__8490 (
            .O(N__36307),
            .I(N__36301));
    InMux I__8489 (
            .O(N__36306),
            .I(N__36301));
    LocalMux I__8488 (
            .O(N__36301),
            .I(N__36295));
    InMux I__8487 (
            .O(N__36300),
            .I(N__36288));
    InMux I__8486 (
            .O(N__36299),
            .I(N__36288));
    InMux I__8485 (
            .O(N__36298),
            .I(N__36288));
    Span4Mux_h I__8484 (
            .O(N__36295),
            .I(N__36282));
    LocalMux I__8483 (
            .O(N__36288),
            .I(N__36282));
    CascadeMux I__8482 (
            .O(N__36287),
            .I(N__36279));
    Span4Mux_v I__8481 (
            .O(N__36282),
            .I(N__36276));
    InMux I__8480 (
            .O(N__36279),
            .I(N__36273));
    Span4Mux_v I__8479 (
            .O(N__36276),
            .I(N__36269));
    LocalMux I__8478 (
            .O(N__36273),
            .I(N__36266));
    InMux I__8477 (
            .O(N__36272),
            .I(N__36263));
    IoSpan4Mux I__8476 (
            .O(N__36269),
            .I(N__36260));
    Span12Mux_h I__8475 (
            .O(N__36266),
            .I(N__36255));
    LocalMux I__8474 (
            .O(N__36263),
            .I(N__36255));
    Odrv4 I__8473 (
            .O(N__36260),
            .I(port_address_in_2));
    Odrv12 I__8472 (
            .O(N__36255),
            .I(port_address_in_2));
    CascadeMux I__8471 (
            .O(N__36250),
            .I(N__36247));
    InMux I__8470 (
            .O(N__36247),
            .I(N__36244));
    LocalMux I__8469 (
            .O(N__36244),
            .I(N__36239));
    InMux I__8468 (
            .O(N__36243),
            .I(N__36236));
    InMux I__8467 (
            .O(N__36242),
            .I(N__36232));
    Span4Mux_v I__8466 (
            .O(N__36239),
            .I(N__36227));
    LocalMux I__8465 (
            .O(N__36236),
            .I(N__36227));
    CascadeMux I__8464 (
            .O(N__36235),
            .I(N__36223));
    LocalMux I__8463 (
            .O(N__36232),
            .I(N__36220));
    Span4Mux_h I__8462 (
            .O(N__36227),
            .I(N__36217));
    InMux I__8461 (
            .O(N__36226),
            .I(N__36214));
    InMux I__8460 (
            .O(N__36223),
            .I(N__36211));
    Span4Mux_v I__8459 (
            .O(N__36220),
            .I(N__36207));
    Span4Mux_h I__8458 (
            .O(N__36217),
            .I(N__36200));
    LocalMux I__8457 (
            .O(N__36214),
            .I(N__36200));
    LocalMux I__8456 (
            .O(N__36211),
            .I(N__36200));
    CascadeMux I__8455 (
            .O(N__36210),
            .I(N__36197));
    Span4Mux_h I__8454 (
            .O(N__36207),
            .I(N__36192));
    Span4Mux_v I__8453 (
            .O(N__36200),
            .I(N__36189));
    InMux I__8452 (
            .O(N__36197),
            .I(N__36186));
    InMux I__8451 (
            .O(N__36196),
            .I(N__36181));
    InMux I__8450 (
            .O(N__36195),
            .I(N__36181));
    Sp12to4 I__8449 (
            .O(N__36192),
            .I(N__36178));
    Span4Mux_h I__8448 (
            .O(N__36189),
            .I(N__36175));
    LocalMux I__8447 (
            .O(N__36186),
            .I(N__36170));
    LocalMux I__8446 (
            .O(N__36181),
            .I(N__36170));
    Span12Mux_s6_h I__8445 (
            .O(N__36178),
            .I(N__36163));
    Sp12to4 I__8444 (
            .O(N__36175),
            .I(N__36163));
    Span12Mux_h I__8443 (
            .O(N__36170),
            .I(N__36163));
    Odrv12 I__8442 (
            .O(N__36163),
            .I(port_address_in_1));
    InMux I__8441 (
            .O(N__36160),
            .I(N__36157));
    LocalMux I__8440 (
            .O(N__36157),
            .I(N__36149));
    InMux I__8439 (
            .O(N__36156),
            .I(N__36146));
    InMux I__8438 (
            .O(N__36155),
            .I(N__36141));
    InMux I__8437 (
            .O(N__36154),
            .I(N__36141));
    InMux I__8436 (
            .O(N__36153),
            .I(N__36138));
    InMux I__8435 (
            .O(N__36152),
            .I(N__36135));
    Odrv4 I__8434 (
            .O(N__36149),
            .I(M_this_substate_qZ0));
    LocalMux I__8433 (
            .O(N__36146),
            .I(M_this_substate_qZ0));
    LocalMux I__8432 (
            .O(N__36141),
            .I(M_this_substate_qZ0));
    LocalMux I__8431 (
            .O(N__36138),
            .I(M_this_substate_qZ0));
    LocalMux I__8430 (
            .O(N__36135),
            .I(M_this_substate_qZ0));
    InMux I__8429 (
            .O(N__36124),
            .I(N__36121));
    LocalMux I__8428 (
            .O(N__36121),
            .I(this_ppu_M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1));
    CascadeMux I__8427 (
            .O(N__36118),
            .I(M_this_map_address_qc_3_0_cascade_));
    InMux I__8426 (
            .O(N__36115),
            .I(N__36110));
    CascadeMux I__8425 (
            .O(N__36114),
            .I(N__36107));
    InMux I__8424 (
            .O(N__36113),
            .I(N__36104));
    LocalMux I__8423 (
            .O(N__36110),
            .I(N__36101));
    InMux I__8422 (
            .O(N__36107),
            .I(N__36096));
    LocalMux I__8421 (
            .O(N__36104),
            .I(N__36091));
    Span4Mux_h I__8420 (
            .O(N__36101),
            .I(N__36091));
    InMux I__8419 (
            .O(N__36100),
            .I(N__36088));
    InMux I__8418 (
            .O(N__36099),
            .I(N__36085));
    LocalMux I__8417 (
            .O(N__36096),
            .I(M_this_state_qZ0Z_10));
    Odrv4 I__8416 (
            .O(N__36091),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__8415 (
            .O(N__36088),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__8414 (
            .O(N__36085),
            .I(M_this_state_qZ0Z_10));
    InMux I__8413 (
            .O(N__36076),
            .I(N__36073));
    LocalMux I__8412 (
            .O(N__36073),
            .I(N__36070));
    Span4Mux_h I__8411 (
            .O(N__36070),
            .I(N__36067));
    Odrv4 I__8410 (
            .O(N__36067),
            .I(N_169_0));
    IoInMux I__8409 (
            .O(N__36064),
            .I(N__36061));
    LocalMux I__8408 (
            .O(N__36061),
            .I(N__36058));
    IoSpan4Mux I__8407 (
            .O(N__36058),
            .I(N__36055));
    IoSpan4Mux I__8406 (
            .O(N__36055),
            .I(N__36052));
    Span4Mux_s1_h I__8405 (
            .O(N__36052),
            .I(N__36049));
    Span4Mux_h I__8404 (
            .O(N__36049),
            .I(N__36046));
    Odrv4 I__8403 (
            .O(N__36046),
            .I(N_1048_i));
    InMux I__8402 (
            .O(N__36043),
            .I(N__36040));
    LocalMux I__8401 (
            .O(N__36040),
            .I(N__36037));
    Span4Mux_h I__8400 (
            .O(N__36037),
            .I(N__36034));
    Span4Mux_v I__8399 (
            .O(N__36034),
            .I(N__36031));
    Odrv4 I__8398 (
            .O(N__36031),
            .I(\this_spr_ram.mem_out_bus5_1 ));
    InMux I__8397 (
            .O(N__36028),
            .I(N__36025));
    LocalMux I__8396 (
            .O(N__36025),
            .I(N__36022));
    Span4Mux_v I__8395 (
            .O(N__36022),
            .I(N__36019));
    Span4Mux_v I__8394 (
            .O(N__36019),
            .I(N__36016));
    Odrv4 I__8393 (
            .O(N__36016),
            .I(\this_spr_ram.mem_out_bus1_1 ));
    InMux I__8392 (
            .O(N__36013),
            .I(N__36010));
    LocalMux I__8391 (
            .O(N__36010),
            .I(N__36007));
    Span4Mux_v I__8390 (
            .O(N__36007),
            .I(N__36004));
    Odrv4 I__8389 (
            .O(N__36004),
            .I(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0 ));
    InMux I__8388 (
            .O(N__36001),
            .I(N__35995));
    InMux I__8387 (
            .O(N__36000),
            .I(N__35995));
    LocalMux I__8386 (
            .O(N__35995),
            .I(\this_ppu.N_1257 ));
    InMux I__8385 (
            .O(N__35992),
            .I(N__35989));
    LocalMux I__8384 (
            .O(N__35989),
            .I(N__35985));
    InMux I__8383 (
            .O(N__35988),
            .I(N__35982));
    Span4Mux_v I__8382 (
            .O(N__35985),
            .I(N__35977));
    LocalMux I__8381 (
            .O(N__35982),
            .I(N__35977));
    Span4Mux_h I__8380 (
            .O(N__35977),
            .I(N__35973));
    InMux I__8379 (
            .O(N__35976),
            .I(N__35970));
    Odrv4 I__8378 (
            .O(N__35973),
            .I(\this_ppu.N_1322 ));
    LocalMux I__8377 (
            .O(N__35970),
            .I(\this_ppu.N_1322 ));
    InMux I__8376 (
            .O(N__35965),
            .I(N__35961));
    InMux I__8375 (
            .O(N__35964),
            .I(N__35957));
    LocalMux I__8374 (
            .O(N__35961),
            .I(N__35954));
    InMux I__8373 (
            .O(N__35960),
            .I(N__35951));
    LocalMux I__8372 (
            .O(N__35957),
            .I(N__35946));
    Span4Mux_h I__8371 (
            .O(N__35954),
            .I(N__35943));
    LocalMux I__8370 (
            .O(N__35951),
            .I(N__35940));
    InMux I__8369 (
            .O(N__35950),
            .I(N__35937));
    InMux I__8368 (
            .O(N__35949),
            .I(N__35933));
    Span4Mux_v I__8367 (
            .O(N__35946),
            .I(N__35930));
    Span4Mux_v I__8366 (
            .O(N__35943),
            .I(N__35925));
    Span4Mux_h I__8365 (
            .O(N__35940),
            .I(N__35925));
    LocalMux I__8364 (
            .O(N__35937),
            .I(N__35922));
    InMux I__8363 (
            .O(N__35936),
            .I(N__35919));
    LocalMux I__8362 (
            .O(N__35933),
            .I(N__35915));
    Span4Mux_v I__8361 (
            .O(N__35930),
            .I(N__35911));
    Span4Mux_v I__8360 (
            .O(N__35925),
            .I(N__35906));
    Span4Mux_h I__8359 (
            .O(N__35922),
            .I(N__35906));
    LocalMux I__8358 (
            .O(N__35919),
            .I(N__35903));
    InMux I__8357 (
            .O(N__35918),
            .I(N__35900));
    Span4Mux_h I__8356 (
            .O(N__35915),
            .I(N__35897));
    InMux I__8355 (
            .O(N__35914),
            .I(N__35894));
    Sp12to4 I__8354 (
            .O(N__35911),
            .I(N__35891));
    Span4Mux_v I__8353 (
            .O(N__35906),
            .I(N__35886));
    Span4Mux_h I__8352 (
            .O(N__35903),
            .I(N__35886));
    LocalMux I__8351 (
            .O(N__35900),
            .I(N__35883));
    Span4Mux_v I__8350 (
            .O(N__35897),
            .I(N__35878));
    LocalMux I__8349 (
            .O(N__35894),
            .I(N__35878));
    Span12Mux_h I__8348 (
            .O(N__35891),
            .I(N__35875));
    Span4Mux_v I__8347 (
            .O(N__35886),
            .I(N__35868));
    Span4Mux_h I__8346 (
            .O(N__35883),
            .I(N__35868));
    Span4Mux_h I__8345 (
            .O(N__35878),
            .I(N__35868));
    Odrv12 I__8344 (
            .O(N__35875),
            .I(M_this_spr_ram_write_data_1));
    Odrv4 I__8343 (
            .O(N__35868),
            .I(M_this_spr_ram_write_data_1));
    IoInMux I__8342 (
            .O(N__35863),
            .I(N__35860));
    LocalMux I__8341 (
            .O(N__35860),
            .I(N__35857));
    Span4Mux_s3_h I__8340 (
            .O(N__35857),
            .I(N__35854));
    Span4Mux_h I__8339 (
            .O(N__35854),
            .I(N__35851));
    Span4Mux_h I__8338 (
            .O(N__35851),
            .I(N__35848));
    Sp12to4 I__8337 (
            .O(N__35848),
            .I(N__35842));
    InMux I__8336 (
            .O(N__35847),
            .I(N__35834));
    InMux I__8335 (
            .O(N__35846),
            .I(N__35834));
    InMux I__8334 (
            .O(N__35845),
            .I(N__35831));
    Span12Mux_v I__8333 (
            .O(N__35842),
            .I(N__35827));
    InMux I__8332 (
            .O(N__35841),
            .I(N__35822));
    InMux I__8331 (
            .O(N__35840),
            .I(N__35822));
    InMux I__8330 (
            .O(N__35839),
            .I(N__35819));
    LocalMux I__8329 (
            .O(N__35834),
            .I(N__35814));
    LocalMux I__8328 (
            .O(N__35831),
            .I(N__35814));
    InMux I__8327 (
            .O(N__35830),
            .I(N__35811));
    Odrv12 I__8326 (
            .O(N__35827),
            .I(led_c_1));
    LocalMux I__8325 (
            .O(N__35822),
            .I(led_c_1));
    LocalMux I__8324 (
            .O(N__35819),
            .I(led_c_1));
    Odrv4 I__8323 (
            .O(N__35814),
            .I(led_c_1));
    LocalMux I__8322 (
            .O(N__35811),
            .I(led_c_1));
    CascadeMux I__8321 (
            .O(N__35800),
            .I(N_1416_cascade_));
    CascadeMux I__8320 (
            .O(N__35797),
            .I(N__35794));
    InMux I__8319 (
            .O(N__35794),
            .I(N__35788));
    InMux I__8318 (
            .O(N__35793),
            .I(N__35788));
    LocalMux I__8317 (
            .O(N__35788),
            .I(N_1151_3));
    InMux I__8316 (
            .O(N__35785),
            .I(N__35778));
    InMux I__8315 (
            .O(N__35784),
            .I(N__35774));
    InMux I__8314 (
            .O(N__35783),
            .I(N__35770));
    InMux I__8313 (
            .O(N__35782),
            .I(N__35767));
    InMux I__8312 (
            .O(N__35781),
            .I(N__35764));
    LocalMux I__8311 (
            .O(N__35778),
            .I(N__35760));
    InMux I__8310 (
            .O(N__35777),
            .I(N__35757));
    LocalMux I__8309 (
            .O(N__35774),
            .I(N__35754));
    InMux I__8308 (
            .O(N__35773),
            .I(N__35751));
    LocalMux I__8307 (
            .O(N__35770),
            .I(N__35748));
    LocalMux I__8306 (
            .O(N__35767),
            .I(N__35743));
    LocalMux I__8305 (
            .O(N__35764),
            .I(N__35743));
    InMux I__8304 (
            .O(N__35763),
            .I(N__35740));
    Span4Mux_h I__8303 (
            .O(N__35760),
            .I(N__35733));
    LocalMux I__8302 (
            .O(N__35757),
            .I(N__35733));
    Span4Mux_v I__8301 (
            .O(N__35754),
            .I(N__35733));
    LocalMux I__8300 (
            .O(N__35751),
            .I(N__35726));
    Span4Mux_v I__8299 (
            .O(N__35748),
            .I(N__35726));
    Span4Mux_v I__8298 (
            .O(N__35743),
            .I(N__35726));
    LocalMux I__8297 (
            .O(N__35740),
            .I(\this_ppu.N_787_0 ));
    Odrv4 I__8296 (
            .O(N__35733),
            .I(\this_ppu.N_787_0 ));
    Odrv4 I__8295 (
            .O(N__35726),
            .I(\this_ppu.N_787_0 ));
    InMux I__8294 (
            .O(N__35719),
            .I(N__35716));
    LocalMux I__8293 (
            .O(N__35716),
            .I(\this_ppu.M_this_state_q_srsts_0_0_a2_1_sxZ0Z_0 ));
    CascadeMux I__8292 (
            .O(N__35713),
            .I(N__35706));
    InMux I__8291 (
            .O(N__35712),
            .I(N__35698));
    InMux I__8290 (
            .O(N__35711),
            .I(N__35698));
    InMux I__8289 (
            .O(N__35710),
            .I(N__35698));
    InMux I__8288 (
            .O(N__35709),
            .I(N__35693));
    InMux I__8287 (
            .O(N__35706),
            .I(N__35693));
    CascadeMux I__8286 (
            .O(N__35705),
            .I(N__35690));
    LocalMux I__8285 (
            .O(N__35698),
            .I(N__35685));
    LocalMux I__8284 (
            .O(N__35693),
            .I(N__35685));
    InMux I__8283 (
            .O(N__35690),
            .I(N__35681));
    Span4Mux_h I__8282 (
            .O(N__35685),
            .I(N__35678));
    InMux I__8281 (
            .O(N__35684),
            .I(N__35675));
    LocalMux I__8280 (
            .O(N__35681),
            .I(N__35672));
    Odrv4 I__8279 (
            .O(N__35678),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__8278 (
            .O(N__35675),
            .I(\this_vga_signals.vaddress_6 ));
    Odrv4 I__8277 (
            .O(N__35672),
            .I(\this_vga_signals.vaddress_6 ));
    InMux I__8276 (
            .O(N__35665),
            .I(N__35660));
    InMux I__8275 (
            .O(N__35664),
            .I(N__35657));
    InMux I__8274 (
            .O(N__35663),
            .I(N__35653));
    LocalMux I__8273 (
            .O(N__35660),
            .I(N__35648));
    LocalMux I__8272 (
            .O(N__35657),
            .I(N__35648));
    InMux I__8271 (
            .O(N__35656),
            .I(N__35645));
    LocalMux I__8270 (
            .O(N__35653),
            .I(N__35642));
    Span4Mux_h I__8269 (
            .O(N__35648),
            .I(N__35637));
    LocalMux I__8268 (
            .O(N__35645),
            .I(N__35637));
    Span4Mux_h I__8267 (
            .O(N__35642),
            .I(N__35634));
    Odrv4 I__8266 (
            .O(N__35637),
            .I(\this_vga_signals.vaddress_5 ));
    Odrv4 I__8265 (
            .O(N__35634),
            .I(\this_vga_signals.vaddress_5 ));
    CascadeMux I__8264 (
            .O(N__35629),
            .I(N__35626));
    InMux I__8263 (
            .O(N__35626),
            .I(N__35623));
    LocalMux I__8262 (
            .O(N__35623),
            .I(N__35620));
    Odrv4 I__8261 (
            .O(N__35620),
            .I(\this_vga_signals.g2_1_0 ));
    CascadeMux I__8260 (
            .O(N__35617),
            .I(N__35612));
    CascadeMux I__8259 (
            .O(N__35616),
            .I(N__35605));
    InMux I__8258 (
            .O(N__35615),
            .I(N__35595));
    InMux I__8257 (
            .O(N__35612),
            .I(N__35595));
    InMux I__8256 (
            .O(N__35611),
            .I(N__35595));
    InMux I__8255 (
            .O(N__35610),
            .I(N__35592));
    InMux I__8254 (
            .O(N__35609),
            .I(N__35587));
    InMux I__8253 (
            .O(N__35608),
            .I(N__35587));
    InMux I__8252 (
            .O(N__35605),
            .I(N__35582));
    InMux I__8251 (
            .O(N__35604),
            .I(N__35582));
    InMux I__8250 (
            .O(N__35603),
            .I(N__35577));
    InMux I__8249 (
            .O(N__35602),
            .I(N__35577));
    LocalMux I__8248 (
            .O(N__35595),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_4 ));
    LocalMux I__8247 (
            .O(N__35592),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_4 ));
    LocalMux I__8246 (
            .O(N__35587),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_4 ));
    LocalMux I__8245 (
            .O(N__35582),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_4 ));
    LocalMux I__8244 (
            .O(N__35577),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_4 ));
    InMux I__8243 (
            .O(N__35566),
            .I(N__35563));
    LocalMux I__8242 (
            .O(N__35563),
            .I(N__35560));
    Odrv12 I__8241 (
            .O(N__35560),
            .I(\this_vga_signals.mult1_un47_sum_2_1 ));
    InMux I__8240 (
            .O(N__35557),
            .I(N__35554));
    LocalMux I__8239 (
            .O(N__35554),
            .I(N__35549));
    InMux I__8238 (
            .O(N__35553),
            .I(N__35545));
    InMux I__8237 (
            .O(N__35552),
            .I(N__35542));
    Span4Mux_h I__8236 (
            .O(N__35549),
            .I(N__35539));
    InMux I__8235 (
            .O(N__35548),
            .I(N__35536));
    LocalMux I__8234 (
            .O(N__35545),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__8233 (
            .O(N__35542),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    Odrv4 I__8232 (
            .O(N__35539),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__8231 (
            .O(N__35536),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    InMux I__8230 (
            .O(N__35527),
            .I(N__35524));
    LocalMux I__8229 (
            .O(N__35524),
            .I(\this_vga_signals.if_N_7_0_0 ));
    CascadeMux I__8228 (
            .O(N__35521),
            .I(N__35511));
    CascadeMux I__8227 (
            .O(N__35520),
            .I(N__35508));
    CascadeMux I__8226 (
            .O(N__35519),
            .I(N__35505));
    InMux I__8225 (
            .O(N__35518),
            .I(N__35498));
    InMux I__8224 (
            .O(N__35517),
            .I(N__35498));
    InMux I__8223 (
            .O(N__35516),
            .I(N__35498));
    InMux I__8222 (
            .O(N__35515),
            .I(N__35495));
    InMux I__8221 (
            .O(N__35514),
            .I(N__35492));
    InMux I__8220 (
            .O(N__35511),
            .I(N__35486));
    InMux I__8219 (
            .O(N__35508),
            .I(N__35483));
    InMux I__8218 (
            .O(N__35505),
            .I(N__35480));
    LocalMux I__8217 (
            .O(N__35498),
            .I(N__35477));
    LocalMux I__8216 (
            .O(N__35495),
            .I(N__35472));
    LocalMux I__8215 (
            .O(N__35492),
            .I(N__35472));
    CascadeMux I__8214 (
            .O(N__35491),
            .I(N__35469));
    CascadeMux I__8213 (
            .O(N__35490),
            .I(N__35466));
    InMux I__8212 (
            .O(N__35489),
            .I(N__35461));
    LocalMux I__8211 (
            .O(N__35486),
            .I(N__35453));
    LocalMux I__8210 (
            .O(N__35483),
            .I(N__35453));
    LocalMux I__8209 (
            .O(N__35480),
            .I(N__35453));
    Span4Mux_h I__8208 (
            .O(N__35477),
            .I(N__35448));
    Span4Mux_h I__8207 (
            .O(N__35472),
            .I(N__35448));
    InMux I__8206 (
            .O(N__35469),
            .I(N__35443));
    InMux I__8205 (
            .O(N__35466),
            .I(N__35443));
    InMux I__8204 (
            .O(N__35465),
            .I(N__35440));
    InMux I__8203 (
            .O(N__35464),
            .I(N__35437));
    LocalMux I__8202 (
            .O(N__35461),
            .I(N__35434));
    InMux I__8201 (
            .O(N__35460),
            .I(N__35431));
    Span12Mux_h I__8200 (
            .O(N__35453),
            .I(N__35426));
    Sp12to4 I__8199 (
            .O(N__35448),
            .I(N__35426));
    LocalMux I__8198 (
            .O(N__35443),
            .I(N__35423));
    LocalMux I__8197 (
            .O(N__35440),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__8196 (
            .O(N__35437),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__8195 (
            .O(N__35434),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__8194 (
            .O(N__35431),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv12 I__8193 (
            .O(N__35426),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__8192 (
            .O(N__35423),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    InMux I__8191 (
            .O(N__35410),
            .I(N__35402));
    InMux I__8190 (
            .O(N__35409),
            .I(N__35393));
    InMux I__8189 (
            .O(N__35408),
            .I(N__35393));
    InMux I__8188 (
            .O(N__35407),
            .I(N__35387));
    InMux I__8187 (
            .O(N__35406),
            .I(N__35387));
    CascadeMux I__8186 (
            .O(N__35405),
            .I(N__35381));
    LocalMux I__8185 (
            .O(N__35402),
            .I(N__35377));
    InMux I__8184 (
            .O(N__35401),
            .I(N__35370));
    InMux I__8183 (
            .O(N__35400),
            .I(N__35370));
    InMux I__8182 (
            .O(N__35399),
            .I(N__35370));
    InMux I__8181 (
            .O(N__35398),
            .I(N__35367));
    LocalMux I__8180 (
            .O(N__35393),
            .I(N__35364));
    InMux I__8179 (
            .O(N__35392),
            .I(N__35361));
    LocalMux I__8178 (
            .O(N__35387),
            .I(N__35358));
    InMux I__8177 (
            .O(N__35386),
            .I(N__35353));
    InMux I__8176 (
            .O(N__35385),
            .I(N__35353));
    InMux I__8175 (
            .O(N__35384),
            .I(N__35346));
    InMux I__8174 (
            .O(N__35381),
            .I(N__35346));
    InMux I__8173 (
            .O(N__35380),
            .I(N__35346));
    Odrv4 I__8172 (
            .O(N__35377),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__8171 (
            .O(N__35370),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__8170 (
            .O(N__35367),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv12 I__8169 (
            .O(N__35364),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__8168 (
            .O(N__35361),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__8167 (
            .O(N__35358),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__8166 (
            .O(N__35353),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__8165 (
            .O(N__35346),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    InMux I__8164 (
            .O(N__35329),
            .I(N__35326));
    LocalMux I__8163 (
            .O(N__35326),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d_0_0 ));
    InMux I__8162 (
            .O(N__35323),
            .I(N__35311));
    InMux I__8161 (
            .O(N__35322),
            .I(N__35308));
    InMux I__8160 (
            .O(N__35321),
            .I(N__35297));
    InMux I__8159 (
            .O(N__35320),
            .I(N__35294));
    InMux I__8158 (
            .O(N__35319),
            .I(N__35290));
    InMux I__8157 (
            .O(N__35318),
            .I(N__35287));
    InMux I__8156 (
            .O(N__35317),
            .I(N__35279));
    InMux I__8155 (
            .O(N__35316),
            .I(N__35279));
    InMux I__8154 (
            .O(N__35315),
            .I(N__35279));
    InMux I__8153 (
            .O(N__35314),
            .I(N__35276));
    LocalMux I__8152 (
            .O(N__35311),
            .I(N__35271));
    LocalMux I__8151 (
            .O(N__35308),
            .I(N__35271));
    InMux I__8150 (
            .O(N__35307),
            .I(N__35266));
    InMux I__8149 (
            .O(N__35306),
            .I(N__35266));
    InMux I__8148 (
            .O(N__35305),
            .I(N__35263));
    InMux I__8147 (
            .O(N__35304),
            .I(N__35260));
    InMux I__8146 (
            .O(N__35303),
            .I(N__35257));
    InMux I__8145 (
            .O(N__35302),
            .I(N__35252));
    InMux I__8144 (
            .O(N__35301),
            .I(N__35252));
    CascadeMux I__8143 (
            .O(N__35300),
            .I(N__35249));
    LocalMux I__8142 (
            .O(N__35297),
            .I(N__35245));
    LocalMux I__8141 (
            .O(N__35294),
            .I(N__35242));
    CascadeMux I__8140 (
            .O(N__35293),
            .I(N__35237));
    LocalMux I__8139 (
            .O(N__35290),
            .I(N__35232));
    LocalMux I__8138 (
            .O(N__35287),
            .I(N__35232));
    InMux I__8137 (
            .O(N__35286),
            .I(N__35229));
    LocalMux I__8136 (
            .O(N__35279),
            .I(N__35220));
    LocalMux I__8135 (
            .O(N__35276),
            .I(N__35220));
    Span4Mux_v I__8134 (
            .O(N__35271),
            .I(N__35220));
    LocalMux I__8133 (
            .O(N__35266),
            .I(N__35220));
    LocalMux I__8132 (
            .O(N__35263),
            .I(N__35216));
    LocalMux I__8131 (
            .O(N__35260),
            .I(N__35211));
    LocalMux I__8130 (
            .O(N__35257),
            .I(N__35211));
    LocalMux I__8129 (
            .O(N__35252),
            .I(N__35208));
    InMux I__8128 (
            .O(N__35249),
            .I(N__35205));
    InMux I__8127 (
            .O(N__35248),
            .I(N__35202));
    Span4Mux_v I__8126 (
            .O(N__35245),
            .I(N__35197));
    Span4Mux_v I__8125 (
            .O(N__35242),
            .I(N__35197));
    InMux I__8124 (
            .O(N__35241),
            .I(N__35190));
    InMux I__8123 (
            .O(N__35240),
            .I(N__35190));
    InMux I__8122 (
            .O(N__35237),
            .I(N__35190));
    Sp12to4 I__8121 (
            .O(N__35232),
            .I(N__35185));
    LocalMux I__8120 (
            .O(N__35229),
            .I(N__35185));
    Span4Mux_h I__8119 (
            .O(N__35220),
            .I(N__35182));
    InMux I__8118 (
            .O(N__35219),
            .I(N__35179));
    Span4Mux_h I__8117 (
            .O(N__35216),
            .I(N__35170));
    Span4Mux_h I__8116 (
            .O(N__35211),
            .I(N__35170));
    Span4Mux_h I__8115 (
            .O(N__35208),
            .I(N__35170));
    LocalMux I__8114 (
            .O(N__35205),
            .I(N__35170));
    LocalMux I__8113 (
            .O(N__35202),
            .I(this_vga_signals_M_vcounter_q_4));
    Odrv4 I__8112 (
            .O(N__35197),
            .I(this_vga_signals_M_vcounter_q_4));
    LocalMux I__8111 (
            .O(N__35190),
            .I(this_vga_signals_M_vcounter_q_4));
    Odrv12 I__8110 (
            .O(N__35185),
            .I(this_vga_signals_M_vcounter_q_4));
    Odrv4 I__8109 (
            .O(N__35182),
            .I(this_vga_signals_M_vcounter_q_4));
    LocalMux I__8108 (
            .O(N__35179),
            .I(this_vga_signals_M_vcounter_q_4));
    Odrv4 I__8107 (
            .O(N__35170),
            .I(this_vga_signals_M_vcounter_q_4));
    CascadeMux I__8106 (
            .O(N__35155),
            .I(N__35147));
    CascadeMux I__8105 (
            .O(N__35154),
            .I(N__35143));
    InMux I__8104 (
            .O(N__35153),
            .I(N__35138));
    InMux I__8103 (
            .O(N__35152),
            .I(N__35130));
    InMux I__8102 (
            .O(N__35151),
            .I(N__35127));
    InMux I__8101 (
            .O(N__35150),
            .I(N__35124));
    InMux I__8100 (
            .O(N__35147),
            .I(N__35121));
    InMux I__8099 (
            .O(N__35146),
            .I(N__35118));
    InMux I__8098 (
            .O(N__35143),
            .I(N__35115));
    InMux I__8097 (
            .O(N__35142),
            .I(N__35110));
    InMux I__8096 (
            .O(N__35141),
            .I(N__35110));
    LocalMux I__8095 (
            .O(N__35138),
            .I(N__35107));
    InMux I__8094 (
            .O(N__35137),
            .I(N__35104));
    CascadeMux I__8093 (
            .O(N__35136),
            .I(N__35101));
    CascadeMux I__8092 (
            .O(N__35135),
            .I(N__35096));
    InMux I__8091 (
            .O(N__35134),
            .I(N__35093));
    CascadeMux I__8090 (
            .O(N__35133),
            .I(N__35090));
    LocalMux I__8089 (
            .O(N__35130),
            .I(N__35086));
    LocalMux I__8088 (
            .O(N__35127),
            .I(N__35079));
    LocalMux I__8087 (
            .O(N__35124),
            .I(N__35079));
    LocalMux I__8086 (
            .O(N__35121),
            .I(N__35079));
    LocalMux I__8085 (
            .O(N__35118),
            .I(N__35076));
    LocalMux I__8084 (
            .O(N__35115),
            .I(N__35072));
    LocalMux I__8083 (
            .O(N__35110),
            .I(N__35065));
    Span4Mux_v I__8082 (
            .O(N__35107),
            .I(N__35065));
    LocalMux I__8081 (
            .O(N__35104),
            .I(N__35065));
    InMux I__8080 (
            .O(N__35101),
            .I(N__35060));
    InMux I__8079 (
            .O(N__35100),
            .I(N__35060));
    InMux I__8078 (
            .O(N__35099),
            .I(N__35057));
    InMux I__8077 (
            .O(N__35096),
            .I(N__35054));
    LocalMux I__8076 (
            .O(N__35093),
            .I(N__35051));
    InMux I__8075 (
            .O(N__35090),
            .I(N__35046));
    InMux I__8074 (
            .O(N__35089),
            .I(N__35046));
    Span4Mux_v I__8073 (
            .O(N__35086),
            .I(N__35039));
    Span4Mux_h I__8072 (
            .O(N__35079),
            .I(N__35039));
    Span4Mux_v I__8071 (
            .O(N__35076),
            .I(N__35039));
    InMux I__8070 (
            .O(N__35075),
            .I(N__35036));
    Span4Mux_h I__8069 (
            .O(N__35072),
            .I(N__35029));
    Span4Mux_h I__8068 (
            .O(N__35065),
            .I(N__35029));
    LocalMux I__8067 (
            .O(N__35060),
            .I(N__35029));
    LocalMux I__8066 (
            .O(N__35057),
            .I(this_vga_signals_M_vcounter_q_7));
    LocalMux I__8065 (
            .O(N__35054),
            .I(this_vga_signals_M_vcounter_q_7));
    Odrv4 I__8064 (
            .O(N__35051),
            .I(this_vga_signals_M_vcounter_q_7));
    LocalMux I__8063 (
            .O(N__35046),
            .I(this_vga_signals_M_vcounter_q_7));
    Odrv4 I__8062 (
            .O(N__35039),
            .I(this_vga_signals_M_vcounter_q_7));
    LocalMux I__8061 (
            .O(N__35036),
            .I(this_vga_signals_M_vcounter_q_7));
    Odrv4 I__8060 (
            .O(N__35029),
            .I(this_vga_signals_M_vcounter_q_7));
    InMux I__8059 (
            .O(N__35014),
            .I(N__35009));
    CascadeMux I__8058 (
            .O(N__35013),
            .I(N__35006));
    InMux I__8057 (
            .O(N__35012),
            .I(N__35001));
    LocalMux I__8056 (
            .O(N__35009),
            .I(N__34996));
    InMux I__8055 (
            .O(N__35006),
            .I(N__34987));
    CascadeMux I__8054 (
            .O(N__35005),
            .I(N__34983));
    InMux I__8053 (
            .O(N__35004),
            .I(N__34980));
    LocalMux I__8052 (
            .O(N__35001),
            .I(N__34977));
    InMux I__8051 (
            .O(N__35000),
            .I(N__34974));
    CascadeMux I__8050 (
            .O(N__34999),
            .I(N__34968));
    Span4Mux_h I__8049 (
            .O(N__34996),
            .I(N__34963));
    InMux I__8048 (
            .O(N__34995),
            .I(N__34960));
    InMux I__8047 (
            .O(N__34994),
            .I(N__34955));
    InMux I__8046 (
            .O(N__34993),
            .I(N__34955));
    InMux I__8045 (
            .O(N__34992),
            .I(N__34948));
    InMux I__8044 (
            .O(N__34991),
            .I(N__34948));
    InMux I__8043 (
            .O(N__34990),
            .I(N__34948));
    LocalMux I__8042 (
            .O(N__34987),
            .I(N__34939));
    InMux I__8041 (
            .O(N__34986),
            .I(N__34935));
    InMux I__8040 (
            .O(N__34983),
            .I(N__34932));
    LocalMux I__8039 (
            .O(N__34980),
            .I(N__34929));
    Span4Mux_h I__8038 (
            .O(N__34977),
            .I(N__34924));
    LocalMux I__8037 (
            .O(N__34974),
            .I(N__34924));
    InMux I__8036 (
            .O(N__34973),
            .I(N__34921));
    InMux I__8035 (
            .O(N__34972),
            .I(N__34916));
    InMux I__8034 (
            .O(N__34971),
            .I(N__34916));
    InMux I__8033 (
            .O(N__34968),
            .I(N__34913));
    InMux I__8032 (
            .O(N__34967),
            .I(N__34908));
    InMux I__8031 (
            .O(N__34966),
            .I(N__34908));
    Span4Mux_h I__8030 (
            .O(N__34963),
            .I(N__34901));
    LocalMux I__8029 (
            .O(N__34960),
            .I(N__34901));
    LocalMux I__8028 (
            .O(N__34955),
            .I(N__34901));
    LocalMux I__8027 (
            .O(N__34948),
            .I(N__34898));
    InMux I__8026 (
            .O(N__34947),
            .I(N__34894));
    CascadeMux I__8025 (
            .O(N__34946),
            .I(N__34891));
    CascadeMux I__8024 (
            .O(N__34945),
            .I(N__34888));
    CascadeMux I__8023 (
            .O(N__34944),
            .I(N__34885));
    CascadeMux I__8022 (
            .O(N__34943),
            .I(N__34882));
    CascadeMux I__8021 (
            .O(N__34942),
            .I(N__34876));
    Span4Mux_v I__8020 (
            .O(N__34939),
            .I(N__34873));
    CascadeMux I__8019 (
            .O(N__34938),
            .I(N__34870));
    LocalMux I__8018 (
            .O(N__34935),
            .I(N__34865));
    LocalMux I__8017 (
            .O(N__34932),
            .I(N__34865));
    Span4Mux_v I__8016 (
            .O(N__34929),
            .I(N__34858));
    Span4Mux_v I__8015 (
            .O(N__34924),
            .I(N__34858));
    LocalMux I__8014 (
            .O(N__34921),
            .I(N__34858));
    LocalMux I__8013 (
            .O(N__34916),
            .I(N__34855));
    LocalMux I__8012 (
            .O(N__34913),
            .I(N__34846));
    LocalMux I__8011 (
            .O(N__34908),
            .I(N__34846));
    Span4Mux_h I__8010 (
            .O(N__34901),
            .I(N__34846));
    Span4Mux_v I__8009 (
            .O(N__34898),
            .I(N__34846));
    CascadeMux I__8008 (
            .O(N__34897),
            .I(N__34843));
    LocalMux I__8007 (
            .O(N__34894),
            .I(N__34839));
    InMux I__8006 (
            .O(N__34891),
            .I(N__34836));
    InMux I__8005 (
            .O(N__34888),
            .I(N__34831));
    InMux I__8004 (
            .O(N__34885),
            .I(N__34831));
    InMux I__8003 (
            .O(N__34882),
            .I(N__34826));
    InMux I__8002 (
            .O(N__34881),
            .I(N__34826));
    InMux I__8001 (
            .O(N__34880),
            .I(N__34823));
    InMux I__8000 (
            .O(N__34879),
            .I(N__34820));
    InMux I__7999 (
            .O(N__34876),
            .I(N__34817));
    Span4Mux_h I__7998 (
            .O(N__34873),
            .I(N__34814));
    InMux I__7997 (
            .O(N__34870),
            .I(N__34811));
    Span4Mux_v I__7996 (
            .O(N__34865),
            .I(N__34804));
    Span4Mux_h I__7995 (
            .O(N__34858),
            .I(N__34804));
    Span4Mux_v I__7994 (
            .O(N__34855),
            .I(N__34804));
    Span4Mux_h I__7993 (
            .O(N__34846),
            .I(N__34801));
    InMux I__7992 (
            .O(N__34843),
            .I(N__34796));
    InMux I__7991 (
            .O(N__34842),
            .I(N__34796));
    Span12Mux_v I__7990 (
            .O(N__34839),
            .I(N__34787));
    LocalMux I__7989 (
            .O(N__34836),
            .I(N__34787));
    LocalMux I__7988 (
            .O(N__34831),
            .I(N__34787));
    LocalMux I__7987 (
            .O(N__34826),
            .I(N__34787));
    LocalMux I__7986 (
            .O(N__34823),
            .I(this_vga_signals_M_vcounter_q_5));
    LocalMux I__7985 (
            .O(N__34820),
            .I(this_vga_signals_M_vcounter_q_5));
    LocalMux I__7984 (
            .O(N__34817),
            .I(this_vga_signals_M_vcounter_q_5));
    Odrv4 I__7983 (
            .O(N__34814),
            .I(this_vga_signals_M_vcounter_q_5));
    LocalMux I__7982 (
            .O(N__34811),
            .I(this_vga_signals_M_vcounter_q_5));
    Odrv4 I__7981 (
            .O(N__34804),
            .I(this_vga_signals_M_vcounter_q_5));
    Odrv4 I__7980 (
            .O(N__34801),
            .I(this_vga_signals_M_vcounter_q_5));
    LocalMux I__7979 (
            .O(N__34796),
            .I(this_vga_signals_M_vcounter_q_5));
    Odrv12 I__7978 (
            .O(N__34787),
            .I(this_vga_signals_M_vcounter_q_5));
    CascadeMux I__7977 (
            .O(N__34768),
            .I(N__34765));
    InMux I__7976 (
            .O(N__34765),
            .I(N__34762));
    LocalMux I__7975 (
            .O(N__34762),
            .I(N__34759));
    Span4Mux_v I__7974 (
            .O(N__34759),
            .I(N__34755));
    InMux I__7973 (
            .O(N__34758),
            .I(N__34752));
    Span4Mux_h I__7972 (
            .O(N__34755),
            .I(N__34739));
    LocalMux I__7971 (
            .O(N__34752),
            .I(N__34739));
    InMux I__7970 (
            .O(N__34751),
            .I(N__34736));
    InMux I__7969 (
            .O(N__34750),
            .I(N__34732));
    InMux I__7968 (
            .O(N__34749),
            .I(N__34729));
    InMux I__7967 (
            .O(N__34748),
            .I(N__34726));
    InMux I__7966 (
            .O(N__34747),
            .I(N__34723));
    InMux I__7965 (
            .O(N__34746),
            .I(N__34720));
    InMux I__7964 (
            .O(N__34745),
            .I(N__34717));
    InMux I__7963 (
            .O(N__34744),
            .I(N__34713));
    Span4Mux_v I__7962 (
            .O(N__34739),
            .I(N__34710));
    LocalMux I__7961 (
            .O(N__34736),
            .I(N__34707));
    InMux I__7960 (
            .O(N__34735),
            .I(N__34700));
    LocalMux I__7959 (
            .O(N__34732),
            .I(N__34697));
    LocalMux I__7958 (
            .O(N__34729),
            .I(N__34692));
    LocalMux I__7957 (
            .O(N__34726),
            .I(N__34692));
    LocalMux I__7956 (
            .O(N__34723),
            .I(N__34685));
    LocalMux I__7955 (
            .O(N__34720),
            .I(N__34685));
    LocalMux I__7954 (
            .O(N__34717),
            .I(N__34685));
    InMux I__7953 (
            .O(N__34716),
            .I(N__34682));
    LocalMux I__7952 (
            .O(N__34713),
            .I(N__34679));
    Span4Mux_h I__7951 (
            .O(N__34710),
            .I(N__34676));
    Span12Mux_h I__7950 (
            .O(N__34707),
            .I(N__34673));
    InMux I__7949 (
            .O(N__34706),
            .I(N__34670));
    InMux I__7948 (
            .O(N__34705),
            .I(N__34667));
    InMux I__7947 (
            .O(N__34704),
            .I(N__34662));
    InMux I__7946 (
            .O(N__34703),
            .I(N__34662));
    LocalMux I__7945 (
            .O(N__34700),
            .I(N__34651));
    Span4Mux_h I__7944 (
            .O(N__34697),
            .I(N__34651));
    Span4Mux_h I__7943 (
            .O(N__34692),
            .I(N__34651));
    Span4Mux_v I__7942 (
            .O(N__34685),
            .I(N__34651));
    LocalMux I__7941 (
            .O(N__34682),
            .I(N__34651));
    Span4Mux_v I__7940 (
            .O(N__34679),
            .I(N__34648));
    Odrv4 I__7939 (
            .O(N__34676),
            .I(this_vga_signals_M_vcounter_q_6));
    Odrv12 I__7938 (
            .O(N__34673),
            .I(this_vga_signals_M_vcounter_q_6));
    LocalMux I__7937 (
            .O(N__34670),
            .I(this_vga_signals_M_vcounter_q_6));
    LocalMux I__7936 (
            .O(N__34667),
            .I(this_vga_signals_M_vcounter_q_6));
    LocalMux I__7935 (
            .O(N__34662),
            .I(this_vga_signals_M_vcounter_q_6));
    Odrv4 I__7934 (
            .O(N__34651),
            .I(this_vga_signals_M_vcounter_q_6));
    Odrv4 I__7933 (
            .O(N__34648),
            .I(this_vga_signals_M_vcounter_q_6));
    CascadeMux I__7932 (
            .O(N__34633),
            .I(N__34630));
    InMux I__7931 (
            .O(N__34630),
            .I(N__34627));
    LocalMux I__7930 (
            .O(N__34627),
            .I(\this_vga_signals.vaddress_0_0_7 ));
    CascadeMux I__7929 (
            .O(N__34624),
            .I(N__34621));
    InMux I__7928 (
            .O(N__34621),
            .I(N__34618));
    LocalMux I__7927 (
            .O(N__34618),
            .I(N__34615));
    Span4Mux_h I__7926 (
            .O(N__34615),
            .I(N__34611));
    CascadeMux I__7925 (
            .O(N__34614),
            .I(N__34608));
    Span4Mux_h I__7924 (
            .O(N__34611),
            .I(N__34605));
    InMux I__7923 (
            .O(N__34608),
            .I(N__34602));
    Odrv4 I__7922 (
            .O(N__34605),
            .I(M_this_scroll_qZ0Z_6));
    LocalMux I__7921 (
            .O(N__34602),
            .I(M_this_scroll_qZ0Z_6));
    InMux I__7920 (
            .O(N__34597),
            .I(N__34594));
    LocalMux I__7919 (
            .O(N__34594),
            .I(N__34591));
    Span4Mux_h I__7918 (
            .O(N__34591),
            .I(N__34588));
    Span4Mux_h I__7917 (
            .O(N__34588),
            .I(N__34585));
    Odrv4 I__7916 (
            .O(N__34585),
            .I(\this_ppu.M_screen_y_q_esr_RNILD7F7Z0Z_6 ));
    InMux I__7915 (
            .O(N__34582),
            .I(N__34579));
    LocalMux I__7914 (
            .O(N__34579),
            .I(N__34573));
    InMux I__7913 (
            .O(N__34578),
            .I(N__34570));
    InMux I__7912 (
            .O(N__34577),
            .I(N__34567));
    InMux I__7911 (
            .O(N__34576),
            .I(N__34562));
    Span4Mux_s3_v I__7910 (
            .O(N__34573),
            .I(N__34557));
    LocalMux I__7909 (
            .O(N__34570),
            .I(N__34557));
    LocalMux I__7908 (
            .O(N__34567),
            .I(N__34554));
    InMux I__7907 (
            .O(N__34566),
            .I(N__34550));
    InMux I__7906 (
            .O(N__34565),
            .I(N__34547));
    LocalMux I__7905 (
            .O(N__34562),
            .I(N__34544));
    Span4Mux_v I__7904 (
            .O(N__34557),
            .I(N__34541));
    Span4Mux_h I__7903 (
            .O(N__34554),
            .I(N__34538));
    InMux I__7902 (
            .O(N__34553),
            .I(N__34535));
    LocalMux I__7901 (
            .O(N__34550),
            .I(N__34532));
    LocalMux I__7900 (
            .O(N__34547),
            .I(N__34529));
    Span12Mux_s10_h I__7899 (
            .O(N__34544),
            .I(N__34525));
    Sp12to4 I__7898 (
            .O(N__34541),
            .I(N__34522));
    Sp12to4 I__7897 (
            .O(N__34538),
            .I(N__34519));
    LocalMux I__7896 (
            .O(N__34535),
            .I(N__34516));
    Span4Mux_v I__7895 (
            .O(N__34532),
            .I(N__34511));
    Span4Mux_h I__7894 (
            .O(N__34529),
            .I(N__34511));
    InMux I__7893 (
            .O(N__34528),
            .I(N__34508));
    Span12Mux_v I__7892 (
            .O(N__34525),
            .I(N__34505));
    Span12Mux_h I__7891 (
            .O(N__34522),
            .I(N__34498));
    Span12Mux_v I__7890 (
            .O(N__34519),
            .I(N__34498));
    Span12Mux_s10_h I__7889 (
            .O(N__34516),
            .I(N__34498));
    Span4Mux_v I__7888 (
            .O(N__34511),
            .I(N__34493));
    LocalMux I__7887 (
            .O(N__34508),
            .I(N__34493));
    Odrv12 I__7886 (
            .O(N__34505),
            .I(M_this_spr_ram_write_data_3));
    Odrv12 I__7885 (
            .O(N__34498),
            .I(M_this_spr_ram_write_data_3));
    Odrv4 I__7884 (
            .O(N__34493),
            .I(M_this_spr_ram_write_data_3));
    InMux I__7883 (
            .O(N__34486),
            .I(N__34483));
    LocalMux I__7882 (
            .O(N__34483),
            .I(N__34480));
    Odrv4 I__7881 (
            .O(N__34480),
            .I(\this_ppu.M_this_state_q_srsts_0_0_a2_1_xZ0Z_0 ));
    InMux I__7880 (
            .O(N__34477),
            .I(N__34473));
    InMux I__7879 (
            .O(N__34476),
            .I(N__34470));
    LocalMux I__7878 (
            .O(N__34473),
            .I(N__34464));
    LocalMux I__7877 (
            .O(N__34470),
            .I(N__34464));
    InMux I__7876 (
            .O(N__34469),
            .I(N__34461));
    Span4Mux_v I__7875 (
            .O(N__34464),
            .I(N__34458));
    LocalMux I__7874 (
            .O(N__34461),
            .I(N__34455));
    Span4Mux_h I__7873 (
            .O(N__34458),
            .I(N__34451));
    Span12Mux_h I__7872 (
            .O(N__34455),
            .I(N__34448));
    InMux I__7871 (
            .O(N__34454),
            .I(N__34445));
    Odrv4 I__7870 (
            .O(N__34451),
            .I(\this_ppu.N_798_0 ));
    Odrv12 I__7869 (
            .O(N__34448),
            .I(\this_ppu.N_798_0 ));
    LocalMux I__7868 (
            .O(N__34445),
            .I(\this_ppu.N_798_0 ));
    InMux I__7867 (
            .O(N__34438),
            .I(N__34434));
    InMux I__7866 (
            .O(N__34437),
            .I(N__34431));
    LocalMux I__7865 (
            .O(N__34434),
            .I(N__34427));
    LocalMux I__7864 (
            .O(N__34431),
            .I(N__34424));
    InMux I__7863 (
            .O(N__34430),
            .I(N__34421));
    Span4Mux_v I__7862 (
            .O(N__34427),
            .I(N__34418));
    Span4Mux_v I__7861 (
            .O(N__34424),
            .I(N__34413));
    LocalMux I__7860 (
            .O(N__34421),
            .I(N__34413));
    Span4Mux_h I__7859 (
            .O(N__34418),
            .I(N__34408));
    Span4Mux_h I__7858 (
            .O(N__34413),
            .I(N__34408));
    Odrv4 I__7857 (
            .O(N__34408),
            .I(\this_ppu.N_1426 ));
    InMux I__7856 (
            .O(N__34405),
            .I(N__34402));
    LocalMux I__7855 (
            .O(N__34402),
            .I(N__34399));
    Span4Mux_h I__7854 (
            .O(N__34399),
            .I(N__34396));
    Span4Mux_h I__7853 (
            .O(N__34396),
            .I(N__34393));
    Span4Mux_h I__7852 (
            .O(N__34393),
            .I(N__34390));
    Span4Mux_h I__7851 (
            .O(N__34390),
            .I(N__34387));
    Odrv4 I__7850 (
            .O(N__34387),
            .I(M_this_ppu_vram_data_3));
    InMux I__7849 (
            .O(N__34384),
            .I(N__34381));
    LocalMux I__7848 (
            .O(N__34381),
            .I(M_this_spr_ram_read_data_2));
    CascadeMux I__7847 (
            .O(N__34378),
            .I(M_this_spr_ram_read_data_1_cascade_));
    InMux I__7846 (
            .O(N__34375),
            .I(N__34371));
    InMux I__7845 (
            .O(N__34374),
            .I(N__34365));
    LocalMux I__7844 (
            .O(N__34371),
            .I(N__34362));
    InMux I__7843 (
            .O(N__34370),
            .I(N__34357));
    InMux I__7842 (
            .O(N__34369),
            .I(N__34357));
    InMux I__7841 (
            .O(N__34368),
            .I(N__34354));
    LocalMux I__7840 (
            .O(N__34365),
            .I(N__34351));
    Span12Mux_h I__7839 (
            .O(N__34362),
            .I(N__34348));
    LocalMux I__7838 (
            .O(N__34357),
            .I(N__34341));
    LocalMux I__7837 (
            .O(N__34354),
            .I(N__34341));
    Span12Mux_v I__7836 (
            .O(N__34351),
            .I(N__34341));
    Odrv12 I__7835 (
            .O(N__34348),
            .I(\this_ppu.N_1000_0 ));
    Odrv12 I__7834 (
            .O(N__34341),
            .I(\this_ppu.N_1000_0 ));
    InMux I__7833 (
            .O(N__34336),
            .I(N__34333));
    LocalMux I__7832 (
            .O(N__34333),
            .I(M_this_spr_ram_read_data_1));
    InMux I__7831 (
            .O(N__34330),
            .I(N__34327));
    LocalMux I__7830 (
            .O(N__34327),
            .I(N__34324));
    Span4Mux_v I__7829 (
            .O(N__34324),
            .I(N__34321));
    Span4Mux_h I__7828 (
            .O(N__34321),
            .I(N__34318));
    Sp12to4 I__7827 (
            .O(N__34318),
            .I(N__34315));
    Odrv12 I__7826 (
            .O(N__34315),
            .I(M_this_ppu_vram_data_1));
    InMux I__7825 (
            .O(N__34312),
            .I(N__34309));
    LocalMux I__7824 (
            .O(N__34309),
            .I(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0 ));
    InMux I__7823 (
            .O(N__34306),
            .I(N__34303));
    LocalMux I__7822 (
            .O(N__34303),
            .I(N__34300));
    Span4Mux_h I__7821 (
            .O(N__34300),
            .I(N__34297));
    Span4Mux_h I__7820 (
            .O(N__34297),
            .I(N__34293));
    InMux I__7819 (
            .O(N__34296),
            .I(N__34290));
    Odrv4 I__7818 (
            .O(N__34293),
            .I(M_this_spr_ram_read_data_0));
    LocalMux I__7817 (
            .O(N__34290),
            .I(M_this_spr_ram_read_data_0));
    InMux I__7816 (
            .O(N__34285),
            .I(N__34281));
    InMux I__7815 (
            .O(N__34284),
            .I(N__34278));
    LocalMux I__7814 (
            .O(N__34281),
            .I(N__34274));
    LocalMux I__7813 (
            .O(N__34278),
            .I(N__34271));
    InMux I__7812 (
            .O(N__34277),
            .I(N__34268));
    Span4Mux_h I__7811 (
            .O(N__34274),
            .I(N__34265));
    Span4Mux_v I__7810 (
            .O(N__34271),
            .I(N__34262));
    LocalMux I__7809 (
            .O(N__34268),
            .I(N__34259));
    Odrv4 I__7808 (
            .O(N__34265),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    Odrv4 I__7807 (
            .O(N__34262),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    Odrv4 I__7806 (
            .O(N__34259),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    CEMux I__7805 (
            .O(N__34252),
            .I(N__34231));
    CEMux I__7804 (
            .O(N__34251),
            .I(N__34231));
    CEMux I__7803 (
            .O(N__34250),
            .I(N__34231));
    CEMux I__7802 (
            .O(N__34249),
            .I(N__34231));
    CEMux I__7801 (
            .O(N__34248),
            .I(N__34231));
    CEMux I__7800 (
            .O(N__34247),
            .I(N__34231));
    CEMux I__7799 (
            .O(N__34246),
            .I(N__34231));
    GlobalMux I__7798 (
            .O(N__34231),
            .I(N__34228));
    gio2CtrlBuf I__7797 (
            .O(N__34228),
            .I(\this_vga_signals.N_1307_0_g ));
    InMux I__7796 (
            .O(N__34225),
            .I(N__34222));
    LocalMux I__7795 (
            .O(N__34222),
            .I(N__34211));
    SRMux I__7794 (
            .O(N__34221),
            .I(N__34192));
    SRMux I__7793 (
            .O(N__34220),
            .I(N__34192));
    SRMux I__7792 (
            .O(N__34219),
            .I(N__34192));
    SRMux I__7791 (
            .O(N__34218),
            .I(N__34192));
    SRMux I__7790 (
            .O(N__34217),
            .I(N__34192));
    SRMux I__7789 (
            .O(N__34216),
            .I(N__34192));
    SRMux I__7788 (
            .O(N__34215),
            .I(N__34192));
    SRMux I__7787 (
            .O(N__34214),
            .I(N__34192));
    Glb2LocalMux I__7786 (
            .O(N__34211),
            .I(N__34192));
    GlobalMux I__7785 (
            .O(N__34192),
            .I(N__34189));
    gio2CtrlBuf I__7784 (
            .O(N__34189),
            .I(\this_vga_signals.N_1637_g ));
    InMux I__7783 (
            .O(N__34186),
            .I(N__34183));
    LocalMux I__7782 (
            .O(N__34183),
            .I(N__34180));
    Odrv4 I__7781 (
            .O(N__34180),
            .I(\this_vga_signals.N_5_i_0 ));
    CascadeMux I__7780 (
            .O(N__34177),
            .I(\this_vga_signals.N_5_i_0_cascade_ ));
    InMux I__7779 (
            .O(N__34174),
            .I(N__34171));
    LocalMux I__7778 (
            .O(N__34171),
            .I(N__34168));
    Span4Mux_v I__7777 (
            .O(N__34168),
            .I(N__34165));
    Odrv4 I__7776 (
            .O(N__34165),
            .I(\this_vga_signals.mult1_un47_sum_0_1 ));
    InMux I__7775 (
            .O(N__34162),
            .I(N__34159));
    LocalMux I__7774 (
            .O(N__34159),
            .I(N__34156));
    Odrv12 I__7773 (
            .O(N__34156),
            .I(\this_vga_signals.g0_21_1 ));
    InMux I__7772 (
            .O(N__34153),
            .I(N__34149));
    InMux I__7771 (
            .O(N__34152),
            .I(N__34146));
    LocalMux I__7770 (
            .O(N__34149),
            .I(\this_vga_signals.mult1_un47_sum_axb1 ));
    LocalMux I__7769 (
            .O(N__34146),
            .I(\this_vga_signals.mult1_un47_sum_axb1 ));
    InMux I__7768 (
            .O(N__34141),
            .I(N__34138));
    LocalMux I__7767 (
            .O(N__34138),
            .I(N__34133));
    CascadeMux I__7766 (
            .O(N__34137),
            .I(N__34127));
    CascadeMux I__7765 (
            .O(N__34136),
            .I(N__34120));
    Span4Mux_h I__7764 (
            .O(N__34133),
            .I(N__34115));
    InMux I__7763 (
            .O(N__34132),
            .I(N__34110));
    InMux I__7762 (
            .O(N__34131),
            .I(N__34110));
    InMux I__7761 (
            .O(N__34130),
            .I(N__34101));
    InMux I__7760 (
            .O(N__34127),
            .I(N__34101));
    InMux I__7759 (
            .O(N__34126),
            .I(N__34101));
    InMux I__7758 (
            .O(N__34125),
            .I(N__34101));
    InMux I__7757 (
            .O(N__34124),
            .I(N__34098));
    InMux I__7756 (
            .O(N__34123),
            .I(N__34095));
    InMux I__7755 (
            .O(N__34120),
            .I(N__34088));
    InMux I__7754 (
            .O(N__34119),
            .I(N__34088));
    InMux I__7753 (
            .O(N__34118),
            .I(N__34088));
    Odrv4 I__7752 (
            .O(N__34115),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    LocalMux I__7751 (
            .O(N__34110),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    LocalMux I__7750 (
            .O(N__34101),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    LocalMux I__7749 (
            .O(N__34098),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    LocalMux I__7748 (
            .O(N__34095),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    LocalMux I__7747 (
            .O(N__34088),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    InMux I__7746 (
            .O(N__34075),
            .I(N__34061));
    InMux I__7745 (
            .O(N__34074),
            .I(N__34061));
    InMux I__7744 (
            .O(N__34073),
            .I(N__34061));
    InMux I__7743 (
            .O(N__34072),
            .I(N__34058));
    InMux I__7742 (
            .O(N__34071),
            .I(N__34053));
    InMux I__7741 (
            .O(N__34070),
            .I(N__34053));
    InMux I__7740 (
            .O(N__34069),
            .I(N__34048));
    InMux I__7739 (
            .O(N__34068),
            .I(N__34048));
    LocalMux I__7738 (
            .O(N__34061),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_3 ));
    LocalMux I__7737 (
            .O(N__34058),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_3 ));
    LocalMux I__7736 (
            .O(N__34053),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_3 ));
    LocalMux I__7735 (
            .O(N__34048),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_3 ));
    InMux I__7734 (
            .O(N__34039),
            .I(N__34036));
    LocalMux I__7733 (
            .O(N__34036),
            .I(N__34033));
    Span4Mux_h I__7732 (
            .O(N__34033),
            .I(N__34030));
    Odrv4 I__7731 (
            .O(N__34030),
            .I(\this_vga_signals.mult1_un47_sum_1_1 ));
    InMux I__7730 (
            .O(N__34027),
            .I(N__34024));
    LocalMux I__7729 (
            .O(N__34024),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_6 ));
    InMux I__7728 (
            .O(N__34021),
            .I(N__34018));
    LocalMux I__7727 (
            .O(N__34018),
            .I(N__34015));
    Span4Mux_h I__7726 (
            .O(N__34015),
            .I(N__34012));
    Span4Mux_v I__7725 (
            .O(N__34012),
            .I(N__34009));
    Odrv4 I__7724 (
            .O(N__34009),
            .I(\this_spr_ram.mem_out_bus4_2 ));
    InMux I__7723 (
            .O(N__34006),
            .I(N__34003));
    LocalMux I__7722 (
            .O(N__34003),
            .I(N__34000));
    Span4Mux_h I__7721 (
            .O(N__34000),
            .I(N__33997));
    Span4Mux_v I__7720 (
            .O(N__33997),
            .I(N__33994));
    Span4Mux_v I__7719 (
            .O(N__33994),
            .I(N__33991));
    Odrv4 I__7718 (
            .O(N__33991),
            .I(\this_spr_ram.mem_out_bus0_2 ));
    CascadeMux I__7717 (
            .O(N__33988),
            .I(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0_cascade_ ));
    CascadeMux I__7716 (
            .O(N__33985),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ));
    CascadeMux I__7715 (
            .O(N__33982),
            .I(M_this_spr_ram_read_data_2_cascade_));
    InMux I__7714 (
            .O(N__33979),
            .I(N__33976));
    LocalMux I__7713 (
            .O(N__33976),
            .I(N__33973));
    Span12Mux_s9_h I__7712 (
            .O(N__33973),
            .I(N__33970));
    Span12Mux_h I__7711 (
            .O(N__33970),
            .I(N__33967));
    Odrv12 I__7710 (
            .O(N__33967),
            .I(M_this_ppu_vram_data_2));
    InMux I__7709 (
            .O(N__33964),
            .I(N__33961));
    LocalMux I__7708 (
            .O(N__33961),
            .I(N__33958));
    Span4Mux_v I__7707 (
            .O(N__33958),
            .I(N__33955));
    Span4Mux_h I__7706 (
            .O(N__33955),
            .I(N__33952));
    Odrv4 I__7705 (
            .O(N__33952),
            .I(\this_spr_ram.mem_out_bus5_0 ));
    InMux I__7704 (
            .O(N__33949),
            .I(N__33946));
    LocalMux I__7703 (
            .O(N__33946),
            .I(N__33943));
    Span4Mux_v I__7702 (
            .O(N__33943),
            .I(N__33940));
    Span4Mux_h I__7701 (
            .O(N__33940),
            .I(N__33937));
    Span4Mux_v I__7700 (
            .O(N__33937),
            .I(N__33934));
    Odrv4 I__7699 (
            .O(N__33934),
            .I(\this_spr_ram.mem_out_bus1_0 ));
    InMux I__7698 (
            .O(N__33931),
            .I(N__33928));
    LocalMux I__7697 (
            .O(N__33928),
            .I(N__33925));
    Span4Mux_h I__7696 (
            .O(N__33925),
            .I(N__33922));
    Odrv4 I__7695 (
            .O(N__33922),
            .I(\this_spr_ram.mem_out_bus4_1 ));
    InMux I__7694 (
            .O(N__33919),
            .I(N__33916));
    LocalMux I__7693 (
            .O(N__33916),
            .I(N__33913));
    Span4Mux_h I__7692 (
            .O(N__33913),
            .I(N__33910));
    Span4Mux_v I__7691 (
            .O(N__33910),
            .I(N__33907));
    Span4Mux_v I__7690 (
            .O(N__33907),
            .I(N__33904));
    Span4Mux_v I__7689 (
            .O(N__33904),
            .I(N__33901));
    Odrv4 I__7688 (
            .O(N__33901),
            .I(\this_spr_ram.mem_out_bus0_1 ));
    CascadeMux I__7687 (
            .O(N__33898),
            .I(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0_cascade_ ));
    CascadeMux I__7686 (
            .O(N__33895),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ));
    CascadeMux I__7685 (
            .O(N__33892),
            .I(N__33887));
    CascadeMux I__7684 (
            .O(N__33891),
            .I(N__33882));
    CascadeMux I__7683 (
            .O(N__33890),
            .I(N__33877));
    InMux I__7682 (
            .O(N__33887),
            .I(N__33873));
    CascadeMux I__7681 (
            .O(N__33886),
            .I(N__33870));
    CascadeMux I__7680 (
            .O(N__33885),
            .I(N__33867));
    InMux I__7679 (
            .O(N__33882),
            .I(N__33864));
    CascadeMux I__7678 (
            .O(N__33881),
            .I(N__33861));
    CascadeMux I__7677 (
            .O(N__33880),
            .I(N__33857));
    InMux I__7676 (
            .O(N__33877),
            .I(N__33853));
    CascadeMux I__7675 (
            .O(N__33876),
            .I(N__33850));
    LocalMux I__7674 (
            .O(N__33873),
            .I(N__33846));
    InMux I__7673 (
            .O(N__33870),
            .I(N__33843));
    InMux I__7672 (
            .O(N__33867),
            .I(N__33840));
    LocalMux I__7671 (
            .O(N__33864),
            .I(N__33837));
    InMux I__7670 (
            .O(N__33861),
            .I(N__33834));
    CascadeMux I__7669 (
            .O(N__33860),
            .I(N__33831));
    InMux I__7668 (
            .O(N__33857),
            .I(N__33827));
    CascadeMux I__7667 (
            .O(N__33856),
            .I(N__33824));
    LocalMux I__7666 (
            .O(N__33853),
            .I(N__33821));
    InMux I__7665 (
            .O(N__33850),
            .I(N__33818));
    CascadeMux I__7664 (
            .O(N__33849),
            .I(N__33815));
    Span4Mux_s1_v I__7663 (
            .O(N__33846),
            .I(N__33806));
    LocalMux I__7662 (
            .O(N__33843),
            .I(N__33806));
    LocalMux I__7661 (
            .O(N__33840),
            .I(N__33806));
    Span4Mux_h I__7660 (
            .O(N__33837),
            .I(N__33801));
    LocalMux I__7659 (
            .O(N__33834),
            .I(N__33801));
    InMux I__7658 (
            .O(N__33831),
            .I(N__33798));
    CascadeMux I__7657 (
            .O(N__33830),
            .I(N__33795));
    LocalMux I__7656 (
            .O(N__33827),
            .I(N__33791));
    InMux I__7655 (
            .O(N__33824),
            .I(N__33788));
    Span4Mux_v I__7654 (
            .O(N__33821),
            .I(N__33783));
    LocalMux I__7653 (
            .O(N__33818),
            .I(N__33783));
    InMux I__7652 (
            .O(N__33815),
            .I(N__33780));
    CascadeMux I__7651 (
            .O(N__33814),
            .I(N__33777));
    CascadeMux I__7650 (
            .O(N__33813),
            .I(N__33774));
    Span4Mux_v I__7649 (
            .O(N__33806),
            .I(N__33770));
    Span4Mux_v I__7648 (
            .O(N__33801),
            .I(N__33765));
    LocalMux I__7647 (
            .O(N__33798),
            .I(N__33765));
    InMux I__7646 (
            .O(N__33795),
            .I(N__33762));
    CascadeMux I__7645 (
            .O(N__33794),
            .I(N__33759));
    Span4Mux_v I__7644 (
            .O(N__33791),
            .I(N__33754));
    LocalMux I__7643 (
            .O(N__33788),
            .I(N__33754));
    Span4Mux_v I__7642 (
            .O(N__33783),
            .I(N__33749));
    LocalMux I__7641 (
            .O(N__33780),
            .I(N__33749));
    InMux I__7640 (
            .O(N__33777),
            .I(N__33746));
    InMux I__7639 (
            .O(N__33774),
            .I(N__33743));
    CascadeMux I__7638 (
            .O(N__33773),
            .I(N__33740));
    Sp12to4 I__7637 (
            .O(N__33770),
            .I(N__33737));
    Span4Mux_h I__7636 (
            .O(N__33765),
            .I(N__33732));
    LocalMux I__7635 (
            .O(N__33762),
            .I(N__33732));
    InMux I__7634 (
            .O(N__33759),
            .I(N__33729));
    Span4Mux_v I__7633 (
            .O(N__33754),
            .I(N__33722));
    Span4Mux_h I__7632 (
            .O(N__33749),
            .I(N__33722));
    LocalMux I__7631 (
            .O(N__33746),
            .I(N__33722));
    LocalMux I__7630 (
            .O(N__33743),
            .I(N__33719));
    InMux I__7629 (
            .O(N__33740),
            .I(N__33716));
    Span12Mux_h I__7628 (
            .O(N__33737),
            .I(N__33713));
    Span4Mux_v I__7627 (
            .O(N__33732),
            .I(N__33708));
    LocalMux I__7626 (
            .O(N__33729),
            .I(N__33708));
    Span4Mux_v I__7625 (
            .O(N__33722),
            .I(N__33701));
    Span4Mux_v I__7624 (
            .O(N__33719),
            .I(N__33701));
    LocalMux I__7623 (
            .O(N__33716),
            .I(N__33701));
    Span12Mux_v I__7622 (
            .O(N__33713),
            .I(N__33697));
    Span4Mux_h I__7621 (
            .O(N__33708),
            .I(N__33692));
    Span4Mux_h I__7620 (
            .O(N__33701),
            .I(N__33692));
    InMux I__7619 (
            .O(N__33700),
            .I(N__33689));
    Odrv12 I__7618 (
            .O(N__33697),
            .I(M_this_spr_address_qZ0Z_8));
    Odrv4 I__7617 (
            .O(N__33692),
            .I(M_this_spr_address_qZ0Z_8));
    LocalMux I__7616 (
            .O(N__33689),
            .I(M_this_spr_address_qZ0Z_8));
    InMux I__7615 (
            .O(N__33682),
            .I(bfn_22_15_0_));
    CascadeMux I__7614 (
            .O(N__33679),
            .I(N__33675));
    CascadeMux I__7613 (
            .O(N__33678),
            .I(N__33670));
    InMux I__7612 (
            .O(N__33675),
            .I(N__33666));
    CascadeMux I__7611 (
            .O(N__33674),
            .I(N__33663));
    CascadeMux I__7610 (
            .O(N__33673),
            .I(N__33659));
    InMux I__7609 (
            .O(N__33670),
            .I(N__33655));
    CascadeMux I__7608 (
            .O(N__33669),
            .I(N__33652));
    LocalMux I__7607 (
            .O(N__33666),
            .I(N__33646));
    InMux I__7606 (
            .O(N__33663),
            .I(N__33643));
    CascadeMux I__7605 (
            .O(N__33662),
            .I(N__33640));
    InMux I__7604 (
            .O(N__33659),
            .I(N__33637));
    CascadeMux I__7603 (
            .O(N__33658),
            .I(N__33634));
    LocalMux I__7602 (
            .O(N__33655),
            .I(N__33630));
    InMux I__7601 (
            .O(N__33652),
            .I(N__33627));
    CascadeMux I__7600 (
            .O(N__33651),
            .I(N__33624));
    CascadeMux I__7599 (
            .O(N__33650),
            .I(N__33621));
    CascadeMux I__7598 (
            .O(N__33649),
            .I(N__33617));
    Span4Mux_s1_v I__7597 (
            .O(N__33646),
            .I(N__33611));
    LocalMux I__7596 (
            .O(N__33643),
            .I(N__33611));
    InMux I__7595 (
            .O(N__33640),
            .I(N__33608));
    LocalMux I__7594 (
            .O(N__33637),
            .I(N__33604));
    InMux I__7593 (
            .O(N__33634),
            .I(N__33601));
    CascadeMux I__7592 (
            .O(N__33633),
            .I(N__33598));
    Span4Mux_h I__7591 (
            .O(N__33630),
            .I(N__33592));
    LocalMux I__7590 (
            .O(N__33627),
            .I(N__33592));
    InMux I__7589 (
            .O(N__33624),
            .I(N__33589));
    InMux I__7588 (
            .O(N__33621),
            .I(N__33586));
    CascadeMux I__7587 (
            .O(N__33620),
            .I(N__33583));
    InMux I__7586 (
            .O(N__33617),
            .I(N__33580));
    CascadeMux I__7585 (
            .O(N__33616),
            .I(N__33577));
    Span4Mux_v I__7584 (
            .O(N__33611),
            .I(N__33573));
    LocalMux I__7583 (
            .O(N__33608),
            .I(N__33570));
    CascadeMux I__7582 (
            .O(N__33607),
            .I(N__33567));
    Span4Mux_v I__7581 (
            .O(N__33604),
            .I(N__33562));
    LocalMux I__7580 (
            .O(N__33601),
            .I(N__33562));
    InMux I__7579 (
            .O(N__33598),
            .I(N__33559));
    CascadeMux I__7578 (
            .O(N__33597),
            .I(N__33556));
    Span4Mux_v I__7577 (
            .O(N__33592),
            .I(N__33549));
    LocalMux I__7576 (
            .O(N__33589),
            .I(N__33549));
    LocalMux I__7575 (
            .O(N__33586),
            .I(N__33549));
    InMux I__7574 (
            .O(N__33583),
            .I(N__33546));
    LocalMux I__7573 (
            .O(N__33580),
            .I(N__33543));
    InMux I__7572 (
            .O(N__33577),
            .I(N__33540));
    CascadeMux I__7571 (
            .O(N__33576),
            .I(N__33537));
    Sp12to4 I__7570 (
            .O(N__33573),
            .I(N__33534));
    Span12Mux_s9_h I__7569 (
            .O(N__33570),
            .I(N__33531));
    InMux I__7568 (
            .O(N__33567),
            .I(N__33528));
    Span4Mux_h I__7567 (
            .O(N__33562),
            .I(N__33523));
    LocalMux I__7566 (
            .O(N__33559),
            .I(N__33523));
    InMux I__7565 (
            .O(N__33556),
            .I(N__33520));
    Span4Mux_v I__7564 (
            .O(N__33549),
            .I(N__33517));
    LocalMux I__7563 (
            .O(N__33546),
            .I(N__33514));
    Span4Mux_v I__7562 (
            .O(N__33543),
            .I(N__33509));
    LocalMux I__7561 (
            .O(N__33540),
            .I(N__33509));
    InMux I__7560 (
            .O(N__33537),
            .I(N__33506));
    Span12Mux_h I__7559 (
            .O(N__33534),
            .I(N__33503));
    Span12Mux_h I__7558 (
            .O(N__33531),
            .I(N__33500));
    LocalMux I__7557 (
            .O(N__33528),
            .I(N__33497));
    Span4Mux_v I__7556 (
            .O(N__33523),
            .I(N__33492));
    LocalMux I__7555 (
            .O(N__33520),
            .I(N__33492));
    Span4Mux_v I__7554 (
            .O(N__33517),
            .I(N__33483));
    Span4Mux_v I__7553 (
            .O(N__33514),
            .I(N__33483));
    Span4Mux_v I__7552 (
            .O(N__33509),
            .I(N__33483));
    LocalMux I__7551 (
            .O(N__33506),
            .I(N__33483));
    Span12Mux_v I__7550 (
            .O(N__33503),
            .I(N__33479));
    Span12Mux_v I__7549 (
            .O(N__33500),
            .I(N__33474));
    Span12Mux_s10_h I__7548 (
            .O(N__33497),
            .I(N__33474));
    Span4Mux_h I__7547 (
            .O(N__33492),
            .I(N__33469));
    Span4Mux_h I__7546 (
            .O(N__33483),
            .I(N__33469));
    InMux I__7545 (
            .O(N__33482),
            .I(N__33466));
    Odrv12 I__7544 (
            .O(N__33479),
            .I(M_this_spr_address_qZ0Z_9));
    Odrv12 I__7543 (
            .O(N__33474),
            .I(M_this_spr_address_qZ0Z_9));
    Odrv4 I__7542 (
            .O(N__33469),
            .I(M_this_spr_address_qZ0Z_9));
    LocalMux I__7541 (
            .O(N__33466),
            .I(M_this_spr_address_qZ0Z_9));
    InMux I__7540 (
            .O(N__33457),
            .I(un1_M_this_spr_address_q_cry_8));
    CascadeMux I__7539 (
            .O(N__33454),
            .I(N__33449));
    CascadeMux I__7538 (
            .O(N__33453),
            .I(N__33445));
    CascadeMux I__7537 (
            .O(N__33452),
            .I(N__33440));
    InMux I__7536 (
            .O(N__33449),
            .I(N__33437));
    CascadeMux I__7535 (
            .O(N__33448),
            .I(N__33434));
    InMux I__7534 (
            .O(N__33445),
            .I(N__33427));
    CascadeMux I__7533 (
            .O(N__33444),
            .I(N__33424));
    CascadeMux I__7532 (
            .O(N__33443),
            .I(N__33420));
    InMux I__7531 (
            .O(N__33440),
            .I(N__33416));
    LocalMux I__7530 (
            .O(N__33437),
            .I(N__33413));
    InMux I__7529 (
            .O(N__33434),
            .I(N__33410));
    CascadeMux I__7528 (
            .O(N__33433),
            .I(N__33407));
    CascadeMux I__7527 (
            .O(N__33432),
            .I(N__33404));
    CascadeMux I__7526 (
            .O(N__33431),
            .I(N__33399));
    CascadeMux I__7525 (
            .O(N__33430),
            .I(N__33396));
    LocalMux I__7524 (
            .O(N__33427),
            .I(N__33393));
    InMux I__7523 (
            .O(N__33424),
            .I(N__33390));
    CascadeMux I__7522 (
            .O(N__33423),
            .I(N__33387));
    InMux I__7521 (
            .O(N__33420),
            .I(N__33383));
    CascadeMux I__7520 (
            .O(N__33419),
            .I(N__33380));
    LocalMux I__7519 (
            .O(N__33416),
            .I(N__33373));
    Span4Mux_s1_v I__7518 (
            .O(N__33413),
            .I(N__33373));
    LocalMux I__7517 (
            .O(N__33410),
            .I(N__33373));
    InMux I__7516 (
            .O(N__33407),
            .I(N__33369));
    InMux I__7515 (
            .O(N__33404),
            .I(N__33366));
    CascadeMux I__7514 (
            .O(N__33403),
            .I(N__33363));
    CascadeMux I__7513 (
            .O(N__33402),
            .I(N__33360));
    InMux I__7512 (
            .O(N__33399),
            .I(N__33357));
    InMux I__7511 (
            .O(N__33396),
            .I(N__33354));
    Span4Mux_v I__7510 (
            .O(N__33393),
            .I(N__33349));
    LocalMux I__7509 (
            .O(N__33390),
            .I(N__33349));
    InMux I__7508 (
            .O(N__33387),
            .I(N__33346));
    CascadeMux I__7507 (
            .O(N__33386),
            .I(N__33343));
    LocalMux I__7506 (
            .O(N__33383),
            .I(N__33340));
    InMux I__7505 (
            .O(N__33380),
            .I(N__33337));
    Span4Mux_v I__7504 (
            .O(N__33373),
            .I(N__33334));
    CascadeMux I__7503 (
            .O(N__33372),
            .I(N__33331));
    LocalMux I__7502 (
            .O(N__33369),
            .I(N__33328));
    LocalMux I__7501 (
            .O(N__33366),
            .I(N__33325));
    InMux I__7500 (
            .O(N__33363),
            .I(N__33322));
    InMux I__7499 (
            .O(N__33360),
            .I(N__33319));
    LocalMux I__7498 (
            .O(N__33357),
            .I(N__33316));
    LocalMux I__7497 (
            .O(N__33354),
            .I(N__33313));
    Span4Mux_h I__7496 (
            .O(N__33349),
            .I(N__33310));
    LocalMux I__7495 (
            .O(N__33346),
            .I(N__33307));
    InMux I__7494 (
            .O(N__33343),
            .I(N__33304));
    Span4Mux_v I__7493 (
            .O(N__33340),
            .I(N__33299));
    LocalMux I__7492 (
            .O(N__33337),
            .I(N__33299));
    Span4Mux_h I__7491 (
            .O(N__33334),
            .I(N__33296));
    InMux I__7490 (
            .O(N__33331),
            .I(N__33293));
    Span4Mux_v I__7489 (
            .O(N__33328),
            .I(N__33286));
    Span4Mux_v I__7488 (
            .O(N__33325),
            .I(N__33286));
    LocalMux I__7487 (
            .O(N__33322),
            .I(N__33286));
    LocalMux I__7486 (
            .O(N__33319),
            .I(N__33281));
    Span4Mux_v I__7485 (
            .O(N__33316),
            .I(N__33281));
    Span4Mux_h I__7484 (
            .O(N__33313),
            .I(N__33276));
    Span4Mux_v I__7483 (
            .O(N__33310),
            .I(N__33276));
    Span4Mux_v I__7482 (
            .O(N__33307),
            .I(N__33271));
    LocalMux I__7481 (
            .O(N__33304),
            .I(N__33271));
    Span4Mux_h I__7480 (
            .O(N__33299),
            .I(N__33268));
    Sp12to4 I__7479 (
            .O(N__33296),
            .I(N__33265));
    LocalMux I__7478 (
            .O(N__33293),
            .I(N__33261));
    Span4Mux_h I__7477 (
            .O(N__33286),
            .I(N__33254));
    Span4Mux_h I__7476 (
            .O(N__33281),
            .I(N__33254));
    Span4Mux_v I__7475 (
            .O(N__33276),
            .I(N__33254));
    Span4Mux_h I__7474 (
            .O(N__33271),
            .I(N__33249));
    Span4Mux_v I__7473 (
            .O(N__33268),
            .I(N__33249));
    Span12Mux_v I__7472 (
            .O(N__33265),
            .I(N__33246));
    InMux I__7471 (
            .O(N__33264),
            .I(N__33243));
    Span4Mux_h I__7470 (
            .O(N__33261),
            .I(N__33236));
    Span4Mux_v I__7469 (
            .O(N__33254),
            .I(N__33236));
    Span4Mux_v I__7468 (
            .O(N__33249),
            .I(N__33236));
    Span12Mux_h I__7467 (
            .O(N__33246),
            .I(N__33233));
    LocalMux I__7466 (
            .O(N__33243),
            .I(M_this_spr_address_qZ0Z_10));
    Odrv4 I__7465 (
            .O(N__33236),
            .I(M_this_spr_address_qZ0Z_10));
    Odrv12 I__7464 (
            .O(N__33233),
            .I(M_this_spr_address_qZ0Z_10));
    InMux I__7463 (
            .O(N__33226),
            .I(un1_M_this_spr_address_q_cry_9));
    InMux I__7462 (
            .O(N__33223),
            .I(un1_M_this_spr_address_q_cry_10));
    InMux I__7461 (
            .O(N__33220),
            .I(un1_M_this_spr_address_q_cry_11));
    InMux I__7460 (
            .O(N__33217),
            .I(N__33195));
    InMux I__7459 (
            .O(N__33216),
            .I(N__33195));
    InMux I__7458 (
            .O(N__33215),
            .I(N__33195));
    InMux I__7457 (
            .O(N__33214),
            .I(N__33195));
    InMux I__7456 (
            .O(N__33213),
            .I(N__33186));
    InMux I__7455 (
            .O(N__33212),
            .I(N__33186));
    InMux I__7454 (
            .O(N__33211),
            .I(N__33186));
    InMux I__7453 (
            .O(N__33210),
            .I(N__33186));
    InMux I__7452 (
            .O(N__33209),
            .I(N__33181));
    InMux I__7451 (
            .O(N__33208),
            .I(N__33181));
    InMux I__7450 (
            .O(N__33207),
            .I(N__33172));
    InMux I__7449 (
            .O(N__33206),
            .I(N__33172));
    InMux I__7448 (
            .O(N__33205),
            .I(N__33172));
    InMux I__7447 (
            .O(N__33204),
            .I(N__33172));
    LocalMux I__7446 (
            .O(N__33195),
            .I(N__33165));
    LocalMux I__7445 (
            .O(N__33186),
            .I(N__33165));
    LocalMux I__7444 (
            .O(N__33181),
            .I(N__33160));
    LocalMux I__7443 (
            .O(N__33172),
            .I(N__33160));
    CascadeMux I__7442 (
            .O(N__33171),
            .I(N__33157));
    CascadeMux I__7441 (
            .O(N__33170),
            .I(N__33154));
    Span4Mux_v I__7440 (
            .O(N__33165),
            .I(N__33151));
    Span4Mux_h I__7439 (
            .O(N__33160),
            .I(N__33148));
    InMux I__7438 (
            .O(N__33157),
            .I(N__33145));
    InMux I__7437 (
            .O(N__33154),
            .I(N__33142));
    Sp12to4 I__7436 (
            .O(N__33151),
            .I(N__33139));
    Span4Mux_v I__7435 (
            .O(N__33148),
            .I(N__33136));
    LocalMux I__7434 (
            .O(N__33145),
            .I(N__33133));
    LocalMux I__7433 (
            .O(N__33142),
            .I(N__33128));
    Span12Mux_h I__7432 (
            .O(N__33139),
            .I(N__33128));
    Span4Mux_h I__7431 (
            .O(N__33136),
            .I(N__33125));
    Odrv12 I__7430 (
            .O(N__33133),
            .I(N_1005_0));
    Odrv12 I__7429 (
            .O(N__33128),
            .I(N_1005_0));
    Odrv4 I__7428 (
            .O(N__33125),
            .I(N_1005_0));
    InMux I__7427 (
            .O(N__33118),
            .I(un1_M_this_spr_address_q_cry_12));
    InMux I__7426 (
            .O(N__33115),
            .I(N__33112));
    LocalMux I__7425 (
            .O(N__33112),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_5 ));
    InMux I__7424 (
            .O(N__33109),
            .I(N__33106));
    LocalMux I__7423 (
            .O(N__33106),
            .I(N__33103));
    Span4Mux_v I__7422 (
            .O(N__33103),
            .I(N__33100));
    Sp12to4 I__7421 (
            .O(N__33100),
            .I(N__33097));
    Span12Mux_h I__7420 (
            .O(N__33097),
            .I(N__33094));
    Odrv12 I__7419 (
            .O(N__33094),
            .I(\this_ppu.oam_cache.mem_6 ));
    InMux I__7418 (
            .O(N__33091),
            .I(N__33084));
    InMux I__7417 (
            .O(N__33090),
            .I(N__33081));
    InMux I__7416 (
            .O(N__33089),
            .I(N__33076));
    InMux I__7415 (
            .O(N__33088),
            .I(N__33076));
    CascadeMux I__7414 (
            .O(N__33087),
            .I(N__33070));
    LocalMux I__7413 (
            .O(N__33084),
            .I(N__33063));
    LocalMux I__7412 (
            .O(N__33081),
            .I(N__33063));
    LocalMux I__7411 (
            .O(N__33076),
            .I(N__33063));
    InMux I__7410 (
            .O(N__33075),
            .I(N__33056));
    InMux I__7409 (
            .O(N__33074),
            .I(N__33056));
    InMux I__7408 (
            .O(N__33073),
            .I(N__33056));
    InMux I__7407 (
            .O(N__33070),
            .I(N__33053));
    Span4Mux_v I__7406 (
            .O(N__33063),
            .I(N__33048));
    LocalMux I__7405 (
            .O(N__33056),
            .I(N__33043));
    LocalMux I__7404 (
            .O(N__33053),
            .I(N__33043));
    InMux I__7403 (
            .O(N__33052),
            .I(N__33038));
    InMux I__7402 (
            .O(N__33051),
            .I(N__33038));
    Span4Mux_h I__7401 (
            .O(N__33048),
            .I(N__33031));
    Span4Mux_v I__7400 (
            .O(N__33043),
            .I(N__33031));
    LocalMux I__7399 (
            .O(N__33038),
            .I(N__33031));
    Span4Mux_h I__7398 (
            .O(N__33031),
            .I(N__33028));
    Span4Mux_h I__7397 (
            .O(N__33028),
            .I(N__33025));
    Odrv4 I__7396 (
            .O(N__33025),
            .I(port_address_in_4));
    CascadeMux I__7395 (
            .O(N__33022),
            .I(N__33016));
    InMux I__7394 (
            .O(N__33021),
            .I(N__33008));
    InMux I__7393 (
            .O(N__33020),
            .I(N__33008));
    InMux I__7392 (
            .O(N__33019),
            .I(N__33005));
    InMux I__7391 (
            .O(N__33016),
            .I(N__33000));
    InMux I__7390 (
            .O(N__33015),
            .I(N__33000));
    InMux I__7389 (
            .O(N__33014),
            .I(N__32995));
    InMux I__7388 (
            .O(N__33013),
            .I(N__32995));
    LocalMux I__7387 (
            .O(N__33008),
            .I(N__32990));
    LocalMux I__7386 (
            .O(N__33005),
            .I(N__32990));
    LocalMux I__7385 (
            .O(N__33000),
            .I(N__32982));
    LocalMux I__7384 (
            .O(N__32995),
            .I(N__32982));
    Span4Mux_v I__7383 (
            .O(N__32990),
            .I(N__32977));
    InMux I__7382 (
            .O(N__32989),
            .I(N__32970));
    InMux I__7381 (
            .O(N__32988),
            .I(N__32970));
    InMux I__7380 (
            .O(N__32987),
            .I(N__32970));
    Span4Mux_v I__7379 (
            .O(N__32982),
            .I(N__32967));
    InMux I__7378 (
            .O(N__32981),
            .I(N__32962));
    InMux I__7377 (
            .O(N__32980),
            .I(N__32962));
    Sp12to4 I__7376 (
            .O(N__32977),
            .I(N__32953));
    LocalMux I__7375 (
            .O(N__32970),
            .I(N__32953));
    Sp12to4 I__7374 (
            .O(N__32967),
            .I(N__32953));
    LocalMux I__7373 (
            .O(N__32962),
            .I(N__32953));
    Span12Mux_h I__7372 (
            .O(N__32953),
            .I(N__32950));
    Odrv12 I__7371 (
            .O(N__32950),
            .I(port_address_in_0));
    CascadeMux I__7370 (
            .O(N__32947),
            .I(N__32944));
    InMux I__7369 (
            .O(N__32944),
            .I(N__32939));
    CascadeMux I__7368 (
            .O(N__32943),
            .I(N__32936));
    CascadeMux I__7367 (
            .O(N__32942),
            .I(N__32929));
    LocalMux I__7366 (
            .O(N__32939),
            .I(N__32924));
    InMux I__7365 (
            .O(N__32936),
            .I(N__32921));
    InMux I__7364 (
            .O(N__32935),
            .I(N__32916));
    InMux I__7363 (
            .O(N__32934),
            .I(N__32916));
    InMux I__7362 (
            .O(N__32933),
            .I(N__32913));
    InMux I__7361 (
            .O(N__32932),
            .I(N__32908));
    InMux I__7360 (
            .O(N__32929),
            .I(N__32908));
    InMux I__7359 (
            .O(N__32928),
            .I(N__32903));
    InMux I__7358 (
            .O(N__32927),
            .I(N__32903));
    Span4Mux_h I__7357 (
            .O(N__32924),
            .I(N__32890));
    LocalMux I__7356 (
            .O(N__32921),
            .I(N__32890));
    LocalMux I__7355 (
            .O(N__32916),
            .I(N__32890));
    LocalMux I__7354 (
            .O(N__32913),
            .I(N__32890));
    LocalMux I__7353 (
            .O(N__32908),
            .I(N__32890));
    LocalMux I__7352 (
            .O(N__32903),
            .I(N__32890));
    Span4Mux_v I__7351 (
            .O(N__32890),
            .I(N__32887));
    Span4Mux_h I__7350 (
            .O(N__32887),
            .I(N__32884));
    Span4Mux_v I__7349 (
            .O(N__32884),
            .I(N__32881));
    Sp12to4 I__7348 (
            .O(N__32881),
            .I(N__32878));
    Span12Mux_h I__7347 (
            .O(N__32878),
            .I(N__32874));
    InMux I__7346 (
            .O(N__32877),
            .I(N__32871));
    Odrv12 I__7345 (
            .O(N__32874),
            .I(port_rw_in));
    LocalMux I__7344 (
            .O(N__32871),
            .I(port_rw_in));
    CascadeMux I__7343 (
            .O(N__32866),
            .I(N__32863));
    InMux I__7342 (
            .O(N__32863),
            .I(N__32860));
    LocalMux I__7341 (
            .O(N__32860),
            .I(N__32857));
    Span4Mux_h I__7340 (
            .O(N__32857),
            .I(N__32853));
    InMux I__7339 (
            .O(N__32856),
            .I(N__32850));
    Odrv4 I__7338 (
            .O(N__32853),
            .I(N_1422));
    LocalMux I__7337 (
            .O(N__32850),
            .I(N_1422));
    CascadeMux I__7336 (
            .O(N__32845),
            .I(N__32840));
    CascadeMux I__7335 (
            .O(N__32844),
            .I(N__32834));
    CascadeMux I__7334 (
            .O(N__32843),
            .I(N__32831));
    InMux I__7333 (
            .O(N__32840),
            .I(N__32827));
    CascadeMux I__7332 (
            .O(N__32839),
            .I(N__32824));
    CascadeMux I__7331 (
            .O(N__32838),
            .I(N__32820));
    CascadeMux I__7330 (
            .O(N__32837),
            .I(N__32817));
    InMux I__7329 (
            .O(N__32834),
            .I(N__32812));
    InMux I__7328 (
            .O(N__32831),
            .I(N__32809));
    CascadeMux I__7327 (
            .O(N__32830),
            .I(N__32806));
    LocalMux I__7326 (
            .O(N__32827),
            .I(N__32803));
    InMux I__7325 (
            .O(N__32824),
            .I(N__32800));
    CascadeMux I__7324 (
            .O(N__32823),
            .I(N__32797));
    InMux I__7323 (
            .O(N__32820),
            .I(N__32793));
    InMux I__7322 (
            .O(N__32817),
            .I(N__32790));
    CascadeMux I__7321 (
            .O(N__32816),
            .I(N__32787));
    CascadeMux I__7320 (
            .O(N__32815),
            .I(N__32784));
    LocalMux I__7319 (
            .O(N__32812),
            .I(N__32779));
    LocalMux I__7318 (
            .O(N__32809),
            .I(N__32776));
    InMux I__7317 (
            .O(N__32806),
            .I(N__32773));
    Span4Mux_h I__7316 (
            .O(N__32803),
            .I(N__32768));
    LocalMux I__7315 (
            .O(N__32800),
            .I(N__32768));
    InMux I__7314 (
            .O(N__32797),
            .I(N__32765));
    CascadeMux I__7313 (
            .O(N__32796),
            .I(N__32762));
    LocalMux I__7312 (
            .O(N__32793),
            .I(N__32758));
    LocalMux I__7311 (
            .O(N__32790),
            .I(N__32755));
    InMux I__7310 (
            .O(N__32787),
            .I(N__32752));
    InMux I__7309 (
            .O(N__32784),
            .I(N__32749));
    CascadeMux I__7308 (
            .O(N__32783),
            .I(N__32746));
    CascadeMux I__7307 (
            .O(N__32782),
            .I(N__32743));
    Span4Mux_s2_v I__7306 (
            .O(N__32779),
            .I(N__32735));
    Span4Mux_h I__7305 (
            .O(N__32776),
            .I(N__32735));
    LocalMux I__7304 (
            .O(N__32773),
            .I(N__32735));
    Span4Mux_v I__7303 (
            .O(N__32768),
            .I(N__32730));
    LocalMux I__7302 (
            .O(N__32765),
            .I(N__32730));
    InMux I__7301 (
            .O(N__32762),
            .I(N__32727));
    CascadeMux I__7300 (
            .O(N__32761),
            .I(N__32724));
    Span4Mux_v I__7299 (
            .O(N__32758),
            .I(N__32715));
    Span4Mux_v I__7298 (
            .O(N__32755),
            .I(N__32715));
    LocalMux I__7297 (
            .O(N__32752),
            .I(N__32715));
    LocalMux I__7296 (
            .O(N__32749),
            .I(N__32715));
    InMux I__7295 (
            .O(N__32746),
            .I(N__32712));
    InMux I__7294 (
            .O(N__32743),
            .I(N__32709));
    CascadeMux I__7293 (
            .O(N__32742),
            .I(N__32706));
    Span4Mux_v I__7292 (
            .O(N__32735),
            .I(N__32703));
    Span4Mux_h I__7291 (
            .O(N__32730),
            .I(N__32697));
    LocalMux I__7290 (
            .O(N__32727),
            .I(N__32697));
    InMux I__7289 (
            .O(N__32724),
            .I(N__32694));
    Span4Mux_v I__7288 (
            .O(N__32715),
            .I(N__32687));
    LocalMux I__7287 (
            .O(N__32712),
            .I(N__32687));
    LocalMux I__7286 (
            .O(N__32709),
            .I(N__32687));
    InMux I__7285 (
            .O(N__32706),
            .I(N__32684));
    Sp12to4 I__7284 (
            .O(N__32703),
            .I(N__32681));
    CascadeMux I__7283 (
            .O(N__32702),
            .I(N__32678));
    Span4Mux_v I__7282 (
            .O(N__32697),
            .I(N__32673));
    LocalMux I__7281 (
            .O(N__32694),
            .I(N__32673));
    Span4Mux_v I__7280 (
            .O(N__32687),
            .I(N__32668));
    LocalMux I__7279 (
            .O(N__32684),
            .I(N__32668));
    Span12Mux_h I__7278 (
            .O(N__32681),
            .I(N__32665));
    InMux I__7277 (
            .O(N__32678),
            .I(N__32662));
    Span4Mux_h I__7276 (
            .O(N__32673),
            .I(N__32656));
    Span4Mux_h I__7275 (
            .O(N__32668),
            .I(N__32656));
    Span12Mux_v I__7274 (
            .O(N__32665),
            .I(N__32651));
    LocalMux I__7273 (
            .O(N__32662),
            .I(N__32651));
    InMux I__7272 (
            .O(N__32661),
            .I(N__32648));
    Odrv4 I__7271 (
            .O(N__32656),
            .I(M_this_spr_address_qZ0Z_0));
    Odrv12 I__7270 (
            .O(N__32651),
            .I(M_this_spr_address_qZ0Z_0));
    LocalMux I__7269 (
            .O(N__32648),
            .I(M_this_spr_address_qZ0Z_0));
    CascadeMux I__7268 (
            .O(N__32641),
            .I(N__32638));
    InMux I__7267 (
            .O(N__32638),
            .I(N__32627));
    CascadeMux I__7266 (
            .O(N__32637),
            .I(N__32624));
    CascadeMux I__7265 (
            .O(N__32636),
            .I(N__32620));
    CascadeMux I__7264 (
            .O(N__32635),
            .I(N__32617));
    CascadeMux I__7263 (
            .O(N__32634),
            .I(N__32614));
    CascadeMux I__7262 (
            .O(N__32633),
            .I(N__32610));
    CascadeMux I__7261 (
            .O(N__32632),
            .I(N__32606));
    CascadeMux I__7260 (
            .O(N__32631),
            .I(N__32603));
    CascadeMux I__7259 (
            .O(N__32630),
            .I(N__32598));
    LocalMux I__7258 (
            .O(N__32627),
            .I(N__32595));
    InMux I__7257 (
            .O(N__32624),
            .I(N__32592));
    CascadeMux I__7256 (
            .O(N__32623),
            .I(N__32589));
    InMux I__7255 (
            .O(N__32620),
            .I(N__32586));
    InMux I__7254 (
            .O(N__32617),
            .I(N__32583));
    InMux I__7253 (
            .O(N__32614),
            .I(N__32580));
    CascadeMux I__7252 (
            .O(N__32613),
            .I(N__32576));
    InMux I__7251 (
            .O(N__32610),
            .I(N__32573));
    CascadeMux I__7250 (
            .O(N__32609),
            .I(N__32570));
    InMux I__7249 (
            .O(N__32606),
            .I(N__32567));
    InMux I__7248 (
            .O(N__32603),
            .I(N__32564));
    CascadeMux I__7247 (
            .O(N__32602),
            .I(N__32561));
    CascadeMux I__7246 (
            .O(N__32601),
            .I(N__32558));
    InMux I__7245 (
            .O(N__32598),
            .I(N__32555));
    Span4Mux_v I__7244 (
            .O(N__32595),
            .I(N__32550));
    LocalMux I__7243 (
            .O(N__32592),
            .I(N__32550));
    InMux I__7242 (
            .O(N__32589),
            .I(N__32547));
    LocalMux I__7241 (
            .O(N__32586),
            .I(N__32544));
    LocalMux I__7240 (
            .O(N__32583),
            .I(N__32541));
    LocalMux I__7239 (
            .O(N__32580),
            .I(N__32538));
    CascadeMux I__7238 (
            .O(N__32579),
            .I(N__32534));
    InMux I__7237 (
            .O(N__32576),
            .I(N__32531));
    LocalMux I__7236 (
            .O(N__32573),
            .I(N__32528));
    InMux I__7235 (
            .O(N__32570),
            .I(N__32525));
    LocalMux I__7234 (
            .O(N__32567),
            .I(N__32520));
    LocalMux I__7233 (
            .O(N__32564),
            .I(N__32520));
    InMux I__7232 (
            .O(N__32561),
            .I(N__32517));
    InMux I__7231 (
            .O(N__32558),
            .I(N__32514));
    LocalMux I__7230 (
            .O(N__32555),
            .I(N__32511));
    Span4Mux_h I__7229 (
            .O(N__32550),
            .I(N__32508));
    LocalMux I__7228 (
            .O(N__32547),
            .I(N__32505));
    Span4Mux_h I__7227 (
            .O(N__32544),
            .I(N__32502));
    Span4Mux_h I__7226 (
            .O(N__32541),
            .I(N__32499));
    Span4Mux_h I__7225 (
            .O(N__32538),
            .I(N__32496));
    CascadeMux I__7224 (
            .O(N__32537),
            .I(N__32493));
    InMux I__7223 (
            .O(N__32534),
            .I(N__32490));
    LocalMux I__7222 (
            .O(N__32531),
            .I(N__32487));
    Span4Mux_v I__7221 (
            .O(N__32528),
            .I(N__32482));
    LocalMux I__7220 (
            .O(N__32525),
            .I(N__32482));
    Span4Mux_v I__7219 (
            .O(N__32520),
            .I(N__32477));
    LocalMux I__7218 (
            .O(N__32517),
            .I(N__32477));
    LocalMux I__7217 (
            .O(N__32514),
            .I(N__32474));
    Span4Mux_h I__7216 (
            .O(N__32511),
            .I(N__32471));
    Span4Mux_h I__7215 (
            .O(N__32508),
            .I(N__32466));
    Span4Mux_h I__7214 (
            .O(N__32505),
            .I(N__32466));
    Sp12to4 I__7213 (
            .O(N__32502),
            .I(N__32459));
    Sp12to4 I__7212 (
            .O(N__32499),
            .I(N__32459));
    Sp12to4 I__7211 (
            .O(N__32496),
            .I(N__32459));
    InMux I__7210 (
            .O(N__32493),
            .I(N__32456));
    LocalMux I__7209 (
            .O(N__32490),
            .I(N__32453));
    Span4Mux_h I__7208 (
            .O(N__32487),
            .I(N__32448));
    Span4Mux_h I__7207 (
            .O(N__32482),
            .I(N__32448));
    Span4Mux_h I__7206 (
            .O(N__32477),
            .I(N__32445));
    Span4Mux_h I__7205 (
            .O(N__32474),
            .I(N__32442));
    Sp12to4 I__7204 (
            .O(N__32471),
            .I(N__32436));
    Sp12to4 I__7203 (
            .O(N__32466),
            .I(N__32436));
    Span12Mux_s9_v I__7202 (
            .O(N__32459),
            .I(N__32433));
    LocalMux I__7201 (
            .O(N__32456),
            .I(N__32430));
    Span4Mux_h I__7200 (
            .O(N__32453),
            .I(N__32425));
    Span4Mux_v I__7199 (
            .O(N__32448),
            .I(N__32425));
    Span4Mux_v I__7198 (
            .O(N__32445),
            .I(N__32422));
    Sp12to4 I__7197 (
            .O(N__32442),
            .I(N__32419));
    InMux I__7196 (
            .O(N__32441),
            .I(N__32416));
    Span12Mux_s9_v I__7195 (
            .O(N__32436),
            .I(N__32411));
    Span12Mux_h I__7194 (
            .O(N__32433),
            .I(N__32411));
    Odrv4 I__7193 (
            .O(N__32430),
            .I(M_this_spr_address_qZ0Z_1));
    Odrv4 I__7192 (
            .O(N__32425),
            .I(M_this_spr_address_qZ0Z_1));
    Odrv4 I__7191 (
            .O(N__32422),
            .I(M_this_spr_address_qZ0Z_1));
    Odrv12 I__7190 (
            .O(N__32419),
            .I(M_this_spr_address_qZ0Z_1));
    LocalMux I__7189 (
            .O(N__32416),
            .I(M_this_spr_address_qZ0Z_1));
    Odrv12 I__7188 (
            .O(N__32411),
            .I(M_this_spr_address_qZ0Z_1));
    InMux I__7187 (
            .O(N__32398),
            .I(un1_M_this_spr_address_q_cry_0));
    CascadeMux I__7186 (
            .O(N__32395),
            .I(N__32392));
    InMux I__7185 (
            .O(N__32392),
            .I(N__32387));
    CascadeMux I__7184 (
            .O(N__32391),
            .I(N__32384));
    CascadeMux I__7183 (
            .O(N__32390),
            .I(N__32381));
    LocalMux I__7182 (
            .O(N__32387),
            .I(N__32376));
    InMux I__7181 (
            .O(N__32384),
            .I(N__32373));
    InMux I__7180 (
            .O(N__32381),
            .I(N__32369));
    CascadeMux I__7179 (
            .O(N__32380),
            .I(N__32366));
    CascadeMux I__7178 (
            .O(N__32379),
            .I(N__32362));
    Span4Mux_h I__7177 (
            .O(N__32376),
            .I(N__32355));
    LocalMux I__7176 (
            .O(N__32373),
            .I(N__32355));
    CascadeMux I__7175 (
            .O(N__32372),
            .I(N__32352));
    LocalMux I__7174 (
            .O(N__32369),
            .I(N__32349));
    InMux I__7173 (
            .O(N__32366),
            .I(N__32346));
    CascadeMux I__7172 (
            .O(N__32365),
            .I(N__32343));
    InMux I__7171 (
            .O(N__32362),
            .I(N__32339));
    CascadeMux I__7170 (
            .O(N__32361),
            .I(N__32336));
    CascadeMux I__7169 (
            .O(N__32360),
            .I(N__32333));
    Span4Mux_v I__7168 (
            .O(N__32355),
            .I(N__32328));
    InMux I__7167 (
            .O(N__32352),
            .I(N__32325));
    Span4Mux_v I__7166 (
            .O(N__32349),
            .I(N__32320));
    LocalMux I__7165 (
            .O(N__32346),
            .I(N__32320));
    InMux I__7164 (
            .O(N__32343),
            .I(N__32317));
    CascadeMux I__7163 (
            .O(N__32342),
            .I(N__32314));
    LocalMux I__7162 (
            .O(N__32339),
            .I(N__32310));
    InMux I__7161 (
            .O(N__32336),
            .I(N__32307));
    InMux I__7160 (
            .O(N__32333),
            .I(N__32304));
    CascadeMux I__7159 (
            .O(N__32332),
            .I(N__32301));
    CascadeMux I__7158 (
            .O(N__32331),
            .I(N__32298));
    Sp12to4 I__7157 (
            .O(N__32328),
            .I(N__32293));
    LocalMux I__7156 (
            .O(N__32325),
            .I(N__32290));
    Span4Mux_h I__7155 (
            .O(N__32320),
            .I(N__32285));
    LocalMux I__7154 (
            .O(N__32317),
            .I(N__32285));
    InMux I__7153 (
            .O(N__32314),
            .I(N__32282));
    CascadeMux I__7152 (
            .O(N__32313),
            .I(N__32279));
    Span4Mux_v I__7151 (
            .O(N__32310),
            .I(N__32272));
    LocalMux I__7150 (
            .O(N__32307),
            .I(N__32272));
    LocalMux I__7149 (
            .O(N__32304),
            .I(N__32272));
    InMux I__7148 (
            .O(N__32301),
            .I(N__32269));
    InMux I__7147 (
            .O(N__32298),
            .I(N__32266));
    CascadeMux I__7146 (
            .O(N__32297),
            .I(N__32263));
    CascadeMux I__7145 (
            .O(N__32296),
            .I(N__32260));
    Span12Mux_h I__7144 (
            .O(N__32293),
            .I(N__32254));
    Span12Mux_s9_h I__7143 (
            .O(N__32290),
            .I(N__32254));
    Span4Mux_v I__7142 (
            .O(N__32285),
            .I(N__32249));
    LocalMux I__7141 (
            .O(N__32282),
            .I(N__32249));
    InMux I__7140 (
            .O(N__32279),
            .I(N__32246));
    Span4Mux_v I__7139 (
            .O(N__32272),
            .I(N__32239));
    LocalMux I__7138 (
            .O(N__32269),
            .I(N__32239));
    LocalMux I__7137 (
            .O(N__32266),
            .I(N__32239));
    InMux I__7136 (
            .O(N__32263),
            .I(N__32236));
    InMux I__7135 (
            .O(N__32260),
            .I(N__32233));
    CascadeMux I__7134 (
            .O(N__32259),
            .I(N__32230));
    Span12Mux_v I__7133 (
            .O(N__32254),
            .I(N__32227));
    Span4Mux_h I__7132 (
            .O(N__32249),
            .I(N__32222));
    LocalMux I__7131 (
            .O(N__32246),
            .I(N__32222));
    Span4Mux_v I__7130 (
            .O(N__32239),
            .I(N__32215));
    LocalMux I__7129 (
            .O(N__32236),
            .I(N__32215));
    LocalMux I__7128 (
            .O(N__32233),
            .I(N__32215));
    InMux I__7127 (
            .O(N__32230),
            .I(N__32212));
    Span12Mux_h I__7126 (
            .O(N__32227),
            .I(N__32208));
    Span4Mux_v I__7125 (
            .O(N__32222),
            .I(N__32201));
    Span4Mux_v I__7124 (
            .O(N__32215),
            .I(N__32201));
    LocalMux I__7123 (
            .O(N__32212),
            .I(N__32201));
    InMux I__7122 (
            .O(N__32211),
            .I(N__32198));
    Odrv12 I__7121 (
            .O(N__32208),
            .I(M_this_spr_address_qZ0Z_2));
    Odrv4 I__7120 (
            .O(N__32201),
            .I(M_this_spr_address_qZ0Z_2));
    LocalMux I__7119 (
            .O(N__32198),
            .I(M_this_spr_address_qZ0Z_2));
    InMux I__7118 (
            .O(N__32191),
            .I(un1_M_this_spr_address_q_cry_1));
    CascadeMux I__7117 (
            .O(N__32188),
            .I(N__32184));
    CascadeMux I__7116 (
            .O(N__32187),
            .I(N__32179));
    InMux I__7115 (
            .O(N__32184),
            .I(N__32176));
    CascadeMux I__7114 (
            .O(N__32183),
            .I(N__32173));
    CascadeMux I__7113 (
            .O(N__32182),
            .I(N__32167));
    InMux I__7112 (
            .O(N__32179),
            .I(N__32163));
    LocalMux I__7111 (
            .O(N__32176),
            .I(N__32160));
    InMux I__7110 (
            .O(N__32173),
            .I(N__32157));
    CascadeMux I__7109 (
            .O(N__32172),
            .I(N__32154));
    CascadeMux I__7108 (
            .O(N__32171),
            .I(N__32151));
    CascadeMux I__7107 (
            .O(N__32170),
            .I(N__32146));
    InMux I__7106 (
            .O(N__32167),
            .I(N__32143));
    CascadeMux I__7105 (
            .O(N__32166),
            .I(N__32140));
    LocalMux I__7104 (
            .O(N__32163),
            .I(N__32135));
    Span4Mux_h I__7103 (
            .O(N__32160),
            .I(N__32132));
    LocalMux I__7102 (
            .O(N__32157),
            .I(N__32129));
    InMux I__7101 (
            .O(N__32154),
            .I(N__32126));
    InMux I__7100 (
            .O(N__32151),
            .I(N__32123));
    CascadeMux I__7099 (
            .O(N__32150),
            .I(N__32120));
    CascadeMux I__7098 (
            .O(N__32149),
            .I(N__32117));
    InMux I__7097 (
            .O(N__32146),
            .I(N__32113));
    LocalMux I__7096 (
            .O(N__32143),
            .I(N__32110));
    InMux I__7095 (
            .O(N__32140),
            .I(N__32107));
    CascadeMux I__7094 (
            .O(N__32139),
            .I(N__32104));
    CascadeMux I__7093 (
            .O(N__32138),
            .I(N__32101));
    Span4Mux_h I__7092 (
            .O(N__32135),
            .I(N__32096));
    Span4Mux_v I__7091 (
            .O(N__32132),
            .I(N__32091));
    Span4Mux_h I__7090 (
            .O(N__32129),
            .I(N__32091));
    LocalMux I__7089 (
            .O(N__32126),
            .I(N__32088));
    LocalMux I__7088 (
            .O(N__32123),
            .I(N__32085));
    InMux I__7087 (
            .O(N__32120),
            .I(N__32082));
    InMux I__7086 (
            .O(N__32117),
            .I(N__32079));
    CascadeMux I__7085 (
            .O(N__32116),
            .I(N__32076));
    LocalMux I__7084 (
            .O(N__32113),
            .I(N__32073));
    Span4Mux_v I__7083 (
            .O(N__32110),
            .I(N__32068));
    LocalMux I__7082 (
            .O(N__32107),
            .I(N__32068));
    InMux I__7081 (
            .O(N__32104),
            .I(N__32065));
    InMux I__7080 (
            .O(N__32101),
            .I(N__32062));
    CascadeMux I__7079 (
            .O(N__32100),
            .I(N__32059));
    CascadeMux I__7078 (
            .O(N__32099),
            .I(N__32056));
    Sp12to4 I__7077 (
            .O(N__32096),
            .I(N__32050));
    Sp12to4 I__7076 (
            .O(N__32091),
            .I(N__32050));
    Span4Mux_v I__7075 (
            .O(N__32088),
            .I(N__32043));
    Span4Mux_h I__7074 (
            .O(N__32085),
            .I(N__32043));
    LocalMux I__7073 (
            .O(N__32082),
            .I(N__32043));
    LocalMux I__7072 (
            .O(N__32079),
            .I(N__32040));
    InMux I__7071 (
            .O(N__32076),
            .I(N__32037));
    Span4Mux_v I__7070 (
            .O(N__32073),
            .I(N__32028));
    Span4Mux_v I__7069 (
            .O(N__32068),
            .I(N__32028));
    LocalMux I__7068 (
            .O(N__32065),
            .I(N__32028));
    LocalMux I__7067 (
            .O(N__32062),
            .I(N__32028));
    InMux I__7066 (
            .O(N__32059),
            .I(N__32025));
    InMux I__7065 (
            .O(N__32056),
            .I(N__32022));
    CascadeMux I__7064 (
            .O(N__32055),
            .I(N__32019));
    Span12Mux_v I__7063 (
            .O(N__32050),
            .I(N__32016));
    Span4Mux_v I__7062 (
            .O(N__32043),
            .I(N__32009));
    Span4Mux_h I__7061 (
            .O(N__32040),
            .I(N__32009));
    LocalMux I__7060 (
            .O(N__32037),
            .I(N__32009));
    Span4Mux_v I__7059 (
            .O(N__32028),
            .I(N__32002));
    LocalMux I__7058 (
            .O(N__32025),
            .I(N__32002));
    LocalMux I__7057 (
            .O(N__32022),
            .I(N__32002));
    InMux I__7056 (
            .O(N__32019),
            .I(N__31999));
    Span12Mux_h I__7055 (
            .O(N__32016),
            .I(N__31995));
    Span4Mux_v I__7054 (
            .O(N__32009),
            .I(N__31990));
    Span4Mux_v I__7053 (
            .O(N__32002),
            .I(N__31990));
    LocalMux I__7052 (
            .O(N__31999),
            .I(N__31987));
    InMux I__7051 (
            .O(N__31998),
            .I(N__31984));
    Odrv12 I__7050 (
            .O(N__31995),
            .I(M_this_spr_address_qZ0Z_3));
    Odrv4 I__7049 (
            .O(N__31990),
            .I(M_this_spr_address_qZ0Z_3));
    Odrv12 I__7048 (
            .O(N__31987),
            .I(M_this_spr_address_qZ0Z_3));
    LocalMux I__7047 (
            .O(N__31984),
            .I(M_this_spr_address_qZ0Z_3));
    InMux I__7046 (
            .O(N__31975),
            .I(un1_M_this_spr_address_q_cry_2));
    CascadeMux I__7045 (
            .O(N__31972),
            .I(N__31967));
    CascadeMux I__7044 (
            .O(N__31971),
            .I(N__31963));
    CascadeMux I__7043 (
            .O(N__31970),
            .I(N__31958));
    InMux I__7042 (
            .O(N__31967),
            .I(N__31955));
    CascadeMux I__7041 (
            .O(N__31966),
            .I(N__31952));
    InMux I__7040 (
            .O(N__31963),
            .I(N__31949));
    CascadeMux I__7039 (
            .O(N__31962),
            .I(N__31946));
    CascadeMux I__7038 (
            .O(N__31961),
            .I(N__31942));
    InMux I__7037 (
            .O(N__31958),
            .I(N__31937));
    LocalMux I__7036 (
            .O(N__31955),
            .I(N__31934));
    InMux I__7035 (
            .O(N__31952),
            .I(N__31931));
    LocalMux I__7034 (
            .O(N__31949),
            .I(N__31928));
    InMux I__7033 (
            .O(N__31946),
            .I(N__31925));
    CascadeMux I__7032 (
            .O(N__31945),
            .I(N__31922));
    InMux I__7031 (
            .O(N__31942),
            .I(N__31918));
    CascadeMux I__7030 (
            .O(N__31941),
            .I(N__31915));
    CascadeMux I__7029 (
            .O(N__31940),
            .I(N__31912));
    LocalMux I__7028 (
            .O(N__31937),
            .I(N__31906));
    Span4Mux_h I__7027 (
            .O(N__31934),
            .I(N__31903));
    LocalMux I__7026 (
            .O(N__31931),
            .I(N__31900));
    Span4Mux_v I__7025 (
            .O(N__31928),
            .I(N__31895));
    LocalMux I__7024 (
            .O(N__31925),
            .I(N__31895));
    InMux I__7023 (
            .O(N__31922),
            .I(N__31892));
    CascadeMux I__7022 (
            .O(N__31921),
            .I(N__31889));
    LocalMux I__7021 (
            .O(N__31918),
            .I(N__31885));
    InMux I__7020 (
            .O(N__31915),
            .I(N__31882));
    InMux I__7019 (
            .O(N__31912),
            .I(N__31879));
    CascadeMux I__7018 (
            .O(N__31911),
            .I(N__31876));
    CascadeMux I__7017 (
            .O(N__31910),
            .I(N__31873));
    CascadeMux I__7016 (
            .O(N__31909),
            .I(N__31870));
    Span4Mux_h I__7015 (
            .O(N__31906),
            .I(N__31866));
    Span4Mux_v I__7014 (
            .O(N__31903),
            .I(N__31861));
    Span4Mux_h I__7013 (
            .O(N__31900),
            .I(N__31861));
    Span4Mux_h I__7012 (
            .O(N__31895),
            .I(N__31856));
    LocalMux I__7011 (
            .O(N__31892),
            .I(N__31856));
    InMux I__7010 (
            .O(N__31889),
            .I(N__31853));
    CascadeMux I__7009 (
            .O(N__31888),
            .I(N__31850));
    Span4Mux_v I__7008 (
            .O(N__31885),
            .I(N__31843));
    LocalMux I__7007 (
            .O(N__31882),
            .I(N__31843));
    LocalMux I__7006 (
            .O(N__31879),
            .I(N__31843));
    InMux I__7005 (
            .O(N__31876),
            .I(N__31840));
    InMux I__7004 (
            .O(N__31873),
            .I(N__31837));
    InMux I__7003 (
            .O(N__31870),
            .I(N__31834));
    CascadeMux I__7002 (
            .O(N__31869),
            .I(N__31831));
    Sp12to4 I__7001 (
            .O(N__31866),
            .I(N__31825));
    Sp12to4 I__7000 (
            .O(N__31861),
            .I(N__31825));
    Span4Mux_v I__6999 (
            .O(N__31856),
            .I(N__31820));
    LocalMux I__6998 (
            .O(N__31853),
            .I(N__31820));
    InMux I__6997 (
            .O(N__31850),
            .I(N__31817));
    Span4Mux_v I__6996 (
            .O(N__31843),
            .I(N__31812));
    LocalMux I__6995 (
            .O(N__31840),
            .I(N__31812));
    LocalMux I__6994 (
            .O(N__31837),
            .I(N__31809));
    LocalMux I__6993 (
            .O(N__31834),
            .I(N__31806));
    InMux I__6992 (
            .O(N__31831),
            .I(N__31803));
    CascadeMux I__6991 (
            .O(N__31830),
            .I(N__31800));
    Span12Mux_v I__6990 (
            .O(N__31825),
            .I(N__31797));
    Span4Mux_h I__6989 (
            .O(N__31820),
            .I(N__31792));
    LocalMux I__6988 (
            .O(N__31817),
            .I(N__31792));
    Span4Mux_v I__6987 (
            .O(N__31812),
            .I(N__31783));
    Span4Mux_v I__6986 (
            .O(N__31809),
            .I(N__31783));
    Span4Mux_h I__6985 (
            .O(N__31806),
            .I(N__31783));
    LocalMux I__6984 (
            .O(N__31803),
            .I(N__31783));
    InMux I__6983 (
            .O(N__31800),
            .I(N__31780));
    Span12Mux_h I__6982 (
            .O(N__31797),
            .I(N__31776));
    Span4Mux_v I__6981 (
            .O(N__31792),
            .I(N__31769));
    Span4Mux_v I__6980 (
            .O(N__31783),
            .I(N__31769));
    LocalMux I__6979 (
            .O(N__31780),
            .I(N__31769));
    InMux I__6978 (
            .O(N__31779),
            .I(N__31766));
    Odrv12 I__6977 (
            .O(N__31776),
            .I(M_this_spr_address_qZ0Z_4));
    Odrv4 I__6976 (
            .O(N__31769),
            .I(M_this_spr_address_qZ0Z_4));
    LocalMux I__6975 (
            .O(N__31766),
            .I(M_this_spr_address_qZ0Z_4));
    InMux I__6974 (
            .O(N__31759),
            .I(un1_M_this_spr_address_q_cry_3));
    CascadeMux I__6973 (
            .O(N__31756),
            .I(N__31752));
    CascadeMux I__6972 (
            .O(N__31755),
            .I(N__31749));
    InMux I__6971 (
            .O(N__31752),
            .I(N__31743));
    InMux I__6970 (
            .O(N__31749),
            .I(N__31740));
    CascadeMux I__6969 (
            .O(N__31748),
            .I(N__31737));
    CascadeMux I__6968 (
            .O(N__31747),
            .I(N__31732));
    CascadeMux I__6967 (
            .O(N__31746),
            .I(N__31729));
    LocalMux I__6966 (
            .O(N__31743),
            .I(N__31724));
    LocalMux I__6965 (
            .O(N__31740),
            .I(N__31721));
    InMux I__6964 (
            .O(N__31737),
            .I(N__31718));
    CascadeMux I__6963 (
            .O(N__31736),
            .I(N__31715));
    CascadeMux I__6962 (
            .O(N__31735),
            .I(N__31709));
    InMux I__6961 (
            .O(N__31732),
            .I(N__31704));
    InMux I__6960 (
            .O(N__31729),
            .I(N__31701));
    CascadeMux I__6959 (
            .O(N__31728),
            .I(N__31698));
    CascadeMux I__6958 (
            .O(N__31727),
            .I(N__31695));
    Span4Mux_s2_v I__6957 (
            .O(N__31724),
            .I(N__31687));
    Span4Mux_h I__6956 (
            .O(N__31721),
            .I(N__31687));
    LocalMux I__6955 (
            .O(N__31718),
            .I(N__31687));
    InMux I__6954 (
            .O(N__31715),
            .I(N__31684));
    CascadeMux I__6953 (
            .O(N__31714),
            .I(N__31681));
    CascadeMux I__6952 (
            .O(N__31713),
            .I(N__31678));
    CascadeMux I__6951 (
            .O(N__31712),
            .I(N__31675));
    InMux I__6950 (
            .O(N__31709),
            .I(N__31672));
    CascadeMux I__6949 (
            .O(N__31708),
            .I(N__31669));
    CascadeMux I__6948 (
            .O(N__31707),
            .I(N__31666));
    LocalMux I__6947 (
            .O(N__31704),
            .I(N__31661));
    LocalMux I__6946 (
            .O(N__31701),
            .I(N__31661));
    InMux I__6945 (
            .O(N__31698),
            .I(N__31658));
    InMux I__6944 (
            .O(N__31695),
            .I(N__31655));
    CascadeMux I__6943 (
            .O(N__31694),
            .I(N__31652));
    Span4Mux_v I__6942 (
            .O(N__31687),
            .I(N__31649));
    LocalMux I__6941 (
            .O(N__31684),
            .I(N__31645));
    InMux I__6940 (
            .O(N__31681),
            .I(N__31642));
    InMux I__6939 (
            .O(N__31678),
            .I(N__31639));
    InMux I__6938 (
            .O(N__31675),
            .I(N__31636));
    LocalMux I__6937 (
            .O(N__31672),
            .I(N__31633));
    InMux I__6936 (
            .O(N__31669),
            .I(N__31630));
    InMux I__6935 (
            .O(N__31666),
            .I(N__31627));
    Span4Mux_v I__6934 (
            .O(N__31661),
            .I(N__31620));
    LocalMux I__6933 (
            .O(N__31658),
            .I(N__31620));
    LocalMux I__6932 (
            .O(N__31655),
            .I(N__31620));
    InMux I__6931 (
            .O(N__31652),
            .I(N__31617));
    Sp12to4 I__6930 (
            .O(N__31649),
            .I(N__31614));
    CascadeMux I__6929 (
            .O(N__31648),
            .I(N__31611));
    Span12Mux_s6_v I__6928 (
            .O(N__31645),
            .I(N__31606));
    LocalMux I__6927 (
            .O(N__31642),
            .I(N__31606));
    LocalMux I__6926 (
            .O(N__31639),
            .I(N__31601));
    LocalMux I__6925 (
            .O(N__31636),
            .I(N__31601));
    Span4Mux_v I__6924 (
            .O(N__31633),
            .I(N__31596));
    LocalMux I__6923 (
            .O(N__31630),
            .I(N__31596));
    LocalMux I__6922 (
            .O(N__31627),
            .I(N__31593));
    Span4Mux_v I__6921 (
            .O(N__31620),
            .I(N__31588));
    LocalMux I__6920 (
            .O(N__31617),
            .I(N__31588));
    Span12Mux_h I__6919 (
            .O(N__31614),
            .I(N__31585));
    InMux I__6918 (
            .O(N__31611),
            .I(N__31582));
    Span12Mux_v I__6917 (
            .O(N__31606),
            .I(N__31576));
    Span12Mux_v I__6916 (
            .O(N__31601),
            .I(N__31576));
    Span4Mux_h I__6915 (
            .O(N__31596),
            .I(N__31573));
    Span4Mux_h I__6914 (
            .O(N__31593),
            .I(N__31568));
    Span4Mux_h I__6913 (
            .O(N__31588),
            .I(N__31568));
    Span12Mux_v I__6912 (
            .O(N__31585),
            .I(N__31563));
    LocalMux I__6911 (
            .O(N__31582),
            .I(N__31563));
    InMux I__6910 (
            .O(N__31581),
            .I(N__31560));
    Odrv12 I__6909 (
            .O(N__31576),
            .I(M_this_spr_address_qZ0Z_5));
    Odrv4 I__6908 (
            .O(N__31573),
            .I(M_this_spr_address_qZ0Z_5));
    Odrv4 I__6907 (
            .O(N__31568),
            .I(M_this_spr_address_qZ0Z_5));
    Odrv12 I__6906 (
            .O(N__31563),
            .I(M_this_spr_address_qZ0Z_5));
    LocalMux I__6905 (
            .O(N__31560),
            .I(M_this_spr_address_qZ0Z_5));
    InMux I__6904 (
            .O(N__31549),
            .I(un1_M_this_spr_address_q_cry_4));
    CascadeMux I__6903 (
            .O(N__31546),
            .I(N__31540));
    CascadeMux I__6902 (
            .O(N__31545),
            .I(N__31535));
    CascadeMux I__6901 (
            .O(N__31544),
            .I(N__31530));
    CascadeMux I__6900 (
            .O(N__31543),
            .I(N__31527));
    InMux I__6899 (
            .O(N__31540),
            .I(N__31522));
    CascadeMux I__6898 (
            .O(N__31539),
            .I(N__31519));
    CascadeMux I__6897 (
            .O(N__31538),
            .I(N__31516));
    InMux I__6896 (
            .O(N__31535),
            .I(N__31511));
    CascadeMux I__6895 (
            .O(N__31534),
            .I(N__31508));
    CascadeMux I__6894 (
            .O(N__31533),
            .I(N__31505));
    InMux I__6893 (
            .O(N__31530),
            .I(N__31502));
    InMux I__6892 (
            .O(N__31527),
            .I(N__31499));
    CascadeMux I__6891 (
            .O(N__31526),
            .I(N__31496));
    CascadeMux I__6890 (
            .O(N__31525),
            .I(N__31493));
    LocalMux I__6889 (
            .O(N__31522),
            .I(N__31489));
    InMux I__6888 (
            .O(N__31519),
            .I(N__31486));
    InMux I__6887 (
            .O(N__31516),
            .I(N__31483));
    CascadeMux I__6886 (
            .O(N__31515),
            .I(N__31480));
    CascadeMux I__6885 (
            .O(N__31514),
            .I(N__31477));
    LocalMux I__6884 (
            .O(N__31511),
            .I(N__31472));
    InMux I__6883 (
            .O(N__31508),
            .I(N__31469));
    InMux I__6882 (
            .O(N__31505),
            .I(N__31466));
    LocalMux I__6881 (
            .O(N__31502),
            .I(N__31463));
    LocalMux I__6880 (
            .O(N__31499),
            .I(N__31460));
    InMux I__6879 (
            .O(N__31496),
            .I(N__31457));
    InMux I__6878 (
            .O(N__31493),
            .I(N__31454));
    CascadeMux I__6877 (
            .O(N__31492),
            .I(N__31451));
    Span4Mux_v I__6876 (
            .O(N__31489),
            .I(N__31444));
    LocalMux I__6875 (
            .O(N__31486),
            .I(N__31444));
    LocalMux I__6874 (
            .O(N__31483),
            .I(N__31444));
    InMux I__6873 (
            .O(N__31480),
            .I(N__31441));
    InMux I__6872 (
            .O(N__31477),
            .I(N__31438));
    CascadeMux I__6871 (
            .O(N__31476),
            .I(N__31435));
    CascadeMux I__6870 (
            .O(N__31475),
            .I(N__31432));
    Sp12to4 I__6869 (
            .O(N__31472),
            .I(N__31425));
    LocalMux I__6868 (
            .O(N__31469),
            .I(N__31425));
    LocalMux I__6867 (
            .O(N__31466),
            .I(N__31425));
    Span4Mux_v I__6866 (
            .O(N__31463),
            .I(N__31417));
    Span4Mux_h I__6865 (
            .O(N__31460),
            .I(N__31417));
    LocalMux I__6864 (
            .O(N__31457),
            .I(N__31417));
    LocalMux I__6863 (
            .O(N__31454),
            .I(N__31414));
    InMux I__6862 (
            .O(N__31451),
            .I(N__31411));
    Span4Mux_v I__6861 (
            .O(N__31444),
            .I(N__31404));
    LocalMux I__6860 (
            .O(N__31441),
            .I(N__31404));
    LocalMux I__6859 (
            .O(N__31438),
            .I(N__31404));
    InMux I__6858 (
            .O(N__31435),
            .I(N__31401));
    InMux I__6857 (
            .O(N__31432),
            .I(N__31398));
    Span12Mux_s6_v I__6856 (
            .O(N__31425),
            .I(N__31395));
    CascadeMux I__6855 (
            .O(N__31424),
            .I(N__31392));
    Span4Mux_v I__6854 (
            .O(N__31417),
            .I(N__31385));
    Span4Mux_h I__6853 (
            .O(N__31414),
            .I(N__31385));
    LocalMux I__6852 (
            .O(N__31411),
            .I(N__31385));
    Span4Mux_v I__6851 (
            .O(N__31404),
            .I(N__31378));
    LocalMux I__6850 (
            .O(N__31401),
            .I(N__31378));
    LocalMux I__6849 (
            .O(N__31398),
            .I(N__31378));
    Span12Mux_v I__6848 (
            .O(N__31395),
            .I(N__31375));
    InMux I__6847 (
            .O(N__31392),
            .I(N__31372));
    Span4Mux_v I__6846 (
            .O(N__31385),
            .I(N__31366));
    Span4Mux_v I__6845 (
            .O(N__31378),
            .I(N__31366));
    Span12Mux_h I__6844 (
            .O(N__31375),
            .I(N__31361));
    LocalMux I__6843 (
            .O(N__31372),
            .I(N__31361));
    InMux I__6842 (
            .O(N__31371),
            .I(N__31358));
    Odrv4 I__6841 (
            .O(N__31366),
            .I(M_this_spr_address_qZ0Z_6));
    Odrv12 I__6840 (
            .O(N__31361),
            .I(M_this_spr_address_qZ0Z_6));
    LocalMux I__6839 (
            .O(N__31358),
            .I(M_this_spr_address_qZ0Z_6));
    InMux I__6838 (
            .O(N__31351),
            .I(un1_M_this_spr_address_q_cry_5));
    CascadeMux I__6837 (
            .O(N__31348),
            .I(N__31344));
    CascadeMux I__6836 (
            .O(N__31347),
            .I(N__31341));
    InMux I__6835 (
            .O(N__31344),
            .I(N__31334));
    InMux I__6834 (
            .O(N__31341),
            .I(N__31331));
    CascadeMux I__6833 (
            .O(N__31340),
            .I(N__31328));
    CascadeMux I__6832 (
            .O(N__31339),
            .I(N__31325));
    CascadeMux I__6831 (
            .O(N__31338),
            .I(N__31320));
    CascadeMux I__6830 (
            .O(N__31337),
            .I(N__31317));
    LocalMux I__6829 (
            .O(N__31334),
            .I(N__31312));
    LocalMux I__6828 (
            .O(N__31331),
            .I(N__31309));
    InMux I__6827 (
            .O(N__31328),
            .I(N__31306));
    InMux I__6826 (
            .O(N__31325),
            .I(N__31303));
    CascadeMux I__6825 (
            .O(N__31324),
            .I(N__31300));
    CascadeMux I__6824 (
            .O(N__31323),
            .I(N__31297));
    InMux I__6823 (
            .O(N__31320),
            .I(N__31292));
    InMux I__6822 (
            .O(N__31317),
            .I(N__31289));
    CascadeMux I__6821 (
            .O(N__31316),
            .I(N__31286));
    CascadeMux I__6820 (
            .O(N__31315),
            .I(N__31283));
    Span4Mux_s2_v I__6819 (
            .O(N__31312),
            .I(N__31277));
    Span4Mux_h I__6818 (
            .O(N__31309),
            .I(N__31277));
    LocalMux I__6817 (
            .O(N__31306),
            .I(N__31274));
    LocalMux I__6816 (
            .O(N__31303),
            .I(N__31271));
    InMux I__6815 (
            .O(N__31300),
            .I(N__31268));
    InMux I__6814 (
            .O(N__31297),
            .I(N__31265));
    CascadeMux I__6813 (
            .O(N__31296),
            .I(N__31262));
    CascadeMux I__6812 (
            .O(N__31295),
            .I(N__31259));
    LocalMux I__6811 (
            .O(N__31292),
            .I(N__31255));
    LocalMux I__6810 (
            .O(N__31289),
            .I(N__31252));
    InMux I__6809 (
            .O(N__31286),
            .I(N__31249));
    InMux I__6808 (
            .O(N__31283),
            .I(N__31246));
    CascadeMux I__6807 (
            .O(N__31282),
            .I(N__31243));
    Span4Mux_v I__6806 (
            .O(N__31277),
            .I(N__31236));
    Span4Mux_v I__6805 (
            .O(N__31274),
            .I(N__31236));
    Span4Mux_v I__6804 (
            .O(N__31271),
            .I(N__31229));
    LocalMux I__6803 (
            .O(N__31268),
            .I(N__31229));
    LocalMux I__6802 (
            .O(N__31265),
            .I(N__31229));
    InMux I__6801 (
            .O(N__31262),
            .I(N__31226));
    InMux I__6800 (
            .O(N__31259),
            .I(N__31223));
    CascadeMux I__6799 (
            .O(N__31258),
            .I(N__31220));
    Span4Mux_v I__6798 (
            .O(N__31255),
            .I(N__31213));
    Span4Mux_h I__6797 (
            .O(N__31252),
            .I(N__31213));
    LocalMux I__6796 (
            .O(N__31249),
            .I(N__31213));
    LocalMux I__6795 (
            .O(N__31246),
            .I(N__31210));
    InMux I__6794 (
            .O(N__31243),
            .I(N__31207));
    CascadeMux I__6793 (
            .O(N__31242),
            .I(N__31204));
    CascadeMux I__6792 (
            .O(N__31241),
            .I(N__31201));
    Sp12to4 I__6791 (
            .O(N__31236),
            .I(N__31198));
    Span4Mux_v I__6790 (
            .O(N__31229),
            .I(N__31191));
    LocalMux I__6789 (
            .O(N__31226),
            .I(N__31191));
    LocalMux I__6788 (
            .O(N__31223),
            .I(N__31191));
    InMux I__6787 (
            .O(N__31220),
            .I(N__31188));
    Span4Mux_v I__6786 (
            .O(N__31213),
            .I(N__31181));
    Span4Mux_h I__6785 (
            .O(N__31210),
            .I(N__31181));
    LocalMux I__6784 (
            .O(N__31207),
            .I(N__31181));
    InMux I__6783 (
            .O(N__31204),
            .I(N__31178));
    InMux I__6782 (
            .O(N__31201),
            .I(N__31175));
    Span12Mux_h I__6781 (
            .O(N__31198),
            .I(N__31172));
    Span4Mux_v I__6780 (
            .O(N__31191),
            .I(N__31163));
    LocalMux I__6779 (
            .O(N__31188),
            .I(N__31163));
    Span4Mux_v I__6778 (
            .O(N__31181),
            .I(N__31163));
    LocalMux I__6777 (
            .O(N__31178),
            .I(N__31163));
    LocalMux I__6776 (
            .O(N__31175),
            .I(N__31160));
    Span12Mux_v I__6775 (
            .O(N__31172),
            .I(N__31156));
    Span4Mux_v I__6774 (
            .O(N__31163),
            .I(N__31151));
    Span4Mux_h I__6773 (
            .O(N__31160),
            .I(N__31151));
    InMux I__6772 (
            .O(N__31159),
            .I(N__31148));
    Odrv12 I__6771 (
            .O(N__31156),
            .I(M_this_spr_address_qZ0Z_7));
    Odrv4 I__6770 (
            .O(N__31151),
            .I(M_this_spr_address_qZ0Z_7));
    LocalMux I__6769 (
            .O(N__31148),
            .I(M_this_spr_address_qZ0Z_7));
    InMux I__6768 (
            .O(N__31141),
            .I(un1_M_this_spr_address_q_cry_6));
    InMux I__6767 (
            .O(N__31138),
            .I(N__31132));
    InMux I__6766 (
            .O(N__31137),
            .I(N__31132));
    LocalMux I__6765 (
            .O(N__31132),
            .I(\this_ppu.N_1176_1 ));
    InMux I__6764 (
            .O(N__31129),
            .I(N__31126));
    LocalMux I__6763 (
            .O(N__31126),
            .I(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_3 ));
    CascadeMux I__6762 (
            .O(N__31123),
            .I(N__31120));
    InMux I__6761 (
            .O(N__31120),
            .I(N__31117));
    LocalMux I__6760 (
            .O(N__31117),
            .I(N__31114));
    Odrv4 I__6759 (
            .O(N__31114),
            .I(\this_ppu.N_893 ));
    CascadeMux I__6758 (
            .O(N__31111),
            .I(N__31108));
    InMux I__6757 (
            .O(N__31108),
            .I(N__31105));
    LocalMux I__6756 (
            .O(N__31105),
            .I(\this_ppu.N_969 ));
    CascadeMux I__6755 (
            .O(N__31102),
            .I(un1_M_this_state_q_11_0_0_cascade_));
    CascadeMux I__6754 (
            .O(N__31099),
            .I(\this_ppu.un1_M_this_state_q_11_0_0Z0Z_0_cascade_ ));
    InMux I__6753 (
            .O(N__31096),
            .I(N__31093));
    LocalMux I__6752 (
            .O(N__31093),
            .I(\this_ppu.un1_M_this_state_q_11_0_0Z0Z_1 ));
    CascadeMux I__6751 (
            .O(N__31090),
            .I(N__31085));
    InMux I__6750 (
            .O(N__31089),
            .I(N__31080));
    InMux I__6749 (
            .O(N__31088),
            .I(N__31080));
    InMux I__6748 (
            .O(N__31085),
            .I(N__31076));
    LocalMux I__6747 (
            .O(N__31080),
            .I(N__31072));
    InMux I__6746 (
            .O(N__31079),
            .I(N__31069));
    LocalMux I__6745 (
            .O(N__31076),
            .I(N__31060));
    CascadeMux I__6744 (
            .O(N__31075),
            .I(N__31056));
    Span4Mux_v I__6743 (
            .O(N__31072),
            .I(N__31049));
    LocalMux I__6742 (
            .O(N__31069),
            .I(N__31049));
    InMux I__6741 (
            .O(N__31068),
            .I(N__31040));
    InMux I__6740 (
            .O(N__31067),
            .I(N__31040));
    InMux I__6739 (
            .O(N__31066),
            .I(N__31040));
    InMux I__6738 (
            .O(N__31065),
            .I(N__31040));
    InMux I__6737 (
            .O(N__31064),
            .I(N__31035));
    InMux I__6736 (
            .O(N__31063),
            .I(N__31035));
    Span4Mux_v I__6735 (
            .O(N__31060),
            .I(N__31031));
    InMux I__6734 (
            .O(N__31059),
            .I(N__31028));
    InMux I__6733 (
            .O(N__31056),
            .I(N__31025));
    InMux I__6732 (
            .O(N__31055),
            .I(N__31020));
    InMux I__6731 (
            .O(N__31054),
            .I(N__31020));
    Span4Mux_h I__6730 (
            .O(N__31049),
            .I(N__31017));
    LocalMux I__6729 (
            .O(N__31040),
            .I(N__31012));
    LocalMux I__6728 (
            .O(N__31035),
            .I(N__31012));
    InMux I__6727 (
            .O(N__31034),
            .I(N__31009));
    Odrv4 I__6726 (
            .O(N__31031),
            .I(\this_ppu.N_430_1_0 ));
    LocalMux I__6725 (
            .O(N__31028),
            .I(\this_ppu.N_430_1_0 ));
    LocalMux I__6724 (
            .O(N__31025),
            .I(\this_ppu.N_430_1_0 ));
    LocalMux I__6723 (
            .O(N__31020),
            .I(\this_ppu.N_430_1_0 ));
    Odrv4 I__6722 (
            .O(N__31017),
            .I(\this_ppu.N_430_1_0 ));
    Odrv12 I__6721 (
            .O(N__31012),
            .I(\this_ppu.N_430_1_0 ));
    LocalMux I__6720 (
            .O(N__31009),
            .I(\this_ppu.N_430_1_0 ));
    CascadeMux I__6719 (
            .O(N__30994),
            .I(N__30991));
    InMux I__6718 (
            .O(N__30991),
            .I(N__30987));
    InMux I__6717 (
            .O(N__30990),
            .I(N__30984));
    LocalMux I__6716 (
            .O(N__30987),
            .I(N__30981));
    LocalMux I__6715 (
            .O(N__30984),
            .I(N__30978));
    Odrv4 I__6714 (
            .O(N__30981),
            .I(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_2 ));
    Odrv4 I__6713 (
            .O(N__30978),
            .I(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_2 ));
    CascadeMux I__6712 (
            .O(N__30973),
            .I(\this_ppu.N_1158_cascade_ ));
    InMux I__6711 (
            .O(N__30970),
            .I(N__30966));
    InMux I__6710 (
            .O(N__30969),
            .I(N__30963));
    LocalMux I__6709 (
            .O(N__30966),
            .I(N__30960));
    LocalMux I__6708 (
            .O(N__30963),
            .I(\this_ppu.N_1263 ));
    Odrv4 I__6707 (
            .O(N__30960),
            .I(\this_ppu.N_1263 ));
    CascadeMux I__6706 (
            .O(N__30955),
            .I(N__30952));
    InMux I__6705 (
            .O(N__30952),
            .I(N__30949));
    LocalMux I__6704 (
            .O(N__30949),
            .I(N__30946));
    Odrv4 I__6703 (
            .O(N__30946),
            .I(\this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1Z0Z_0 ));
    InMux I__6702 (
            .O(N__30943),
            .I(N__30940));
    LocalMux I__6701 (
            .O(N__30940),
            .I(\this_ppu.M_this_state_q_srsts_0_0_0_tz_0_0 ));
    InMux I__6700 (
            .O(N__30937),
            .I(N__30933));
    InMux I__6699 (
            .O(N__30936),
            .I(N__30930));
    LocalMux I__6698 (
            .O(N__30933),
            .I(N__30925));
    LocalMux I__6697 (
            .O(N__30930),
            .I(N__30922));
    InMux I__6696 (
            .O(N__30929),
            .I(N__30919));
    InMux I__6695 (
            .O(N__30928),
            .I(N__30915));
    Span4Mux_v I__6694 (
            .O(N__30925),
            .I(N__30910));
    Span4Mux_v I__6693 (
            .O(N__30922),
            .I(N__30910));
    LocalMux I__6692 (
            .O(N__30919),
            .I(N__30907));
    InMux I__6691 (
            .O(N__30918),
            .I(N__30904));
    LocalMux I__6690 (
            .O(N__30915),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__6689 (
            .O(N__30910),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__6688 (
            .O(N__30907),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__6687 (
            .O(N__30904),
            .I(M_this_state_qZ0Z_8));
    InMux I__6686 (
            .O(N__30895),
            .I(N__30892));
    LocalMux I__6685 (
            .O(N__30892),
            .I(N__30889));
    Span4Mux_h I__6684 (
            .O(N__30889),
            .I(N__30884));
    InMux I__6683 (
            .O(N__30888),
            .I(N__30881));
    InMux I__6682 (
            .O(N__30887),
            .I(N__30878));
    Odrv4 I__6681 (
            .O(N__30884),
            .I(N_815_0));
    LocalMux I__6680 (
            .O(N__30881),
            .I(N_815_0));
    LocalMux I__6679 (
            .O(N__30878),
            .I(N_815_0));
    IoInMux I__6678 (
            .O(N__30871),
            .I(N__30868));
    LocalMux I__6677 (
            .O(N__30868),
            .I(N__30865));
    IoSpan4Mux I__6676 (
            .O(N__30865),
            .I(N__30862));
    Span4Mux_s3_h I__6675 (
            .O(N__30862),
            .I(N__30859));
    Sp12to4 I__6674 (
            .O(N__30859),
            .I(N__30856));
    Span12Mux_s11_h I__6673 (
            .O(N__30856),
            .I(N__30853));
    Span12Mux_v I__6672 (
            .O(N__30853),
            .I(N__30850));
    Odrv12 I__6671 (
            .O(N__30850),
            .I(led_c_7));
    CascadeMux I__6670 (
            .O(N__30847),
            .I(N__30844));
    InMux I__6669 (
            .O(N__30844),
            .I(N__30841));
    LocalMux I__6668 (
            .O(N__30841),
            .I(\this_ppu.N_807_0 ));
    InMux I__6667 (
            .O(N__30838),
            .I(N__30828));
    InMux I__6666 (
            .O(N__30837),
            .I(N__30828));
    InMux I__6665 (
            .O(N__30836),
            .I(N__30825));
    InMux I__6664 (
            .O(N__30835),
            .I(N__30822));
    InMux I__6663 (
            .O(N__30834),
            .I(N__30819));
    InMux I__6662 (
            .O(N__30833),
            .I(N__30816));
    LocalMux I__6661 (
            .O(N__30828),
            .I(M_this_state_qZ0Z_16));
    LocalMux I__6660 (
            .O(N__30825),
            .I(M_this_state_qZ0Z_16));
    LocalMux I__6659 (
            .O(N__30822),
            .I(M_this_state_qZ0Z_16));
    LocalMux I__6658 (
            .O(N__30819),
            .I(M_this_state_qZ0Z_16));
    LocalMux I__6657 (
            .O(N__30816),
            .I(M_this_state_qZ0Z_16));
    InMux I__6656 (
            .O(N__30805),
            .I(N__30802));
    LocalMux I__6655 (
            .O(N__30802),
            .I(N__30799));
    Odrv12 I__6654 (
            .O(N__30799),
            .I(N_1415));
    CascadeMux I__6653 (
            .O(N__30796),
            .I(N_1415_cascade_));
    InMux I__6652 (
            .O(N__30793),
            .I(N__30785));
    InMux I__6651 (
            .O(N__30792),
            .I(N__30785));
    InMux I__6650 (
            .O(N__30791),
            .I(N__30780));
    InMux I__6649 (
            .O(N__30790),
            .I(N__30780));
    LocalMux I__6648 (
            .O(N__30785),
            .I(\this_ppu.N_1278 ));
    LocalMux I__6647 (
            .O(N__30780),
            .I(\this_ppu.N_1278 ));
    InMux I__6646 (
            .O(N__30775),
            .I(N__30772));
    LocalMux I__6645 (
            .O(N__30772),
            .I(\this_ppu.N_1166 ));
    CascadeMux I__6644 (
            .O(N__30769),
            .I(\this_ppu.N_1263_cascade_ ));
    InMux I__6643 (
            .O(N__30766),
            .I(N__30763));
    LocalMux I__6642 (
            .O(N__30763),
            .I(N__30759));
    InMux I__6641 (
            .O(N__30762),
            .I(N__30756));
    Span4Mux_h I__6640 (
            .O(N__30759),
            .I(N__30752));
    LocalMux I__6639 (
            .O(N__30756),
            .I(N__30749));
    InMux I__6638 (
            .O(N__30755),
            .I(N__30746));
    Span4Mux_v I__6637 (
            .O(N__30752),
            .I(N__30743));
    Span4Mux_v I__6636 (
            .O(N__30749),
            .I(N__30740));
    LocalMux I__6635 (
            .O(N__30746),
            .I(N__30737));
    Odrv4 I__6634 (
            .O(N__30743),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    Odrv4 I__6633 (
            .O(N__30740),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    Odrv12 I__6632 (
            .O(N__30737),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    InMux I__6631 (
            .O(N__30730),
            .I(N__30727));
    LocalMux I__6630 (
            .O(N__30727),
            .I(N__30722));
    InMux I__6629 (
            .O(N__30726),
            .I(N__30719));
    InMux I__6628 (
            .O(N__30725),
            .I(N__30716));
    Span4Mux_v I__6627 (
            .O(N__30722),
            .I(N__30711));
    LocalMux I__6626 (
            .O(N__30719),
            .I(N__30711));
    LocalMux I__6625 (
            .O(N__30716),
            .I(N__30708));
    Span4Mux_v I__6624 (
            .O(N__30711),
            .I(N__30705));
    Odrv12 I__6623 (
            .O(N__30708),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    Odrv4 I__6622 (
            .O(N__30705),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    InMux I__6621 (
            .O(N__30700),
            .I(N__30694));
    InMux I__6620 (
            .O(N__30699),
            .I(N__30694));
    LocalMux I__6619 (
            .O(N__30694),
            .I(N__30689));
    InMux I__6618 (
            .O(N__30693),
            .I(N__30680));
    InMux I__6617 (
            .O(N__30692),
            .I(N__30677));
    Span4Mux_v I__6616 (
            .O(N__30689),
            .I(N__30674));
    InMux I__6615 (
            .O(N__30688),
            .I(N__30671));
    InMux I__6614 (
            .O(N__30687),
            .I(N__30664));
    InMux I__6613 (
            .O(N__30686),
            .I(N__30664));
    InMux I__6612 (
            .O(N__30685),
            .I(N__30661));
    InMux I__6611 (
            .O(N__30684),
            .I(N__30656));
    InMux I__6610 (
            .O(N__30683),
            .I(N__30656));
    LocalMux I__6609 (
            .O(N__30680),
            .I(N__30653));
    LocalMux I__6608 (
            .O(N__30677),
            .I(N__30648));
    Span4Mux_h I__6607 (
            .O(N__30674),
            .I(N__30645));
    LocalMux I__6606 (
            .O(N__30671),
            .I(N__30642));
    InMux I__6605 (
            .O(N__30670),
            .I(N__30639));
    InMux I__6604 (
            .O(N__30669),
            .I(N__30634));
    LocalMux I__6603 (
            .O(N__30664),
            .I(N__30627));
    LocalMux I__6602 (
            .O(N__30661),
            .I(N__30627));
    LocalMux I__6601 (
            .O(N__30656),
            .I(N__30627));
    Span4Mux_v I__6600 (
            .O(N__30653),
            .I(N__30624));
    InMux I__6599 (
            .O(N__30652),
            .I(N__30619));
    InMux I__6598 (
            .O(N__30651),
            .I(N__30619));
    Span4Mux_v I__6597 (
            .O(N__30648),
            .I(N__30610));
    Span4Mux_h I__6596 (
            .O(N__30645),
            .I(N__30610));
    Span4Mux_v I__6595 (
            .O(N__30642),
            .I(N__30610));
    LocalMux I__6594 (
            .O(N__30639),
            .I(N__30610));
    InMux I__6593 (
            .O(N__30638),
            .I(N__30605));
    InMux I__6592 (
            .O(N__30637),
            .I(N__30605));
    LocalMux I__6591 (
            .O(N__30634),
            .I(N__30600));
    Span4Mux_h I__6590 (
            .O(N__30627),
            .I(N__30600));
    Odrv4 I__6589 (
            .O(N__30624),
            .I(this_vga_signals_M_vcounter_q_8));
    LocalMux I__6588 (
            .O(N__30619),
            .I(this_vga_signals_M_vcounter_q_8));
    Odrv4 I__6587 (
            .O(N__30610),
            .I(this_vga_signals_M_vcounter_q_8));
    LocalMux I__6586 (
            .O(N__30605),
            .I(this_vga_signals_M_vcounter_q_8));
    Odrv4 I__6585 (
            .O(N__30600),
            .I(this_vga_signals_M_vcounter_q_8));
    InMux I__6584 (
            .O(N__30589),
            .I(N__30585));
    InMux I__6583 (
            .O(N__30588),
            .I(N__30582));
    LocalMux I__6582 (
            .O(N__30585),
            .I(N__30578));
    LocalMux I__6581 (
            .O(N__30582),
            .I(N__30575));
    InMux I__6580 (
            .O(N__30581),
            .I(N__30572));
    Span4Mux_v I__6579 (
            .O(N__30578),
            .I(N__30568));
    Span4Mux_h I__6578 (
            .O(N__30575),
            .I(N__30562));
    LocalMux I__6577 (
            .O(N__30572),
            .I(N__30562));
    InMux I__6576 (
            .O(N__30571),
            .I(N__30559));
    Span4Mux_h I__6575 (
            .O(N__30568),
            .I(N__30556));
    InMux I__6574 (
            .O(N__30567),
            .I(N__30553));
    Span4Mux_v I__6573 (
            .O(N__30562),
            .I(N__30548));
    LocalMux I__6572 (
            .O(N__30559),
            .I(N__30548));
    Odrv4 I__6571 (
            .O(N__30556),
            .I(N_1001_0));
    LocalMux I__6570 (
            .O(N__30553),
            .I(N_1001_0));
    Odrv4 I__6569 (
            .O(N__30548),
            .I(N_1001_0));
    InMux I__6568 (
            .O(N__30541),
            .I(N__30536));
    InMux I__6567 (
            .O(N__30540),
            .I(N__30527));
    InMux I__6566 (
            .O(N__30539),
            .I(N__30527));
    LocalMux I__6565 (
            .O(N__30536),
            .I(N__30524));
    InMux I__6564 (
            .O(N__30535),
            .I(N__30521));
    InMux I__6563 (
            .O(N__30534),
            .I(N__30517));
    InMux I__6562 (
            .O(N__30533),
            .I(N__30514));
    InMux I__6561 (
            .O(N__30532),
            .I(N__30511));
    LocalMux I__6560 (
            .O(N__30527),
            .I(N__30508));
    Span4Mux_v I__6559 (
            .O(N__30524),
            .I(N__30503));
    LocalMux I__6558 (
            .O(N__30521),
            .I(N__30503));
    InMux I__6557 (
            .O(N__30520),
            .I(N__30498));
    LocalMux I__6556 (
            .O(N__30517),
            .I(N__30487));
    LocalMux I__6555 (
            .O(N__30514),
            .I(N__30487));
    LocalMux I__6554 (
            .O(N__30511),
            .I(N__30487));
    Span4Mux_h I__6553 (
            .O(N__30508),
            .I(N__30487));
    Span4Mux_h I__6552 (
            .O(N__30503),
            .I(N__30487));
    InMux I__6551 (
            .O(N__30502),
            .I(N__30482));
    InMux I__6550 (
            .O(N__30501),
            .I(N__30482));
    LocalMux I__6549 (
            .O(N__30498),
            .I(N_814_0));
    Odrv4 I__6548 (
            .O(N__30487),
            .I(N_814_0));
    LocalMux I__6547 (
            .O(N__30482),
            .I(N_814_0));
    CascadeMux I__6546 (
            .O(N__30475),
            .I(N_1001_0_cascade_));
    CascadeMux I__6545 (
            .O(N__30472),
            .I(N__30469));
    InMux I__6544 (
            .O(N__30469),
            .I(N__30463));
    InMux I__6543 (
            .O(N__30468),
            .I(N__30460));
    InMux I__6542 (
            .O(N__30467),
            .I(N__30448));
    InMux I__6541 (
            .O(N__30466),
            .I(N__30445));
    LocalMux I__6540 (
            .O(N__30463),
            .I(N__30442));
    LocalMux I__6539 (
            .O(N__30460),
            .I(N__30439));
    InMux I__6538 (
            .O(N__30459),
            .I(N__30436));
    InMux I__6537 (
            .O(N__30458),
            .I(N__30433));
    InMux I__6536 (
            .O(N__30457),
            .I(N__30430));
    InMux I__6535 (
            .O(N__30456),
            .I(N__30425));
    InMux I__6534 (
            .O(N__30455),
            .I(N__30422));
    InMux I__6533 (
            .O(N__30454),
            .I(N__30415));
    InMux I__6532 (
            .O(N__30453),
            .I(N__30415));
    InMux I__6531 (
            .O(N__30452),
            .I(N__30412));
    CascadeMux I__6530 (
            .O(N__30451),
            .I(N__30409));
    LocalMux I__6529 (
            .O(N__30448),
            .I(N__30406));
    LocalMux I__6528 (
            .O(N__30445),
            .I(N__30403));
    Span4Mux_h I__6527 (
            .O(N__30442),
            .I(N__30398));
    Span4Mux_v I__6526 (
            .O(N__30439),
            .I(N__30398));
    LocalMux I__6525 (
            .O(N__30436),
            .I(N__30393));
    LocalMux I__6524 (
            .O(N__30433),
            .I(N__30393));
    LocalMux I__6523 (
            .O(N__30430),
            .I(N__30390));
    InMux I__6522 (
            .O(N__30429),
            .I(N__30385));
    InMux I__6521 (
            .O(N__30428),
            .I(N__30385));
    LocalMux I__6520 (
            .O(N__30425),
            .I(N__30380));
    LocalMux I__6519 (
            .O(N__30422),
            .I(N__30380));
    InMux I__6518 (
            .O(N__30421),
            .I(N__30377));
    InMux I__6517 (
            .O(N__30420),
            .I(N__30374));
    LocalMux I__6516 (
            .O(N__30415),
            .I(N__30371));
    LocalMux I__6515 (
            .O(N__30412),
            .I(N__30368));
    InMux I__6514 (
            .O(N__30409),
            .I(N__30365));
    Span4Mux_v I__6513 (
            .O(N__30406),
            .I(N__30356));
    Span4Mux_v I__6512 (
            .O(N__30403),
            .I(N__30356));
    Span4Mux_h I__6511 (
            .O(N__30398),
            .I(N__30356));
    Span4Mux_v I__6510 (
            .O(N__30393),
            .I(N__30356));
    Span4Mux_v I__6509 (
            .O(N__30390),
            .I(N__30349));
    LocalMux I__6508 (
            .O(N__30385),
            .I(N__30349));
    Span4Mux_h I__6507 (
            .O(N__30380),
            .I(N__30349));
    LocalMux I__6506 (
            .O(N__30377),
            .I(N__30346));
    LocalMux I__6505 (
            .O(N__30374),
            .I(N__30343));
    Odrv4 I__6504 (
            .O(N__30371),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv12 I__6503 (
            .O(N__30368),
            .I(this_vga_signals_M_vcounter_q_9));
    LocalMux I__6502 (
            .O(N__30365),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv4 I__6501 (
            .O(N__30356),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv4 I__6500 (
            .O(N__30349),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv12 I__6499 (
            .O(N__30346),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv4 I__6498 (
            .O(N__30343),
            .I(this_vga_signals_M_vcounter_q_9));
    InMux I__6497 (
            .O(N__30328),
            .I(N__30325));
    LocalMux I__6496 (
            .O(N__30325),
            .I(N__30322));
    Odrv12 I__6495 (
            .O(N__30322),
            .I(\this_vga_signals.g4 ));
    CascadeMux I__6494 (
            .O(N__30319),
            .I(\this_ppu.N_1278_cascade_ ));
    InMux I__6493 (
            .O(N__30316),
            .I(N__30310));
    InMux I__6492 (
            .O(N__30315),
            .I(N__30310));
    LocalMux I__6491 (
            .O(N__30310),
            .I(N__30307));
    Span4Mux_h I__6490 (
            .O(N__30307),
            .I(N__30304));
    Odrv4 I__6489 (
            .O(N__30304),
            .I(\this_ppu.N_767_0 ));
    InMux I__6488 (
            .O(N__30301),
            .I(N__30298));
    LocalMux I__6487 (
            .O(N__30298),
            .I(N__30293));
    InMux I__6486 (
            .O(N__30297),
            .I(N__30288));
    InMux I__6485 (
            .O(N__30296),
            .I(N__30288));
    Odrv4 I__6484 (
            .O(N__30293),
            .I(\this_ppu.N_1425 ));
    LocalMux I__6483 (
            .O(N__30288),
            .I(\this_ppu.N_1425 ));
    CascadeMux I__6482 (
            .O(N__30283),
            .I(\this_ppu.N_1149_cascade_ ));
    CascadeMux I__6481 (
            .O(N__30280),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_3_cascade_ ));
    CascadeMux I__6480 (
            .O(N__30277),
            .I(\this_vga_signals.g1_0_0_0_cascade_ ));
    InMux I__6479 (
            .O(N__30274),
            .I(N__30271));
    LocalMux I__6478 (
            .O(N__30271),
            .I(N__30268));
    Span4Mux_v I__6477 (
            .O(N__30268),
            .I(N__30265));
    Sp12to4 I__6476 (
            .O(N__30265),
            .I(N__30262));
    Odrv12 I__6475 (
            .O(N__30262),
            .I(\this_vga_signals.SUM_2_i_i_1_0_3 ));
    InMux I__6474 (
            .O(N__30259),
            .I(N__30256));
    LocalMux I__6473 (
            .O(N__30256),
            .I(N__30253));
    Odrv4 I__6472 (
            .O(N__30253),
            .I(\this_vga_signals.N_5_0_0 ));
    InMux I__6471 (
            .O(N__30250),
            .I(N__30247));
    LocalMux I__6470 (
            .O(N__30247),
            .I(N__30244));
    Odrv4 I__6469 (
            .O(N__30244),
            .I(\this_vga_signals.g1_0_1 ));
    InMux I__6468 (
            .O(N__30241),
            .I(N__30235));
    InMux I__6467 (
            .O(N__30240),
            .I(N__30235));
    LocalMux I__6466 (
            .O(N__30235),
            .I(N__30232));
    Odrv4 I__6465 (
            .O(N__30232),
            .I(\this_vga_signals.N_39_0_0 ));
    CascadeMux I__6464 (
            .O(N__30229),
            .I(\this_vga_signals.g1_3_0_0_cascade_ ));
    InMux I__6463 (
            .O(N__30226),
            .I(N__30223));
    LocalMux I__6462 (
            .O(N__30223),
            .I(\this_vga_signals.N_4_1 ));
    CascadeMux I__6461 (
            .O(N__30220),
            .I(\this_vga_signals.g3_cascade_ ));
    InMux I__6460 (
            .O(N__30217),
            .I(N__30214));
    LocalMux I__6459 (
            .O(N__30214),
            .I(\this_vga_signals.N_5_1 ));
    InMux I__6458 (
            .O(N__30211),
            .I(N__30208));
    LocalMux I__6457 (
            .O(N__30208),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_0_0_1 ));
    InMux I__6456 (
            .O(N__30205),
            .I(N__30202));
    LocalMux I__6455 (
            .O(N__30202),
            .I(N__30199));
    Odrv4 I__6454 (
            .O(N__30199),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    InMux I__6453 (
            .O(N__30196),
            .I(N__30193));
    LocalMux I__6452 (
            .O(N__30193),
            .I(N__30190));
    Odrv4 I__6451 (
            .O(N__30190),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_0_0_1 ));
    InMux I__6450 (
            .O(N__30187),
            .I(N__30183));
    CascadeMux I__6449 (
            .O(N__30186),
            .I(N__30180));
    LocalMux I__6448 (
            .O(N__30183),
            .I(N__30177));
    InMux I__6447 (
            .O(N__30180),
            .I(N__30174));
    Span4Mux_v I__6446 (
            .O(N__30177),
            .I(N__30168));
    LocalMux I__6445 (
            .O(N__30174),
            .I(N__30168));
    InMux I__6444 (
            .O(N__30173),
            .I(N__30165));
    Span4Mux_h I__6443 (
            .O(N__30168),
            .I(N__30162));
    LocalMux I__6442 (
            .O(N__30165),
            .I(\this_vga_signals.N_1264 ));
    Odrv4 I__6441 (
            .O(N__30162),
            .I(\this_vga_signals.N_1264 ));
    InMux I__6440 (
            .O(N__30157),
            .I(N__30153));
    InMux I__6439 (
            .O(N__30156),
            .I(N__30150));
    LocalMux I__6438 (
            .O(N__30153),
            .I(N__30147));
    LocalMux I__6437 (
            .O(N__30150),
            .I(N__30144));
    Span4Mux_v I__6436 (
            .O(N__30147),
            .I(N__30141));
    Span4Mux_h I__6435 (
            .O(N__30144),
            .I(N__30138));
    Odrv4 I__6434 (
            .O(N__30141),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    Odrv4 I__6433 (
            .O(N__30138),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    CascadeMux I__6432 (
            .O(N__30133),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_x1_cascade_ ));
    InMux I__6431 (
            .O(N__30130),
            .I(N__30127));
    LocalMux I__6430 (
            .O(N__30127),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_x0 ));
    InMux I__6429 (
            .O(N__30124),
            .I(N__30121));
    LocalMux I__6428 (
            .O(N__30121),
            .I(N__30118));
    Span4Mux_h I__6427 (
            .O(N__30118),
            .I(N__30115));
    Odrv4 I__6426 (
            .O(N__30115),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1 ));
    InMux I__6425 (
            .O(N__30112),
            .I(N__30109));
    LocalMux I__6424 (
            .O(N__30109),
            .I(N__30104));
    InMux I__6423 (
            .O(N__30108),
            .I(N__30098));
    InMux I__6422 (
            .O(N__30107),
            .I(N__30098));
    Span4Mux_v I__6421 (
            .O(N__30104),
            .I(N__30095));
    InMux I__6420 (
            .O(N__30103),
            .I(N__30092));
    LocalMux I__6419 (
            .O(N__30098),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__6418 (
            .O(N__30095),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__6417 (
            .O(N__30092),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    CascadeMux I__6416 (
            .O(N__30085),
            .I(\this_vga_signals.mult1_un47_sum_c2_0_cascade_ ));
    CascadeMux I__6415 (
            .O(N__30082),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ));
    InMux I__6414 (
            .O(N__30079),
            .I(N__30076));
    LocalMux I__6413 (
            .O(N__30076),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    InMux I__6412 (
            .O(N__30073),
            .I(N__30069));
    InMux I__6411 (
            .O(N__30072),
            .I(N__30066));
    LocalMux I__6410 (
            .O(N__30069),
            .I(N__30063));
    LocalMux I__6409 (
            .O(N__30066),
            .I(N__30060));
    Span4Mux_h I__6408 (
            .O(N__30063),
            .I(N__30057));
    Odrv4 I__6407 (
            .O(N__30060),
            .I(\this_vga_signals.g1_0 ));
    Odrv4 I__6406 (
            .O(N__30057),
            .I(\this_vga_signals.g1_0 ));
    CascadeMux I__6405 (
            .O(N__30052),
            .I(N__30049));
    InMux I__6404 (
            .O(N__30049),
            .I(N__30046));
    LocalMux I__6403 (
            .O(N__30046),
            .I(N__30043));
    Span4Mux_h I__6402 (
            .O(N__30043),
            .I(N__30040));
    Odrv4 I__6401 (
            .O(N__30040),
            .I(\this_vga_signals.g0_0_1 ));
    InMux I__6400 (
            .O(N__30037),
            .I(N__30034));
    LocalMux I__6399 (
            .O(N__30034),
            .I(\this_vga_signals.g0_3_0 ));
    InMux I__6398 (
            .O(N__30031),
            .I(N__30025));
    InMux I__6397 (
            .O(N__30030),
            .I(N__30020));
    InMux I__6396 (
            .O(N__30029),
            .I(N__30020));
    InMux I__6395 (
            .O(N__30028),
            .I(N__30013));
    LocalMux I__6394 (
            .O(N__30025),
            .I(N__30008));
    LocalMux I__6393 (
            .O(N__30020),
            .I(N__30008));
    InMux I__6392 (
            .O(N__30019),
            .I(N__30003));
    InMux I__6391 (
            .O(N__30018),
            .I(N__30003));
    InMux I__6390 (
            .O(N__30017),
            .I(N__29998));
    InMux I__6389 (
            .O(N__30016),
            .I(N__29998));
    LocalMux I__6388 (
            .O(N__30013),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    Odrv4 I__6387 (
            .O(N__30008),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    LocalMux I__6386 (
            .O(N__30003),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    LocalMux I__6385 (
            .O(N__29998),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    InMux I__6384 (
            .O(N__29989),
            .I(N__29984));
    CascadeMux I__6383 (
            .O(N__29988),
            .I(N__29975));
    InMux I__6382 (
            .O(N__29987),
            .I(N__29972));
    LocalMux I__6381 (
            .O(N__29984),
            .I(N__29969));
    InMux I__6380 (
            .O(N__29983),
            .I(N__29964));
    InMux I__6379 (
            .O(N__29982),
            .I(N__29964));
    InMux I__6378 (
            .O(N__29981),
            .I(N__29959));
    InMux I__6377 (
            .O(N__29980),
            .I(N__29959));
    InMux I__6376 (
            .O(N__29979),
            .I(N__29954));
    InMux I__6375 (
            .O(N__29978),
            .I(N__29954));
    InMux I__6374 (
            .O(N__29975),
            .I(N__29951));
    LocalMux I__6373 (
            .O(N__29972),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    Odrv4 I__6372 (
            .O(N__29969),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    LocalMux I__6371 (
            .O(N__29964),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    LocalMux I__6370 (
            .O(N__29959),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    LocalMux I__6369 (
            .O(N__29954),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    LocalMux I__6368 (
            .O(N__29951),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    InMux I__6367 (
            .O(N__29938),
            .I(N__29934));
    CascadeMux I__6366 (
            .O(N__29937),
            .I(N__29931));
    LocalMux I__6365 (
            .O(N__29934),
            .I(N__29926));
    InMux I__6364 (
            .O(N__29931),
            .I(N__29923));
    CascadeMux I__6363 (
            .O(N__29930),
            .I(N__29920));
    InMux I__6362 (
            .O(N__29929),
            .I(N__29917));
    Span4Mux_v I__6361 (
            .O(N__29926),
            .I(N__29912));
    LocalMux I__6360 (
            .O(N__29923),
            .I(N__29912));
    InMux I__6359 (
            .O(N__29920),
            .I(N__29909));
    LocalMux I__6358 (
            .O(N__29917),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    Odrv4 I__6357 (
            .O(N__29912),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__6356 (
            .O(N__29909),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    CascadeMux I__6355 (
            .O(N__29902),
            .I(N__29899));
    InMux I__6354 (
            .O(N__29899),
            .I(N__29896));
    LocalMux I__6353 (
            .O(N__29896),
            .I(N__29893));
    Span4Mux_h I__6352 (
            .O(N__29893),
            .I(N__29890));
    Odrv4 I__6351 (
            .O(N__29890),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_4_1_0 ));
    InMux I__6350 (
            .O(N__29887),
            .I(N__29881));
    InMux I__6349 (
            .O(N__29886),
            .I(N__29881));
    LocalMux I__6348 (
            .O(N__29881),
            .I(N__29877));
    InMux I__6347 (
            .O(N__29880),
            .I(N__29873));
    Span4Mux_h I__6346 (
            .O(N__29877),
            .I(N__29869));
    InMux I__6345 (
            .O(N__29876),
            .I(N__29866));
    LocalMux I__6344 (
            .O(N__29873),
            .I(N__29863));
    InMux I__6343 (
            .O(N__29872),
            .I(N__29860));
    Odrv4 I__6342 (
            .O(N__29869),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__6341 (
            .O(N__29866),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    Odrv12 I__6340 (
            .O(N__29863),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__6339 (
            .O(N__29860),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    InMux I__6338 (
            .O(N__29851),
            .I(N__29844));
    InMux I__6337 (
            .O(N__29850),
            .I(N__29844));
    CascadeMux I__6336 (
            .O(N__29849),
            .I(N__29839));
    LocalMux I__6335 (
            .O(N__29844),
            .I(N__29835));
    InMux I__6334 (
            .O(N__29843),
            .I(N__29832));
    InMux I__6333 (
            .O(N__29842),
            .I(N__29828));
    InMux I__6332 (
            .O(N__29839),
            .I(N__29823));
    InMux I__6331 (
            .O(N__29838),
            .I(N__29823));
    Span4Mux_v I__6330 (
            .O(N__29835),
            .I(N__29818));
    LocalMux I__6329 (
            .O(N__29832),
            .I(N__29818));
    InMux I__6328 (
            .O(N__29831),
            .I(N__29815));
    LocalMux I__6327 (
            .O(N__29828),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__6326 (
            .O(N__29823),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    Odrv4 I__6325 (
            .O(N__29818),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__6324 (
            .O(N__29815),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    CascadeMux I__6323 (
            .O(N__29806),
            .I(\this_vga_signals.mult1_un47_sum_3_3_cascade_ ));
    InMux I__6322 (
            .O(N__29803),
            .I(N__29800));
    LocalMux I__6321 (
            .O(N__29800),
            .I(N__29797));
    Span4Mux_h I__6320 (
            .O(N__29797),
            .I(N__29794));
    Odrv4 I__6319 (
            .O(N__29794),
            .I(\this_vga_signals.mult1_un54_sum_2_0_3 ));
    InMux I__6318 (
            .O(N__29791),
            .I(N__29788));
    LocalMux I__6317 (
            .O(N__29788),
            .I(N__29785));
    Span12Mux_v I__6316 (
            .O(N__29785),
            .I(N__29782));
    Span12Mux_h I__6315 (
            .O(N__29782),
            .I(N__29779));
    Odrv12 I__6314 (
            .O(N__29779),
            .I(\this_ppu.m18_i_o2_0 ));
    CascadeMux I__6313 (
            .O(N__29776),
            .I(N__29773));
    InMux I__6312 (
            .O(N__29773),
            .I(N__29770));
    LocalMux I__6311 (
            .O(N__29770),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_0 ));
    InMux I__6310 (
            .O(N__29767),
            .I(N__29761));
    CascadeMux I__6309 (
            .O(N__29766),
            .I(N__29757));
    InMux I__6308 (
            .O(N__29765),
            .I(N__29750));
    InMux I__6307 (
            .O(N__29764),
            .I(N__29747));
    LocalMux I__6306 (
            .O(N__29761),
            .I(N__29744));
    InMux I__6305 (
            .O(N__29760),
            .I(N__29737));
    InMux I__6304 (
            .O(N__29757),
            .I(N__29737));
    InMux I__6303 (
            .O(N__29756),
            .I(N__29737));
    InMux I__6302 (
            .O(N__29755),
            .I(N__29730));
    InMux I__6301 (
            .O(N__29754),
            .I(N__29730));
    InMux I__6300 (
            .O(N__29753),
            .I(N__29730));
    LocalMux I__6299 (
            .O(N__29750),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__6298 (
            .O(N__29747),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    Odrv4 I__6297 (
            .O(N__29744),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__6296 (
            .O(N__29737),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__6295 (
            .O(N__29730),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    InMux I__6294 (
            .O(N__29719),
            .I(N__29711));
    CascadeMux I__6293 (
            .O(N__29718),
            .I(N__29708));
    InMux I__6292 (
            .O(N__29717),
            .I(N__29698));
    InMux I__6291 (
            .O(N__29716),
            .I(N__29698));
    InMux I__6290 (
            .O(N__29715),
            .I(N__29693));
    InMux I__6289 (
            .O(N__29714),
            .I(N__29693));
    LocalMux I__6288 (
            .O(N__29711),
            .I(N__29690));
    InMux I__6287 (
            .O(N__29708),
            .I(N__29683));
    InMux I__6286 (
            .O(N__29707),
            .I(N__29683));
    InMux I__6285 (
            .O(N__29706),
            .I(N__29683));
    InMux I__6284 (
            .O(N__29705),
            .I(N__29676));
    InMux I__6283 (
            .O(N__29704),
            .I(N__29676));
    InMux I__6282 (
            .O(N__29703),
            .I(N__29676));
    LocalMux I__6281 (
            .O(N__29698),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__6280 (
            .O(N__29693),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    Odrv4 I__6279 (
            .O(N__29690),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__6278 (
            .O(N__29683),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__6277 (
            .O(N__29676),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    InMux I__6276 (
            .O(N__29665),
            .I(N__29662));
    LocalMux I__6275 (
            .O(N__29662),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_3_0_0 ));
    InMux I__6274 (
            .O(N__29659),
            .I(N__29655));
    InMux I__6273 (
            .O(N__29658),
            .I(N__29652));
    LocalMux I__6272 (
            .O(N__29655),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0 ));
    LocalMux I__6271 (
            .O(N__29652),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0 ));
    CascadeMux I__6270 (
            .O(N__29647),
            .I(N_814_0_cascade_));
    CascadeMux I__6269 (
            .O(N__29644),
            .I(N__29639));
    CascadeMux I__6268 (
            .O(N__29643),
            .I(N__29636));
    InMux I__6267 (
            .O(N__29642),
            .I(N__29632));
    InMux I__6266 (
            .O(N__29639),
            .I(N__29627));
    InMux I__6265 (
            .O(N__29636),
            .I(N__29627));
    InMux I__6264 (
            .O(N__29635),
            .I(N__29623));
    LocalMux I__6263 (
            .O(N__29632),
            .I(N__29613));
    LocalMux I__6262 (
            .O(N__29627),
            .I(N__29613));
    InMux I__6261 (
            .O(N__29626),
            .I(N__29610));
    LocalMux I__6260 (
            .O(N__29623),
            .I(N__29607));
    InMux I__6259 (
            .O(N__29622),
            .I(N__29602));
    InMux I__6258 (
            .O(N__29621),
            .I(N__29602));
    InMux I__6257 (
            .O(N__29620),
            .I(N__29599));
    InMux I__6256 (
            .O(N__29619),
            .I(N__29594));
    InMux I__6255 (
            .O(N__29618),
            .I(N__29594));
    Span4Mux_h I__6254 (
            .O(N__29613),
            .I(N__29591));
    LocalMux I__6253 (
            .O(N__29610),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    Odrv12 I__6252 (
            .O(N__29607),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__6251 (
            .O(N__29602),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__6250 (
            .O(N__29599),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__6249 (
            .O(N__29594),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    Odrv4 I__6248 (
            .O(N__29591),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    CascadeMux I__6247 (
            .O(N__29578),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_2_1_cascade_ ));
    CascadeMux I__6246 (
            .O(N__29575),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_2_2_cascade_ ));
    InMux I__6245 (
            .O(N__29572),
            .I(N__29566));
    InMux I__6244 (
            .O(N__29571),
            .I(N__29559));
    InMux I__6243 (
            .O(N__29570),
            .I(N__29559));
    InMux I__6242 (
            .O(N__29569),
            .I(N__29559));
    LocalMux I__6241 (
            .O(N__29566),
            .I(N__29554));
    LocalMux I__6240 (
            .O(N__29559),
            .I(N__29551));
    InMux I__6239 (
            .O(N__29558),
            .I(N__29546));
    InMux I__6238 (
            .O(N__29557),
            .I(N__29546));
    Span4Mux_v I__6237 (
            .O(N__29554),
            .I(N__29539));
    Span4Mux_v I__6236 (
            .O(N__29551),
            .I(N__29539));
    LocalMux I__6235 (
            .O(N__29546),
            .I(N__29539));
    Odrv4 I__6234 (
            .O(N__29539),
            .I(\this_vga_signals.mult1_un47_sum_c3_0 ));
    InMux I__6233 (
            .O(N__29536),
            .I(N__29533));
    LocalMux I__6232 (
            .O(N__29533),
            .I(N__29528));
    CascadeMux I__6231 (
            .O(N__29532),
            .I(N__29524));
    InMux I__6230 (
            .O(N__29531),
            .I(N__29519));
    Span4Mux_h I__6229 (
            .O(N__29528),
            .I(N__29516));
    InMux I__6228 (
            .O(N__29527),
            .I(N__29509));
    InMux I__6227 (
            .O(N__29524),
            .I(N__29509));
    InMux I__6226 (
            .O(N__29523),
            .I(N__29509));
    InMux I__6225 (
            .O(N__29522),
            .I(N__29506));
    LocalMux I__6224 (
            .O(N__29519),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_2_2 ));
    Odrv4 I__6223 (
            .O(N__29516),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_2_2 ));
    LocalMux I__6222 (
            .O(N__29509),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_2_2 ));
    LocalMux I__6221 (
            .O(N__29506),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_2_2 ));
    CascadeMux I__6220 (
            .O(N__29497),
            .I(N__29494));
    InMux I__6219 (
            .O(N__29494),
            .I(N__29491));
    LocalMux I__6218 (
            .O(N__29491),
            .I(N__29485));
    CascadeMux I__6217 (
            .O(N__29490),
            .I(N__29482));
    CascadeMux I__6216 (
            .O(N__29489),
            .I(N__29477));
    InMux I__6215 (
            .O(N__29488),
            .I(N__29473));
    Span4Mux_h I__6214 (
            .O(N__29485),
            .I(N__29470));
    InMux I__6213 (
            .O(N__29482),
            .I(N__29463));
    InMux I__6212 (
            .O(N__29481),
            .I(N__29463));
    InMux I__6211 (
            .O(N__29480),
            .I(N__29463));
    InMux I__6210 (
            .O(N__29477),
            .I(N__29458));
    InMux I__6209 (
            .O(N__29476),
            .I(N__29458));
    LocalMux I__6208 (
            .O(N__29473),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_2_0 ));
    Odrv4 I__6207 (
            .O(N__29470),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_2_0 ));
    LocalMux I__6206 (
            .O(N__29463),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_2_0 ));
    LocalMux I__6205 (
            .O(N__29458),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0_2_0 ));
    CascadeMux I__6204 (
            .O(N__29449),
            .I(N__29446));
    InMux I__6203 (
            .O(N__29446),
            .I(N__29442));
    CascadeMux I__6202 (
            .O(N__29445),
            .I(N__29439));
    LocalMux I__6201 (
            .O(N__29442),
            .I(N__29436));
    InMux I__6200 (
            .O(N__29439),
            .I(N__29433));
    Odrv4 I__6199 (
            .O(N__29436),
            .I(\this_ppu.N_1341 ));
    LocalMux I__6198 (
            .O(N__29433),
            .I(\this_ppu.N_1341 ));
    InMux I__6197 (
            .O(N__29428),
            .I(N__29424));
    InMux I__6196 (
            .O(N__29427),
            .I(N__29419));
    LocalMux I__6195 (
            .O(N__29424),
            .I(N__29415));
    InMux I__6194 (
            .O(N__29423),
            .I(N__29412));
    InMux I__6193 (
            .O(N__29422),
            .I(N__29408));
    LocalMux I__6192 (
            .O(N__29419),
            .I(N__29404));
    InMux I__6191 (
            .O(N__29418),
            .I(N__29401));
    Span4Mux_v I__6190 (
            .O(N__29415),
            .I(N__29396));
    LocalMux I__6189 (
            .O(N__29412),
            .I(N__29396));
    InMux I__6188 (
            .O(N__29411),
            .I(N__29393));
    LocalMux I__6187 (
            .O(N__29408),
            .I(N__29390));
    InMux I__6186 (
            .O(N__29407),
            .I(N__29387));
    Span4Mux_h I__6185 (
            .O(N__29404),
            .I(N__29384));
    LocalMux I__6184 (
            .O(N__29401),
            .I(N__29381));
    Span4Mux_v I__6183 (
            .O(N__29396),
            .I(N__29376));
    LocalMux I__6182 (
            .O(N__29393),
            .I(N__29376));
    Span12Mux_s4_v I__6181 (
            .O(N__29390),
            .I(N__29370));
    LocalMux I__6180 (
            .O(N__29387),
            .I(N__29370));
    Span4Mux_v I__6179 (
            .O(N__29384),
            .I(N__29365));
    Span4Mux_h I__6178 (
            .O(N__29381),
            .I(N__29365));
    Sp12to4 I__6177 (
            .O(N__29376),
            .I(N__29362));
    InMux I__6176 (
            .O(N__29375),
            .I(N__29359));
    Span12Mux_h I__6175 (
            .O(N__29370),
            .I(N__29356));
    Span4Mux_h I__6174 (
            .O(N__29365),
            .I(N__29353));
    Span12Mux_v I__6173 (
            .O(N__29362),
            .I(N__29348));
    LocalMux I__6172 (
            .O(N__29359),
            .I(N__29348));
    Odrv12 I__6171 (
            .O(N__29356),
            .I(M_this_spr_ram_write_data_2));
    Odrv4 I__6170 (
            .O(N__29353),
            .I(M_this_spr_ram_write_data_2));
    Odrv12 I__6169 (
            .O(N__29348),
            .I(M_this_spr_ram_write_data_2));
    InMux I__6168 (
            .O(N__29341),
            .I(N__29338));
    LocalMux I__6167 (
            .O(N__29338),
            .I(N__29335));
    Span4Mux_h I__6166 (
            .O(N__29335),
            .I(N__29332));
    Span4Mux_h I__6165 (
            .O(N__29332),
            .I(N__29329));
    Span4Mux_h I__6164 (
            .O(N__29329),
            .I(N__29326));
    Span4Mux_h I__6163 (
            .O(N__29326),
            .I(N__29323));
    Odrv4 I__6162 (
            .O(N__29323),
            .I(\this_ppu.oam_cache.mem_5 ));
    InMux I__6161 (
            .O(N__29320),
            .I(N__29317));
    LocalMux I__6160 (
            .O(N__29317),
            .I(N__29314));
    Span4Mux_h I__6159 (
            .O(N__29314),
            .I(N__29311));
    Odrv4 I__6158 (
            .O(N__29311),
            .I(\this_vga_signals.mult1_un54_sum_1_3 ));
    CascadeMux I__6157 (
            .O(N__29308),
            .I(\this_vga_signals.mult1_un47_sum_0_3_cascade_ ));
    InMux I__6156 (
            .O(N__29305),
            .I(N__29302));
    LocalMux I__6155 (
            .O(N__29302),
            .I(\this_vga_signals.N_7 ));
    CascadeMux I__6154 (
            .O(N__29299),
            .I(N__29296));
    InMux I__6153 (
            .O(N__29296),
            .I(N__29293));
    LocalMux I__6152 (
            .O(N__29293),
            .I(\this_vga_signals.mult1_un47_sum_2_3 ));
    InMux I__6151 (
            .O(N__29290),
            .I(N__29286));
    InMux I__6150 (
            .O(N__29289),
            .I(N__29282));
    LocalMux I__6149 (
            .O(N__29286),
            .I(N__29278));
    InMux I__6148 (
            .O(N__29285),
            .I(N__29275));
    LocalMux I__6147 (
            .O(N__29282),
            .I(N__29272));
    InMux I__6146 (
            .O(N__29281),
            .I(N__29268));
    Span12Mux_v I__6145 (
            .O(N__29278),
            .I(N__29263));
    LocalMux I__6144 (
            .O(N__29275),
            .I(N__29263));
    Span4Mux_v I__6143 (
            .O(N__29272),
            .I(N__29260));
    InMux I__6142 (
            .O(N__29271),
            .I(N__29257));
    LocalMux I__6141 (
            .O(N__29268),
            .I(M_this_state_qZ0Z_9));
    Odrv12 I__6140 (
            .O(N__29263),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__6139 (
            .O(N__29260),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__6138 (
            .O(N__29257),
            .I(M_this_state_qZ0Z_9));
    InMux I__6137 (
            .O(N__29248),
            .I(N__29245));
    LocalMux I__6136 (
            .O(N__29245),
            .I(N__29241));
    CascadeMux I__6135 (
            .O(N__29244),
            .I(N__29237));
    Span4Mux_v I__6134 (
            .O(N__29241),
            .I(N__29234));
    InMux I__6133 (
            .O(N__29240),
            .I(N__29231));
    InMux I__6132 (
            .O(N__29237),
            .I(N__29228));
    Span4Mux_h I__6131 (
            .O(N__29234),
            .I(N__29223));
    LocalMux I__6130 (
            .O(N__29231),
            .I(N__29223));
    LocalMux I__6129 (
            .O(N__29228),
            .I(N__29216));
    Span4Mux_h I__6128 (
            .O(N__29223),
            .I(N__29216));
    InMux I__6127 (
            .O(N__29222),
            .I(N__29211));
    InMux I__6126 (
            .O(N__29221),
            .I(N__29211));
    Odrv4 I__6125 (
            .O(N__29216),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__6124 (
            .O(N__29211),
            .I(M_this_state_qZ0Z_11));
    CascadeMux I__6123 (
            .O(N__29206),
            .I(N__29202));
    InMux I__6122 (
            .O(N__29205),
            .I(N__29198));
    InMux I__6121 (
            .O(N__29202),
            .I(N__29195));
    InMux I__6120 (
            .O(N__29201),
            .I(N__29191));
    LocalMux I__6119 (
            .O(N__29198),
            .I(N__29185));
    LocalMux I__6118 (
            .O(N__29195),
            .I(N__29185));
    InMux I__6117 (
            .O(N__29194),
            .I(N__29182));
    LocalMux I__6116 (
            .O(N__29191),
            .I(N__29179));
    InMux I__6115 (
            .O(N__29190),
            .I(N__29176));
    Span4Mux_v I__6114 (
            .O(N__29185),
            .I(N__29171));
    LocalMux I__6113 (
            .O(N__29182),
            .I(N__29171));
    Span4Mux_h I__6112 (
            .O(N__29179),
            .I(N__29168));
    LocalMux I__6111 (
            .O(N__29176),
            .I(\this_ppu.N_1301 ));
    Odrv4 I__6110 (
            .O(N__29171),
            .I(\this_ppu.N_1301 ));
    Odrv4 I__6109 (
            .O(N__29168),
            .I(\this_ppu.N_1301 ));
    InMux I__6108 (
            .O(N__29161),
            .I(N__29158));
    LocalMux I__6107 (
            .O(N__29158),
            .I(\this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_15 ));
    CascadeMux I__6106 (
            .O(N__29155),
            .I(N__29152));
    InMux I__6105 (
            .O(N__29152),
            .I(N__29148));
    CascadeMux I__6104 (
            .O(N__29151),
            .I(N__29145));
    LocalMux I__6103 (
            .O(N__29148),
            .I(N__29139));
    InMux I__6102 (
            .O(N__29145),
            .I(N__29136));
    InMux I__6101 (
            .O(N__29144),
            .I(N__29133));
    InMux I__6100 (
            .O(N__29143),
            .I(N__29128));
    InMux I__6099 (
            .O(N__29142),
            .I(N__29128));
    Span4Mux_v I__6098 (
            .O(N__29139),
            .I(N__29121));
    LocalMux I__6097 (
            .O(N__29136),
            .I(N__29121));
    LocalMux I__6096 (
            .O(N__29133),
            .I(N__29121));
    LocalMux I__6095 (
            .O(N__29128),
            .I(M_this_state_qZ0Z_15));
    Odrv4 I__6094 (
            .O(N__29121),
            .I(M_this_state_qZ0Z_15));
    CascadeMux I__6093 (
            .O(N__29116),
            .I(N__29113));
    InMux I__6092 (
            .O(N__29113),
            .I(N__29110));
    LocalMux I__6091 (
            .O(N__29110),
            .I(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_7 ));
    InMux I__6090 (
            .O(N__29107),
            .I(N__29104));
    LocalMux I__6089 (
            .O(N__29104),
            .I(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_11 ));
    CascadeMux I__6088 (
            .O(N__29101),
            .I(N__29098));
    InMux I__6087 (
            .O(N__29098),
            .I(N__29095));
    LocalMux I__6086 (
            .O(N__29095),
            .I(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_8 ));
    CascadeMux I__6085 (
            .O(N__29092),
            .I(\this_ppu.N_807_0_cascade_ ));
    InMux I__6084 (
            .O(N__29089),
            .I(N__29086));
    LocalMux I__6083 (
            .O(N__29086),
            .I(N__29083));
    Span4Mux_v I__6082 (
            .O(N__29083),
            .I(N__29077));
    InMux I__6081 (
            .O(N__29082),
            .I(N__29074));
    InMux I__6080 (
            .O(N__29081),
            .I(N__29069));
    InMux I__6079 (
            .O(N__29080),
            .I(N__29069));
    Odrv4 I__6078 (
            .O(N__29077),
            .I(\this_ppu.N_1002_0 ));
    LocalMux I__6077 (
            .O(N__29074),
            .I(\this_ppu.N_1002_0 ));
    LocalMux I__6076 (
            .O(N__29069),
            .I(\this_ppu.N_1002_0 ));
    InMux I__6075 (
            .O(N__29062),
            .I(N__29059));
    LocalMux I__6074 (
            .O(N__29059),
            .I(\this_ppu.N_235_2_0 ));
    CascadeMux I__6073 (
            .O(N__29056),
            .I(\this_ppu.N_235_2_0_cascade_ ));
    InMux I__6072 (
            .O(N__29053),
            .I(N__29047));
    InMux I__6071 (
            .O(N__29052),
            .I(N__29047));
    LocalMux I__6070 (
            .O(N__29047),
            .I(N__29043));
    InMux I__6069 (
            .O(N__29046),
            .I(N__29038));
    Span4Mux_h I__6068 (
            .O(N__29043),
            .I(N__29035));
    InMux I__6067 (
            .O(N__29042),
            .I(N__29032));
    InMux I__6066 (
            .O(N__29041),
            .I(N__29029));
    LocalMux I__6065 (
            .O(N__29038),
            .I(M_this_state_qZ0Z_7));
    Odrv4 I__6064 (
            .O(N__29035),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__6063 (
            .O(N__29032),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__6062 (
            .O(N__29029),
            .I(M_this_state_qZ0Z_7));
    InMux I__6061 (
            .O(N__29020),
            .I(N__29017));
    LocalMux I__6060 (
            .O(N__29017),
            .I(\this_ppu.N_1162 ));
    InMux I__6059 (
            .O(N__29014),
            .I(N__29011));
    LocalMux I__6058 (
            .O(N__29011),
            .I(\this_vga_signals.g0_5 ));
    CascadeMux I__6057 (
            .O(N__29008),
            .I(N__29004));
    InMux I__6056 (
            .O(N__29007),
            .I(N__28999));
    InMux I__6055 (
            .O(N__29004),
            .I(N__28992));
    InMux I__6054 (
            .O(N__29003),
            .I(N__28992));
    InMux I__6053 (
            .O(N__29002),
            .I(N__28992));
    LocalMux I__6052 (
            .O(N__28999),
            .I(\this_vga_signals.mult1_un61_sum_axb1_0 ));
    LocalMux I__6051 (
            .O(N__28992),
            .I(\this_vga_signals.mult1_un61_sum_axb1_0 ));
    CascadeMux I__6050 (
            .O(N__28987),
            .I(N__28983));
    CascadeMux I__6049 (
            .O(N__28986),
            .I(N__28978));
    InMux I__6048 (
            .O(N__28983),
            .I(N__28972));
    InMux I__6047 (
            .O(N__28982),
            .I(N__28972));
    InMux I__6046 (
            .O(N__28981),
            .I(N__28969));
    InMux I__6045 (
            .O(N__28978),
            .I(N__28964));
    InMux I__6044 (
            .O(N__28977),
            .I(N__28964));
    LocalMux I__6043 (
            .O(N__28972),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__6042 (
            .O(N__28969),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__6041 (
            .O(N__28964),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    InMux I__6040 (
            .O(N__28957),
            .I(N__28954));
    LocalMux I__6039 (
            .O(N__28954),
            .I(N__28951));
    Odrv4 I__6038 (
            .O(N__28951),
            .I(\this_vga_signals.g0_1_0 ));
    InMux I__6037 (
            .O(N__28948),
            .I(N__28944));
    CascadeMux I__6036 (
            .O(N__28947),
            .I(N__28941));
    LocalMux I__6035 (
            .O(N__28944),
            .I(N__28938));
    InMux I__6034 (
            .O(N__28941),
            .I(N__28932));
    Span4Mux_h I__6033 (
            .O(N__28938),
            .I(N__28925));
    InMux I__6032 (
            .O(N__28937),
            .I(N__28918));
    InMux I__6031 (
            .O(N__28936),
            .I(N__28918));
    InMux I__6030 (
            .O(N__28935),
            .I(N__28918));
    LocalMux I__6029 (
            .O(N__28932),
            .I(N__28915));
    InMux I__6028 (
            .O(N__28931),
            .I(N__28910));
    InMux I__6027 (
            .O(N__28930),
            .I(N__28910));
    CascadeMux I__6026 (
            .O(N__28929),
            .I(N__28906));
    InMux I__6025 (
            .O(N__28928),
            .I(N__28900));
    Span4Mux_h I__6024 (
            .O(N__28925),
            .I(N__28897));
    LocalMux I__6023 (
            .O(N__28918),
            .I(N__28894));
    Span4Mux_v I__6022 (
            .O(N__28915),
            .I(N__28891));
    LocalMux I__6021 (
            .O(N__28910),
            .I(N__28888));
    InMux I__6020 (
            .O(N__28909),
            .I(N__28885));
    InMux I__6019 (
            .O(N__28906),
            .I(N__28880));
    InMux I__6018 (
            .O(N__28905),
            .I(N__28880));
    InMux I__6017 (
            .O(N__28904),
            .I(N__28875));
    InMux I__6016 (
            .O(N__28903),
            .I(N__28875));
    LocalMux I__6015 (
            .O(N__28900),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__6014 (
            .O(N__28897),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__6013 (
            .O(N__28894),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__6012 (
            .O(N__28891),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__6011 (
            .O(N__28888),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__6010 (
            .O(N__28885),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__6009 (
            .O(N__28880),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__6008 (
            .O(N__28875),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    InMux I__6007 (
            .O(N__28858),
            .I(N__28852));
    InMux I__6006 (
            .O(N__28857),
            .I(N__28849));
    InMux I__6005 (
            .O(N__28856),
            .I(N__28844));
    InMux I__6004 (
            .O(N__28855),
            .I(N__28844));
    LocalMux I__6003 (
            .O(N__28852),
            .I(\this_vga_signals.mult1_un61_sum_c3_0 ));
    LocalMux I__6002 (
            .O(N__28849),
            .I(\this_vga_signals.mult1_un61_sum_c3_0 ));
    LocalMux I__6001 (
            .O(N__28844),
            .I(\this_vga_signals.mult1_un61_sum_c3_0 ));
    CascadeMux I__6000 (
            .O(N__28837),
            .I(\this_vga_signals.mult1_un68_sum_c2_0_cascade_ ));
    InMux I__5999 (
            .O(N__28834),
            .I(N__28831));
    LocalMux I__5998 (
            .O(N__28831),
            .I(\this_vga_signals.g0_0_3_1 ));
    InMux I__5997 (
            .O(N__28828),
            .I(N__28825));
    LocalMux I__5996 (
            .O(N__28825),
            .I(\this_vga_signals.g0_0_3 ));
    InMux I__5995 (
            .O(N__28822),
            .I(N__28819));
    LocalMux I__5994 (
            .O(N__28819),
            .I(N__28816));
    Odrv4 I__5993 (
            .O(N__28816),
            .I(\this_vga_signals.g1_1 ));
    CascadeMux I__5992 (
            .O(N__28813),
            .I(N__28810));
    InMux I__5991 (
            .O(N__28810),
            .I(N__28807));
    LocalMux I__5990 (
            .O(N__28807),
            .I(N__28804));
    Span4Mux_v I__5989 (
            .O(N__28804),
            .I(N__28801));
    Odrv4 I__5988 (
            .O(N__28801),
            .I(\this_vga_signals.mult1_un54_sum_0_1 ));
    InMux I__5987 (
            .O(N__28798),
            .I(N__28795));
    LocalMux I__5986 (
            .O(N__28795),
            .I(\this_vga_signals.g0_2_0 ));
    InMux I__5985 (
            .O(N__28792),
            .I(N__28789));
    LocalMux I__5984 (
            .O(N__28789),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_0 ));
    InMux I__5983 (
            .O(N__28786),
            .I(N__28781));
    InMux I__5982 (
            .O(N__28785),
            .I(N__28776));
    InMux I__5981 (
            .O(N__28784),
            .I(N__28776));
    LocalMux I__5980 (
            .O(N__28781),
            .I(\this_vga_signals.vaddress_9 ));
    LocalMux I__5979 (
            .O(N__28776),
            .I(\this_vga_signals.vaddress_9 ));
    InMux I__5978 (
            .O(N__28771),
            .I(N__28761));
    InMux I__5977 (
            .O(N__28770),
            .I(N__28761));
    InMux I__5976 (
            .O(N__28769),
            .I(N__28758));
    InMux I__5975 (
            .O(N__28768),
            .I(N__28755));
    InMux I__5974 (
            .O(N__28767),
            .I(N__28750));
    InMux I__5973 (
            .O(N__28766),
            .I(N__28750));
    LocalMux I__5972 (
            .O(N__28761),
            .I(N__28745));
    LocalMux I__5971 (
            .O(N__28758),
            .I(N__28742));
    LocalMux I__5970 (
            .O(N__28755),
            .I(N__28737));
    LocalMux I__5969 (
            .O(N__28750),
            .I(N__28737));
    InMux I__5968 (
            .O(N__28749),
            .I(N__28732));
    InMux I__5967 (
            .O(N__28748),
            .I(N__28732));
    Span4Mux_v I__5966 (
            .O(N__28745),
            .I(N__28729));
    Span4Mux_h I__5965 (
            .O(N__28742),
            .I(N__28726));
    Odrv12 I__5964 (
            .O(N__28737),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_1 ));
    LocalMux I__5963 (
            .O(N__28732),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_1 ));
    Odrv4 I__5962 (
            .O(N__28729),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_1 ));
    Odrv4 I__5961 (
            .O(N__28726),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_1 ));
    CascadeMux I__5960 (
            .O(N__28717),
            .I(N__28714));
    InMux I__5959 (
            .O(N__28714),
            .I(N__28706));
    InMux I__5958 (
            .O(N__28713),
            .I(N__28706));
    InMux I__5957 (
            .O(N__28712),
            .I(N__28697));
    InMux I__5956 (
            .O(N__28711),
            .I(N__28697));
    LocalMux I__5955 (
            .O(N__28706),
            .I(N__28694));
    InMux I__5954 (
            .O(N__28705),
            .I(N__28690));
    InMux I__5953 (
            .O(N__28704),
            .I(N__28683));
    InMux I__5952 (
            .O(N__28703),
            .I(N__28683));
    InMux I__5951 (
            .O(N__28702),
            .I(N__28683));
    LocalMux I__5950 (
            .O(N__28697),
            .I(N__28678));
    Span4Mux_h I__5949 (
            .O(N__28694),
            .I(N__28678));
    InMux I__5948 (
            .O(N__28693),
            .I(N__28675));
    LocalMux I__5947 (
            .O(N__28690),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__5946 (
            .O(N__28683),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    Odrv4 I__5945 (
            .O(N__28678),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    LocalMux I__5944 (
            .O(N__28675),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ));
    InMux I__5943 (
            .O(N__28666),
            .I(N__28661));
    InMux I__5942 (
            .O(N__28665),
            .I(N__28658));
    InMux I__5941 (
            .O(N__28664),
            .I(N__28655));
    LocalMux I__5940 (
            .O(N__28661),
            .I(N__28652));
    LocalMux I__5939 (
            .O(N__28658),
            .I(N__28645));
    LocalMux I__5938 (
            .O(N__28655),
            .I(N__28642));
    Span4Mux_h I__5937 (
            .O(N__28652),
            .I(N__28639));
    InMux I__5936 (
            .O(N__28651),
            .I(N__28634));
    InMux I__5935 (
            .O(N__28650),
            .I(N__28634));
    InMux I__5934 (
            .O(N__28649),
            .I(N__28629));
    InMux I__5933 (
            .O(N__28648),
            .I(N__28629));
    Odrv4 I__5932 (
            .O(N__28645),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    Odrv12 I__5931 (
            .O(N__28642),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    Odrv4 I__5930 (
            .O(N__28639),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    LocalMux I__5929 (
            .O(N__28634),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    LocalMux I__5928 (
            .O(N__28629),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    CascadeMux I__5927 (
            .O(N__28618),
            .I(N__28615));
    InMux I__5926 (
            .O(N__28615),
            .I(N__28612));
    LocalMux I__5925 (
            .O(N__28612),
            .I(N__28609));
    Span4Mux_h I__5924 (
            .O(N__28609),
            .I(N__28606));
    Odrv4 I__5923 (
            .O(N__28606),
            .I(\this_vga_signals.g0_0_x2 ));
    InMux I__5922 (
            .O(N__28603),
            .I(N__28600));
    LocalMux I__5921 (
            .O(N__28600),
            .I(\this_vga_signals.if_m5_i_0_0_0 ));
    InMux I__5920 (
            .O(N__28597),
            .I(N__28594));
    LocalMux I__5919 (
            .O(N__28594),
            .I(\this_vga_signals.mult1_un54_sum_c3_x0 ));
    CascadeMux I__5918 (
            .O(N__28591),
            .I(\this_vga_signals.if_N_7_0_cascade_ ));
    InMux I__5917 (
            .O(N__28588),
            .I(N__28585));
    LocalMux I__5916 (
            .O(N__28585),
            .I(N__28581));
    InMux I__5915 (
            .O(N__28584),
            .I(N__28578));
    Span4Mux_v I__5914 (
            .O(N__28581),
            .I(N__28575));
    LocalMux I__5913 (
            .O(N__28578),
            .I(N__28572));
    Span4Mux_v I__5912 (
            .O(N__28575),
            .I(N__28569));
    Odrv12 I__5911 (
            .O(N__28572),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    Odrv4 I__5910 (
            .O(N__28569),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    CascadeMux I__5909 (
            .O(N__28564),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d_cascade_ ));
    CascadeMux I__5908 (
            .O(N__28561),
            .I(N__28558));
    InMux I__5907 (
            .O(N__28558),
            .I(N__28555));
    LocalMux I__5906 (
            .O(N__28555),
            .I(N__28552));
    Odrv4 I__5905 (
            .O(N__28552),
            .I(\this_vga_signals.mult1_un47_sum_1_3 ));
    InMux I__5904 (
            .O(N__28549),
            .I(N__28546));
    LocalMux I__5903 (
            .O(N__28546),
            .I(N__28543));
    Odrv4 I__5902 (
            .O(N__28543),
            .I(\this_vga_signals.mult1_un54_sum_1_1 ));
    InMux I__5901 (
            .O(N__28540),
            .I(N__28536));
    InMux I__5900 (
            .O(N__28539),
            .I(N__28533));
    LocalMux I__5899 (
            .O(N__28536),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c ));
    LocalMux I__5898 (
            .O(N__28533),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c ));
    CascadeMux I__5897 (
            .O(N__28528),
            .I(\this_vga_signals.mult1_un54_sum_0_3_cascade_ ));
    InMux I__5896 (
            .O(N__28525),
            .I(N__28521));
    InMux I__5895 (
            .O(N__28524),
            .I(N__28518));
    LocalMux I__5894 (
            .O(N__28521),
            .I(N__28513));
    LocalMux I__5893 (
            .O(N__28518),
            .I(N__28510));
    InMux I__5892 (
            .O(N__28517),
            .I(N__28507));
    InMux I__5891 (
            .O(N__28516),
            .I(N__28504));
    Span4Mux_h I__5890 (
            .O(N__28513),
            .I(N__28501));
    Odrv4 I__5889 (
            .O(N__28510),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d ));
    LocalMux I__5888 (
            .O(N__28507),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d ));
    LocalMux I__5887 (
            .O(N__28504),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d ));
    Odrv4 I__5886 (
            .O(N__28501),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d ));
    CascadeMux I__5885 (
            .O(N__28492),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_1_cascade_ ));
    InMux I__5884 (
            .O(N__28489),
            .I(N__28486));
    LocalMux I__5883 (
            .O(N__28486),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0 ));
    InMux I__5882 (
            .O(N__28483),
            .I(N__28480));
    LocalMux I__5881 (
            .O(N__28480),
            .I(N__28477));
    Odrv12 I__5880 (
            .O(N__28477),
            .I(\this_vga_signals.N_3_1_0_1 ));
    CascadeMux I__5879 (
            .O(N__28474),
            .I(N__28471));
    InMux I__5878 (
            .O(N__28471),
            .I(N__28468));
    LocalMux I__5877 (
            .O(N__28468),
            .I(N__28465));
    Span4Mux_h I__5876 (
            .O(N__28465),
            .I(N__28462));
    Odrv4 I__5875 (
            .O(N__28462),
            .I(\this_vga_signals.g0_2_1 ));
    CascadeMux I__5874 (
            .O(N__28459),
            .I(\this_vga_signals.mult1_un54_sum_c2_0_cascade_ ));
    InMux I__5873 (
            .O(N__28456),
            .I(N__28453));
    LocalMux I__5872 (
            .O(N__28453),
            .I(N__28450));
    Odrv4 I__5871 (
            .O(N__28450),
            .I(\this_vga_signals.g0_4 ));
    CascadeMux I__5870 (
            .O(N__28447),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ));
    InMux I__5869 (
            .O(N__28444),
            .I(N__28441));
    LocalMux I__5868 (
            .O(N__28441),
            .I(\this_vga_signals.mult1_un47_sum_4_3 ));
    CascadeMux I__5867 (
            .O(N__28438),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1_cascade_ ));
    CascadeMux I__5866 (
            .O(N__28435),
            .I(N__28432));
    InMux I__5865 (
            .O(N__28432),
            .I(N__28429));
    LocalMux I__5864 (
            .O(N__28429),
            .I(\this_vga_signals.mult1_un54_sum_c3_x1 ));
    InMux I__5863 (
            .O(N__28426),
            .I(N__28420));
    InMux I__5862 (
            .O(N__28425),
            .I(N__28417));
    InMux I__5861 (
            .O(N__28424),
            .I(N__28414));
    InMux I__5860 (
            .O(N__28423),
            .I(N__28411));
    LocalMux I__5859 (
            .O(N__28420),
            .I(N__28408));
    LocalMux I__5858 (
            .O(N__28417),
            .I(N__28403));
    LocalMux I__5857 (
            .O(N__28414),
            .I(N__28403));
    LocalMux I__5856 (
            .O(N__28411),
            .I(N__28400));
    Span4Mux_h I__5855 (
            .O(N__28408),
            .I(N__28397));
    Span4Mux_v I__5854 (
            .O(N__28403),
            .I(N__28392));
    Span4Mux_h I__5853 (
            .O(N__28400),
            .I(N__28392));
    Odrv4 I__5852 (
            .O(N__28397),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_3 ));
    Odrv4 I__5851 (
            .O(N__28392),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_3 ));
    InMux I__5850 (
            .O(N__28387),
            .I(N__28384));
    LocalMux I__5849 (
            .O(N__28384),
            .I(N__28380));
    InMux I__5848 (
            .O(N__28383),
            .I(N__28377));
    Span4Mux_h I__5847 (
            .O(N__28380),
            .I(N__28374));
    LocalMux I__5846 (
            .O(N__28377),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1 ));
    Odrv4 I__5845 (
            .O(N__28374),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1 ));
    InMux I__5844 (
            .O(N__28369),
            .I(N__28366));
    LocalMux I__5843 (
            .O(N__28366),
            .I(\this_vga_signals.N_27_0 ));
    InMux I__5842 (
            .O(N__28363),
            .I(N__28360));
    LocalMux I__5841 (
            .O(N__28360),
            .I(N__28356));
    InMux I__5840 (
            .O(N__28359),
            .I(N__28353));
    Span4Mux_v I__5839 (
            .O(N__28356),
            .I(N__28350));
    LocalMux I__5838 (
            .O(N__28353),
            .I(N__28347));
    Span4Mux_h I__5837 (
            .O(N__28350),
            .I(N__28344));
    Span4Mux_v I__5836 (
            .O(N__28347),
            .I(N__28341));
    Odrv4 I__5835 (
            .O(N__28344),
            .I(\this_vga_signals.N_1247 ));
    Odrv4 I__5834 (
            .O(N__28341),
            .I(\this_vga_signals.N_1247 ));
    CascadeMux I__5833 (
            .O(N__28336),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0_cascade_ ));
    InMux I__5832 (
            .O(N__28333),
            .I(N__28329));
    InMux I__5831 (
            .O(N__28332),
            .I(N__28326));
    LocalMux I__5830 (
            .O(N__28329),
            .I(N__28322));
    LocalMux I__5829 (
            .O(N__28326),
            .I(N__28319));
    InMux I__5828 (
            .O(N__28325),
            .I(N__28316));
    Span12Mux_v I__5827 (
            .O(N__28322),
            .I(N__28313));
    Span4Mux_v I__5826 (
            .O(N__28319),
            .I(N__28310));
    LocalMux I__5825 (
            .O(N__28316),
            .I(N__28307));
    Odrv12 I__5824 (
            .O(N__28313),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    Odrv4 I__5823 (
            .O(N__28310),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    Odrv12 I__5822 (
            .O(N__28307),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    InMux I__5821 (
            .O(N__28300),
            .I(N__28297));
    LocalMux I__5820 (
            .O(N__28297),
            .I(N__28294));
    Span4Mux_v I__5819 (
            .O(N__28294),
            .I(N__28289));
    InMux I__5818 (
            .O(N__28293),
            .I(N__28286));
    InMux I__5817 (
            .O(N__28292),
            .I(N__28283));
    Span4Mux_v I__5816 (
            .O(N__28289),
            .I(N__28280));
    LocalMux I__5815 (
            .O(N__28286),
            .I(N__28275));
    LocalMux I__5814 (
            .O(N__28283),
            .I(N__28275));
    Odrv4 I__5813 (
            .O(N__28280),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    Odrv12 I__5812 (
            .O(N__28275),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    InMux I__5811 (
            .O(N__28270),
            .I(N__28264));
    InMux I__5810 (
            .O(N__28269),
            .I(N__28264));
    LocalMux I__5809 (
            .O(N__28264),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    InMux I__5808 (
            .O(N__28261),
            .I(N__28257));
    CascadeMux I__5807 (
            .O(N__28260),
            .I(N__28254));
    LocalMux I__5806 (
            .O(N__28257),
            .I(N__28250));
    InMux I__5805 (
            .O(N__28254),
            .I(N__28247));
    InMux I__5804 (
            .O(N__28253),
            .I(N__28244));
    Odrv4 I__5803 (
            .O(N__28250),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__5802 (
            .O(N__28247),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__5801 (
            .O(N__28244),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    InMux I__5800 (
            .O(N__28237),
            .I(N__28234));
    LocalMux I__5799 (
            .O(N__28234),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_1_1_1 ));
    InMux I__5798 (
            .O(N__28231),
            .I(N__28224));
    InMux I__5797 (
            .O(N__28230),
            .I(N__28224));
    InMux I__5796 (
            .O(N__28229),
            .I(N__28221));
    LocalMux I__5795 (
            .O(N__28224),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    LocalMux I__5794 (
            .O(N__28221),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    CascadeMux I__5793 (
            .O(N__28216),
            .I(N__28212));
    InMux I__5792 (
            .O(N__28215),
            .I(N__28209));
    InMux I__5791 (
            .O(N__28212),
            .I(N__28206));
    LocalMux I__5790 (
            .O(N__28209),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    LocalMux I__5789 (
            .O(N__28206),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    InMux I__5788 (
            .O(N__28201),
            .I(N__28197));
    InMux I__5787 (
            .O(N__28200),
            .I(N__28191));
    LocalMux I__5786 (
            .O(N__28197),
            .I(N__28188));
    InMux I__5785 (
            .O(N__28196),
            .I(N__28185));
    InMux I__5784 (
            .O(N__28195),
            .I(N__28180));
    InMux I__5783 (
            .O(N__28194),
            .I(N__28180));
    LocalMux I__5782 (
            .O(N__28191),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__5781 (
            .O(N__28188),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__5780 (
            .O(N__28185),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__5779 (
            .O(N__28180),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    CascadeMux I__5778 (
            .O(N__28171),
            .I(\this_vga_signals.mult1_un54_sum_axb1_cascade_ ));
    InMux I__5777 (
            .O(N__28168),
            .I(N__28157));
    InMux I__5776 (
            .O(N__28167),
            .I(N__28157));
    InMux I__5775 (
            .O(N__28166),
            .I(N__28150));
    InMux I__5774 (
            .O(N__28165),
            .I(N__28150));
    InMux I__5773 (
            .O(N__28164),
            .I(N__28150));
    InMux I__5772 (
            .O(N__28163),
            .I(N__28145));
    InMux I__5771 (
            .O(N__28162),
            .I(N__28145));
    LocalMux I__5770 (
            .O(N__28157),
            .I(M_this_state_qZ0Z_18));
    LocalMux I__5769 (
            .O(N__28150),
            .I(M_this_state_qZ0Z_18));
    LocalMux I__5768 (
            .O(N__28145),
            .I(M_this_state_qZ0Z_18));
    InMux I__5767 (
            .O(N__28138),
            .I(N__28135));
    LocalMux I__5766 (
            .O(N__28135),
            .I(N__28132));
    Odrv12 I__5765 (
            .O(N__28132),
            .I(this_ppu_M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0));
    CascadeMux I__5764 (
            .O(N__28129),
            .I(\this_ppu.N_1322_cascade_ ));
    InMux I__5763 (
            .O(N__28126),
            .I(N__28123));
    LocalMux I__5762 (
            .O(N__28123),
            .I(N__28119));
    InMux I__5761 (
            .O(N__28122),
            .I(N__28116));
    Span4Mux_v I__5760 (
            .O(N__28119),
            .I(N__28109));
    LocalMux I__5759 (
            .O(N__28116),
            .I(N__28109));
    InMux I__5758 (
            .O(N__28115),
            .I(N__28106));
    InMux I__5757 (
            .O(N__28114),
            .I(N__28102));
    Span4Mux_v I__5756 (
            .O(N__28109),
            .I(N__28097));
    LocalMux I__5755 (
            .O(N__28106),
            .I(N__28097));
    InMux I__5754 (
            .O(N__28105),
            .I(N__28094));
    LocalMux I__5753 (
            .O(N__28102),
            .I(N__28090));
    Span4Mux_v I__5752 (
            .O(N__28097),
            .I(N__28085));
    LocalMux I__5751 (
            .O(N__28094),
            .I(N__28085));
    InMux I__5750 (
            .O(N__28093),
            .I(N__28082));
    Span4Mux_h I__5749 (
            .O(N__28090),
            .I(N__28077));
    Span4Mux_v I__5748 (
            .O(N__28085),
            .I(N__28072));
    LocalMux I__5747 (
            .O(N__28082),
            .I(N__28072));
    InMux I__5746 (
            .O(N__28081),
            .I(N__28069));
    InMux I__5745 (
            .O(N__28080),
            .I(N__28066));
    Span4Mux_h I__5744 (
            .O(N__28077),
            .I(N__28063));
    Span4Mux_v I__5743 (
            .O(N__28072),
            .I(N__28058));
    LocalMux I__5742 (
            .O(N__28069),
            .I(N__28058));
    LocalMux I__5741 (
            .O(N__28066),
            .I(N__28055));
    Span4Mux_h I__5740 (
            .O(N__28063),
            .I(N__28052));
    Span4Mux_v I__5739 (
            .O(N__28058),
            .I(N__28047));
    Span4Mux_v I__5738 (
            .O(N__28055),
            .I(N__28047));
    Span4Mux_v I__5737 (
            .O(N__28052),
            .I(N__28042));
    Span4Mux_h I__5736 (
            .O(N__28047),
            .I(N__28042));
    Odrv4 I__5735 (
            .O(N__28042),
            .I(M_this_spr_ram_write_data_0));
    InMux I__5734 (
            .O(N__28039),
            .I(N__28035));
    InMux I__5733 (
            .O(N__28038),
            .I(N__28032));
    LocalMux I__5732 (
            .O(N__28035),
            .I(N__28026));
    LocalMux I__5731 (
            .O(N__28032),
            .I(N__28023));
    CascadeMux I__5730 (
            .O(N__28031),
            .I(N__28020));
    InMux I__5729 (
            .O(N__28030),
            .I(N__28015));
    InMux I__5728 (
            .O(N__28029),
            .I(N__28015));
    Span4Mux_h I__5727 (
            .O(N__28026),
            .I(N__28012));
    Span4Mux_h I__5726 (
            .O(N__28023),
            .I(N__28009));
    InMux I__5725 (
            .O(N__28020),
            .I(N__28006));
    LocalMux I__5724 (
            .O(N__28015),
            .I(N__28003));
    Odrv4 I__5723 (
            .O(N__28012),
            .I(this_vga_signals_CO0_0_i_i));
    Odrv4 I__5722 (
            .O(N__28009),
            .I(this_vga_signals_CO0_0_i_i));
    LocalMux I__5721 (
            .O(N__28006),
            .I(this_vga_signals_CO0_0_i_i));
    Odrv4 I__5720 (
            .O(N__28003),
            .I(this_vga_signals_CO0_0_i_i));
    CascadeMux I__5719 (
            .O(N__27994),
            .I(this_vga_signals_CO0_0_i_i_cascade_));
    InMux I__5718 (
            .O(N__27991),
            .I(N__27986));
    CascadeMux I__5717 (
            .O(N__27990),
            .I(N__27983));
    InMux I__5716 (
            .O(N__27989),
            .I(N__27979));
    LocalMux I__5715 (
            .O(N__27986),
            .I(N__27976));
    InMux I__5714 (
            .O(N__27983),
            .I(N__27971));
    InMux I__5713 (
            .O(N__27982),
            .I(N__27971));
    LocalMux I__5712 (
            .O(N__27979),
            .I(\this_vga_signals.vaddress_8 ));
    Odrv4 I__5711 (
            .O(N__27976),
            .I(\this_vga_signals.vaddress_8 ));
    LocalMux I__5710 (
            .O(N__27971),
            .I(\this_vga_signals.vaddress_8 ));
    InMux I__5709 (
            .O(N__27964),
            .I(N__27961));
    LocalMux I__5708 (
            .O(N__27961),
            .I(\this_vga_signals.g1 ));
    InMux I__5707 (
            .O(N__27958),
            .I(N__27953));
    InMux I__5706 (
            .O(N__27957),
            .I(N__27950));
    InMux I__5705 (
            .O(N__27956),
            .I(N__27946));
    LocalMux I__5704 (
            .O(N__27953),
            .I(N__27940));
    LocalMux I__5703 (
            .O(N__27950),
            .I(N__27940));
    InMux I__5702 (
            .O(N__27949),
            .I(N__27937));
    LocalMux I__5701 (
            .O(N__27946),
            .I(N__27934));
    InMux I__5700 (
            .O(N__27945),
            .I(N__27931));
    Span4Mux_v I__5699 (
            .O(N__27940),
            .I(N__27922));
    LocalMux I__5698 (
            .O(N__27937),
            .I(N__27922));
    Span4Mux_h I__5697 (
            .O(N__27934),
            .I(N__27922));
    LocalMux I__5696 (
            .O(N__27931),
            .I(N__27922));
    Odrv4 I__5695 (
            .O(N__27922),
            .I(\this_vga_signals.N_39_0 ));
    CascadeMux I__5694 (
            .O(N__27919),
            .I(N__27916));
    InMux I__5693 (
            .O(N__27916),
            .I(N__27911));
    InMux I__5692 (
            .O(N__27915),
            .I(N__27906));
    InMux I__5691 (
            .O(N__27914),
            .I(N__27903));
    LocalMux I__5690 (
            .O(N__27911),
            .I(N__27900));
    InMux I__5689 (
            .O(N__27910),
            .I(N__27897));
    InMux I__5688 (
            .O(N__27909),
            .I(N__27894));
    LocalMux I__5687 (
            .O(N__27906),
            .I(\this_vga_signals.vaddress_7 ));
    LocalMux I__5686 (
            .O(N__27903),
            .I(\this_vga_signals.vaddress_7 ));
    Odrv4 I__5685 (
            .O(N__27900),
            .I(\this_vga_signals.vaddress_7 ));
    LocalMux I__5684 (
            .O(N__27897),
            .I(\this_vga_signals.vaddress_7 ));
    LocalMux I__5683 (
            .O(N__27894),
            .I(\this_vga_signals.vaddress_7 ));
    InMux I__5682 (
            .O(N__27883),
            .I(N__27880));
    LocalMux I__5681 (
            .O(N__27880),
            .I(\this_vga_signals.N_38_i_0_a2_0_4Z0Z_1 ));
    CascadeMux I__5680 (
            .O(N__27877),
            .I(\this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_17_cascade_ ));
    InMux I__5679 (
            .O(N__27874),
            .I(N__27868));
    InMux I__5678 (
            .O(N__27873),
            .I(N__27865));
    InMux I__5677 (
            .O(N__27872),
            .I(N__27860));
    InMux I__5676 (
            .O(N__27871),
            .I(N__27860));
    LocalMux I__5675 (
            .O(N__27868),
            .I(M_this_state_qZ0Z_17));
    LocalMux I__5674 (
            .O(N__27865),
            .I(M_this_state_qZ0Z_17));
    LocalMux I__5673 (
            .O(N__27860),
            .I(M_this_state_qZ0Z_17));
    InMux I__5672 (
            .O(N__27853),
            .I(N__27850));
    LocalMux I__5671 (
            .O(N__27850),
            .I(N__27847));
    Odrv12 I__5670 (
            .O(N__27847),
            .I(\this_vga_signals.vsync_1_0_a3_0_a3_0 ));
    InMux I__5669 (
            .O(N__27844),
            .I(N__27841));
    LocalMux I__5668 (
            .O(N__27841),
            .I(\this_vga_signals.N_2840_0_0 ));
    InMux I__5667 (
            .O(N__27838),
            .I(N__27835));
    LocalMux I__5666 (
            .O(N__27835),
            .I(\this_vga_signals.N_27_0_0 ));
    CascadeMux I__5665 (
            .O(N__27832),
            .I(\this_vga_signals.vaddress_7_cascade_ ));
    InMux I__5664 (
            .O(N__27829),
            .I(N__27825));
    InMux I__5663 (
            .O(N__27828),
            .I(N__27822));
    LocalMux I__5662 (
            .O(N__27825),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    LocalMux I__5661 (
            .O(N__27822),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    InMux I__5660 (
            .O(N__27817),
            .I(N__27813));
    CascadeMux I__5659 (
            .O(N__27816),
            .I(N__27810));
    LocalMux I__5658 (
            .O(N__27813),
            .I(N__27807));
    InMux I__5657 (
            .O(N__27810),
            .I(N__27804));
    Odrv4 I__5656 (
            .O(N__27807),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__5655 (
            .O(N__27804),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    CascadeMux I__5654 (
            .O(N__27799),
            .I(\this_vga_signals.g1_2_0_cascade_ ));
    InMux I__5653 (
            .O(N__27796),
            .I(N__27793));
    LocalMux I__5652 (
            .O(N__27793),
            .I(N__27790));
    Odrv4 I__5651 (
            .O(N__27790),
            .I(\this_vga_signals.if_m6_i_x2_3 ));
    InMux I__5650 (
            .O(N__27787),
            .I(N__27784));
    LocalMux I__5649 (
            .O(N__27784),
            .I(\this_vga_signals.g1_3 ));
    CascadeMux I__5648 (
            .O(N__27781),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0_ns_1_cascade_ ));
    InMux I__5647 (
            .O(N__27778),
            .I(N__27775));
    LocalMux I__5646 (
            .O(N__27775),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_c_0_1 ));
    InMux I__5645 (
            .O(N__27772),
            .I(N__27769));
    LocalMux I__5644 (
            .O(N__27769),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_1_0 ));
    CascadeMux I__5643 (
            .O(N__27766),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_ ));
    InMux I__5642 (
            .O(N__27763),
            .I(N__27759));
    InMux I__5641 (
            .O(N__27762),
            .I(N__27756));
    LocalMux I__5640 (
            .O(N__27759),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_1_1 ));
    LocalMux I__5639 (
            .O(N__27756),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_1_1 ));
    CascadeMux I__5638 (
            .O(N__27751),
            .I(\this_vga_signals.if_m5_s_cascade_ ));
    CascadeMux I__5637 (
            .O(N__27748),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_1_0_cascade_ ));
    CascadeMux I__5636 (
            .O(N__27745),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ));
    InMux I__5635 (
            .O(N__27742),
            .I(N__27739));
    LocalMux I__5634 (
            .O(N__27739),
            .I(\this_vga_signals.if_m5_d ));
    CascadeMux I__5633 (
            .O(N__27736),
            .I(\this_vga_signals.if_m5_d_cascade_ ));
    InMux I__5632 (
            .O(N__27733),
            .I(N__27730));
    LocalMux I__5631 (
            .O(N__27730),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1 ));
    CascadeMux I__5630 (
            .O(N__27727),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1_cascade_ ));
    CascadeMux I__5629 (
            .O(N__27724),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_x0_cascade_ ));
    InMux I__5628 (
            .O(N__27721),
            .I(N__27718));
    LocalMux I__5627 (
            .O(N__27718),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_x1 ));
    InMux I__5626 (
            .O(N__27715),
            .I(N__27712));
    LocalMux I__5625 (
            .O(N__27712),
            .I(N__27709));
    Span4Mux_v I__5624 (
            .O(N__27709),
            .I(N__27705));
    InMux I__5623 (
            .O(N__27708),
            .I(N__27702));
    Span4Mux_h I__5622 (
            .O(N__27705),
            .I(N__27699));
    LocalMux I__5621 (
            .O(N__27702),
            .I(N__27696));
    Odrv4 I__5620 (
            .O(N__27699),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    Odrv12 I__5619 (
            .O(N__27696),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    CascadeMux I__5618 (
            .O(N__27691),
            .I(\this_vga_signals.N_38_i_0_a2_3_cascade_ ));
    InMux I__5617 (
            .O(N__27688),
            .I(N__27685));
    LocalMux I__5616 (
            .O(N__27685),
            .I(\this_vga_signals.N_38_i_0_a2_0_3 ));
    CascadeMux I__5615 (
            .O(N__27682),
            .I(N__27676));
    CascadeMux I__5614 (
            .O(N__27681),
            .I(N__27672));
    InMux I__5613 (
            .O(N__27680),
            .I(N__27667));
    InMux I__5612 (
            .O(N__27679),
            .I(N__27667));
    InMux I__5611 (
            .O(N__27676),
            .I(N__27664));
    InMux I__5610 (
            .O(N__27675),
            .I(N__27661));
    InMux I__5609 (
            .O(N__27672),
            .I(N__27658));
    LocalMux I__5608 (
            .O(N__27667),
            .I(N__27655));
    LocalMux I__5607 (
            .O(N__27664),
            .I(N__27652));
    LocalMux I__5606 (
            .O(N__27661),
            .I(N__27647));
    LocalMux I__5605 (
            .O(N__27658),
            .I(N__27647));
    Span4Mux_v I__5604 (
            .O(N__27655),
            .I(N__27642));
    Span4Mux_v I__5603 (
            .O(N__27652),
            .I(N__27642));
    Span4Mux_v I__5602 (
            .O(N__27647),
            .I(N__27639));
    Span4Mux_v I__5601 (
            .O(N__27642),
            .I(N__27636));
    Span4Mux_h I__5600 (
            .O(N__27639),
            .I(N__27633));
    Span4Mux_h I__5599 (
            .O(N__27636),
            .I(N__27630));
    Span4Mux_v I__5598 (
            .O(N__27633),
            .I(N__27627));
    Sp12to4 I__5597 (
            .O(N__27630),
            .I(N__27622));
    Sp12to4 I__5596 (
            .O(N__27627),
            .I(N__27622));
    Span12Mux_h I__5595 (
            .O(N__27622),
            .I(N__27619));
    Odrv12 I__5594 (
            .O(N__27619),
            .I(port_enb_c));
    InMux I__5593 (
            .O(N__27616),
            .I(N__27610));
    InMux I__5592 (
            .O(N__27615),
            .I(N__27607));
    InMux I__5591 (
            .O(N__27614),
            .I(N__27604));
    InMux I__5590 (
            .O(N__27613),
            .I(N__27601));
    LocalMux I__5589 (
            .O(N__27610),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__5588 (
            .O(N__27607),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__5587 (
            .O(N__27604),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__5586 (
            .O(N__27601),
            .I(this_start_data_delay_M_last_q));
    InMux I__5585 (
            .O(N__27592),
            .I(N__27589));
    LocalMux I__5584 (
            .O(N__27589),
            .I(N__27582));
    InMux I__5583 (
            .O(N__27588),
            .I(N__27577));
    InMux I__5582 (
            .O(N__27587),
            .I(N__27577));
    InMux I__5581 (
            .O(N__27586),
            .I(N__27572));
    InMux I__5580 (
            .O(N__27585),
            .I(N__27572));
    Odrv4 I__5579 (
            .O(N__27582),
            .I(M_this_delay_clk_out_0));
    LocalMux I__5578 (
            .O(N__27577),
            .I(M_this_delay_clk_out_0));
    LocalMux I__5577 (
            .O(N__27572),
            .I(M_this_delay_clk_out_0));
    CascadeMux I__5576 (
            .O(N__27565),
            .I(N_765_0_cascade_));
    InMux I__5575 (
            .O(N__27562),
            .I(N__27559));
    LocalMux I__5574 (
            .O(N__27559),
            .I(N__27556));
    Odrv4 I__5573 (
            .O(N__27556),
            .I(\this_ppu.N_229_1_0 ));
    CascadeMux I__5572 (
            .O(N__27553),
            .I(\this_ppu.N_229_1_0_cascade_ ));
    InMux I__5571 (
            .O(N__27550),
            .I(N__27532));
    InMux I__5570 (
            .O(N__27549),
            .I(N__27532));
    InMux I__5569 (
            .O(N__27548),
            .I(N__27521));
    InMux I__5568 (
            .O(N__27547),
            .I(N__27521));
    InMux I__5567 (
            .O(N__27546),
            .I(N__27521));
    InMux I__5566 (
            .O(N__27545),
            .I(N__27521));
    InMux I__5565 (
            .O(N__27544),
            .I(N__27521));
    InMux I__5564 (
            .O(N__27543),
            .I(N__27506));
    InMux I__5563 (
            .O(N__27542),
            .I(N__27506));
    InMux I__5562 (
            .O(N__27541),
            .I(N__27506));
    InMux I__5561 (
            .O(N__27540),
            .I(N__27506));
    InMux I__5560 (
            .O(N__27539),
            .I(N__27506));
    InMux I__5559 (
            .O(N__27538),
            .I(N__27506));
    InMux I__5558 (
            .O(N__27537),
            .I(N__27506));
    LocalMux I__5557 (
            .O(N__27532),
            .I(N__27501));
    LocalMux I__5556 (
            .O(N__27521),
            .I(N__27501));
    LocalMux I__5555 (
            .O(N__27506),
            .I(N__27498));
    Span4Mux_h I__5554 (
            .O(N__27501),
            .I(N__27495));
    Odrv4 I__5553 (
            .O(N__27498),
            .I(N_229));
    Odrv4 I__5552 (
            .O(N__27495),
            .I(N_229));
    CascadeMux I__5551 (
            .O(N__27490),
            .I(N__27486));
    InMux I__5550 (
            .O(N__27489),
            .I(N__27483));
    InMux I__5549 (
            .O(N__27486),
            .I(N__27477));
    LocalMux I__5548 (
            .O(N__27483),
            .I(N__27474));
    InMux I__5547 (
            .O(N__27482),
            .I(N__27467));
    InMux I__5546 (
            .O(N__27481),
            .I(N__27467));
    InMux I__5545 (
            .O(N__27480),
            .I(N__27467));
    LocalMux I__5544 (
            .O(N__27477),
            .I(N__27460));
    Span4Mux_h I__5543 (
            .O(N__27474),
            .I(N__27457));
    LocalMux I__5542 (
            .O(N__27467),
            .I(N__27454));
    InMux I__5541 (
            .O(N__27466),
            .I(N__27445));
    InMux I__5540 (
            .O(N__27465),
            .I(N__27445));
    InMux I__5539 (
            .O(N__27464),
            .I(N__27445));
    InMux I__5538 (
            .O(N__27463),
            .I(N__27445));
    Odrv12 I__5537 (
            .O(N__27460),
            .I(N_1423));
    Odrv4 I__5536 (
            .O(N__27457),
            .I(N_1423));
    Odrv4 I__5535 (
            .O(N__27454),
            .I(N_1423));
    LocalMux I__5534 (
            .O(N__27445),
            .I(N_1423));
    CascadeMux I__5533 (
            .O(N__27436),
            .I(\this_vga_signals.SUM_2_i_i_1_0_3_cascade_ ));
    InMux I__5532 (
            .O(N__27433),
            .I(N__27428));
    InMux I__5531 (
            .O(N__27432),
            .I(N__27422));
    InMux I__5530 (
            .O(N__27431),
            .I(N__27419));
    LocalMux I__5529 (
            .O(N__27428),
            .I(N__27416));
    InMux I__5528 (
            .O(N__27427),
            .I(N__27411));
    InMux I__5527 (
            .O(N__27426),
            .I(N__27411));
    InMux I__5526 (
            .O(N__27425),
            .I(N__27408));
    LocalMux I__5525 (
            .O(N__27422),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__5524 (
            .O(N__27419),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__5523 (
            .O(N__27416),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__5522 (
            .O(N__27411),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__5521 (
            .O(N__27408),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    InMux I__5520 (
            .O(N__27397),
            .I(N__27394));
    LocalMux I__5519 (
            .O(N__27394),
            .I(N__27391));
    Span4Mux_v I__5518 (
            .O(N__27391),
            .I(N__27388));
    Odrv4 I__5517 (
            .O(N__27388),
            .I(\this_vga_signals.vsync_1_0_a3_0_a3_5 ));
    InMux I__5516 (
            .O(N__27385),
            .I(N__27379));
    InMux I__5515 (
            .O(N__27384),
            .I(N__27376));
    InMux I__5514 (
            .O(N__27383),
            .I(N__27371));
    InMux I__5513 (
            .O(N__27382),
            .I(N__27371));
    LocalMux I__5512 (
            .O(N__27379),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__5511 (
            .O(N__27376),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__5510 (
            .O(N__27371),
            .I(M_this_state_qZ0Z_12));
    CascadeMux I__5509 (
            .O(N__27364),
            .I(\this_ppu.N_430_1_0_cascade_ ));
    InMux I__5508 (
            .O(N__27361),
            .I(N__27355));
    InMux I__5507 (
            .O(N__27360),
            .I(N__27355));
    LocalMux I__5506 (
            .O(N__27355),
            .I(M_this_state_q_fastZ0Z_13));
    CascadeMux I__5505 (
            .O(N__27352),
            .I(\this_vga_signals.N_38_i_0_a2_3Z0Z_0_cascade_ ));
    CascadeMux I__5504 (
            .O(N__27349),
            .I(\this_vga_signals.N_38_i_0_a2_3_xZ0Z1_cascade_ ));
    InMux I__5503 (
            .O(N__27346),
            .I(N__27336));
    InMux I__5502 (
            .O(N__27345),
            .I(N__27336));
    InMux I__5501 (
            .O(N__27344),
            .I(N__27336));
    InMux I__5500 (
            .O(N__27343),
            .I(N__27330));
    LocalMux I__5499 (
            .O(N__27336),
            .I(N__27323));
    CEMux I__5498 (
            .O(N__27335),
            .I(N__27320));
    InMux I__5497 (
            .O(N__27334),
            .I(N__27317));
    InMux I__5496 (
            .O(N__27333),
            .I(N__27314));
    LocalMux I__5495 (
            .O(N__27330),
            .I(N__27309));
    InMux I__5494 (
            .O(N__27329),
            .I(N__27304));
    InMux I__5493 (
            .O(N__27328),
            .I(N__27304));
    InMux I__5492 (
            .O(N__27327),
            .I(N__27299));
    InMux I__5491 (
            .O(N__27326),
            .I(N__27299));
    Span4Mux_v I__5490 (
            .O(N__27323),
            .I(N__27286));
    LocalMux I__5489 (
            .O(N__27320),
            .I(N__27286));
    LocalMux I__5488 (
            .O(N__27317),
            .I(N__27281));
    LocalMux I__5487 (
            .O(N__27314),
            .I(N__27281));
    InMux I__5486 (
            .O(N__27313),
            .I(N__27274));
    InMux I__5485 (
            .O(N__27312),
            .I(N__27274));
    Span12Mux_v I__5484 (
            .O(N__27309),
            .I(N__27271));
    LocalMux I__5483 (
            .O(N__27304),
            .I(N__27266));
    LocalMux I__5482 (
            .O(N__27299),
            .I(N__27266));
    InMux I__5481 (
            .O(N__27298),
            .I(N__27263));
    InMux I__5480 (
            .O(N__27297),
            .I(N__27260));
    InMux I__5479 (
            .O(N__27296),
            .I(N__27255));
    InMux I__5478 (
            .O(N__27295),
            .I(N__27255));
    InMux I__5477 (
            .O(N__27294),
            .I(N__27246));
    InMux I__5476 (
            .O(N__27293),
            .I(N__27246));
    InMux I__5475 (
            .O(N__27292),
            .I(N__27246));
    InMux I__5474 (
            .O(N__27291),
            .I(N__27246));
    Span4Mux_v I__5473 (
            .O(N__27286),
            .I(N__27243));
    Span4Mux_v I__5472 (
            .O(N__27281),
            .I(N__27240));
    InMux I__5471 (
            .O(N__27280),
            .I(N__27235));
    InMux I__5470 (
            .O(N__27279),
            .I(N__27235));
    LocalMux I__5469 (
            .O(N__27274),
            .I(N__27230));
    Span12Mux_h I__5468 (
            .O(N__27271),
            .I(N__27230));
    Span12Mux_v I__5467 (
            .O(N__27266),
            .I(N__27225));
    LocalMux I__5466 (
            .O(N__27263),
            .I(N__27225));
    LocalMux I__5465 (
            .O(N__27260),
            .I(G_535));
    LocalMux I__5464 (
            .O(N__27255),
            .I(G_535));
    LocalMux I__5463 (
            .O(N__27246),
            .I(G_535));
    Odrv4 I__5462 (
            .O(N__27243),
            .I(G_535));
    Odrv4 I__5461 (
            .O(N__27240),
            .I(G_535));
    LocalMux I__5460 (
            .O(N__27235),
            .I(G_535));
    Odrv12 I__5459 (
            .O(N__27230),
            .I(G_535));
    Odrv12 I__5458 (
            .O(N__27225),
            .I(G_535));
    InMux I__5457 (
            .O(N__27208),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__5456 (
            .O(N__27205),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__5455 (
            .O(N__27202),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__5454 (
            .O(N__27199),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__5453 (
            .O(N__27196),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    InMux I__5452 (
            .O(N__27193),
            .I(bfn_18_22_0_));
    InMux I__5451 (
            .O(N__27190),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    CascadeMux I__5450 (
            .O(N__27187),
            .I(N__27184));
    InMux I__5449 (
            .O(N__27184),
            .I(N__27181));
    LocalMux I__5448 (
            .O(N__27181),
            .I(N__27178));
    Span4Mux_v I__5447 (
            .O(N__27178),
            .I(N__27175));
    Odrv4 I__5446 (
            .O(N__27175),
            .I(\this_vga_signals.g0_0_0 ));
    InMux I__5445 (
            .O(N__27172),
            .I(N__27169));
    LocalMux I__5444 (
            .O(N__27169),
            .I(N__27166));
    Odrv12 I__5443 (
            .O(N__27166),
            .I(\this_vga_signals.IO_port_data_write_0_a2_i_o2_2Z0Z_1 ));
    CascadeMux I__5442 (
            .O(N__27163),
            .I(N__27160));
    InMux I__5441 (
            .O(N__27160),
            .I(N__27157));
    LocalMux I__5440 (
            .O(N__27157),
            .I(N__27154));
    Odrv4 I__5439 (
            .O(N__27154),
            .I(\this_vga_signals.mult1_un54_sum_2_1 ));
    InMux I__5438 (
            .O(N__27151),
            .I(N__27148));
    LocalMux I__5437 (
            .O(N__27148),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0 ));
    InMux I__5436 (
            .O(N__27145),
            .I(N__27142));
    LocalMux I__5435 (
            .O(N__27142),
            .I(\this_ppu.N_1115 ));
    CascadeMux I__5434 (
            .O(N__27139),
            .I(N__27136));
    InMux I__5433 (
            .O(N__27136),
            .I(N__27133));
    LocalMux I__5432 (
            .O(N__27133),
            .I(\this_vga_signals.g0_33_N_3L4 ));
    InMux I__5431 (
            .O(N__27130),
            .I(N__27127));
    LocalMux I__5430 (
            .O(N__27127),
            .I(\this_vga_signals.g0_33_N_4L6 ));
    InMux I__5429 (
            .O(N__27124),
            .I(N__27121));
    LocalMux I__5428 (
            .O(N__27121),
            .I(\this_vga_signals.g0_33_N_5L8 ));
    CascadeMux I__5427 (
            .O(N__27118),
            .I(N__27113));
    InMux I__5426 (
            .O(N__27117),
            .I(N__27110));
    InMux I__5425 (
            .O(N__27116),
            .I(N__27107));
    InMux I__5424 (
            .O(N__27113),
            .I(N__27104));
    LocalMux I__5423 (
            .O(N__27110),
            .I(N__27098));
    LocalMux I__5422 (
            .O(N__27107),
            .I(N__27095));
    LocalMux I__5421 (
            .O(N__27104),
            .I(N__27092));
    InMux I__5420 (
            .O(N__27103),
            .I(N__27089));
    InMux I__5419 (
            .O(N__27102),
            .I(N__27086));
    InMux I__5418 (
            .O(N__27101),
            .I(N__27083));
    Span4Mux_v I__5417 (
            .O(N__27098),
            .I(N__27075));
    Span4Mux_h I__5416 (
            .O(N__27095),
            .I(N__27075));
    Span4Mux_v I__5415 (
            .O(N__27092),
            .I(N__27075));
    LocalMux I__5414 (
            .O(N__27089),
            .I(N__27069));
    LocalMux I__5413 (
            .O(N__27086),
            .I(N__27069));
    LocalMux I__5412 (
            .O(N__27083),
            .I(N__27066));
    InMux I__5411 (
            .O(N__27082),
            .I(N__27063));
    Span4Mux_v I__5410 (
            .O(N__27075),
            .I(N__27058));
    InMux I__5409 (
            .O(N__27074),
            .I(N__27055));
    Span4Mux_h I__5408 (
            .O(N__27069),
            .I(N__27052));
    Span4Mux_v I__5407 (
            .O(N__27066),
            .I(N__27047));
    LocalMux I__5406 (
            .O(N__27063),
            .I(N__27047));
    InMux I__5405 (
            .O(N__27062),
            .I(N__27042));
    InMux I__5404 (
            .O(N__27061),
            .I(N__27042));
    Sp12to4 I__5403 (
            .O(N__27058),
            .I(N__27037));
    LocalMux I__5402 (
            .O(N__27055),
            .I(N__27037));
    Odrv4 I__5401 (
            .O(N__27052),
            .I(\this_vga_signals.M_hcounter_d7_0_i_0_0 ));
    Odrv4 I__5400 (
            .O(N__27047),
            .I(\this_vga_signals.M_hcounter_d7_0_i_0_0 ));
    LocalMux I__5399 (
            .O(N__27042),
            .I(\this_vga_signals.M_hcounter_d7_0_i_0_0 ));
    Odrv12 I__5398 (
            .O(N__27037),
            .I(\this_vga_signals.M_hcounter_d7_0_i_0_0 ));
    InMux I__5397 (
            .O(N__27028),
            .I(N__27023));
    InMux I__5396 (
            .O(N__27027),
            .I(N__27020));
    InMux I__5395 (
            .O(N__27026),
            .I(N__27017));
    LocalMux I__5394 (
            .O(N__27023),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__5393 (
            .O(N__27020),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__5392 (
            .O(N__27017),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    InMux I__5391 (
            .O(N__27010),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    InMux I__5390 (
            .O(N__27007),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__5389 (
            .O(N__27004),
            .I(N__27001));
    LocalMux I__5388 (
            .O(N__27001),
            .I(\this_vga_signals.mult1_un61_sum_axb2_i ));
    CascadeMux I__5387 (
            .O(N__26998),
            .I(N__26995));
    CascadeBuf I__5386 (
            .O(N__26995),
            .I(N__26992));
    CascadeMux I__5385 (
            .O(N__26992),
            .I(N__26989));
    InMux I__5384 (
            .O(N__26989),
            .I(N__26985));
    InMux I__5383 (
            .O(N__26988),
            .I(N__26982));
    LocalMux I__5382 (
            .O(N__26985),
            .I(N__26978));
    LocalMux I__5381 (
            .O(N__26982),
            .I(N__26974));
    CascadeMux I__5380 (
            .O(N__26981),
            .I(N__26971));
    Span4Mux_v I__5379 (
            .O(N__26978),
            .I(N__26967));
    InMux I__5378 (
            .O(N__26977),
            .I(N__26964));
    Span4Mux_h I__5377 (
            .O(N__26974),
            .I(N__26961));
    InMux I__5376 (
            .O(N__26971),
            .I(N__26956));
    InMux I__5375 (
            .O(N__26970),
            .I(N__26956));
    Sp12to4 I__5374 (
            .O(N__26967),
            .I(N__26953));
    LocalMux I__5373 (
            .O(N__26964),
            .I(M_this_oam_address_qZ0Z_3));
    Odrv4 I__5372 (
            .O(N__26961),
            .I(M_this_oam_address_qZ0Z_3));
    LocalMux I__5371 (
            .O(N__26956),
            .I(M_this_oam_address_qZ0Z_3));
    Odrv12 I__5370 (
            .O(N__26953),
            .I(M_this_oam_address_qZ0Z_3));
    InMux I__5369 (
            .O(N__26944),
            .I(N__26940));
    InMux I__5368 (
            .O(N__26943),
            .I(N__26937));
    LocalMux I__5367 (
            .O(N__26940),
            .I(un1_M_this_oam_address_q_c3));
    LocalMux I__5366 (
            .O(N__26937),
            .I(un1_M_this_oam_address_q_c3));
    CascadeMux I__5365 (
            .O(N__26932),
            .I(N__26929));
    CascadeBuf I__5364 (
            .O(N__26929),
            .I(N__26926));
    CascadeMux I__5363 (
            .O(N__26926),
            .I(N__26920));
    CascadeMux I__5362 (
            .O(N__26925),
            .I(N__26917));
    CascadeMux I__5361 (
            .O(N__26924),
            .I(N__26914));
    InMux I__5360 (
            .O(N__26923),
            .I(N__26911));
    InMux I__5359 (
            .O(N__26920),
            .I(N__26908));
    InMux I__5358 (
            .O(N__26917),
            .I(N__26905));
    InMux I__5357 (
            .O(N__26914),
            .I(N__26902));
    LocalMux I__5356 (
            .O(N__26911),
            .I(N__26897));
    LocalMux I__5355 (
            .O(N__26908),
            .I(N__26897));
    LocalMux I__5354 (
            .O(N__26905),
            .I(M_this_oam_address_qZ0Z_4));
    LocalMux I__5353 (
            .O(N__26902),
            .I(M_this_oam_address_qZ0Z_4));
    Odrv12 I__5352 (
            .O(N__26897),
            .I(M_this_oam_address_qZ0Z_4));
    CascadeMux I__5351 (
            .O(N__26890),
            .I(N__26884));
    CascadeMux I__5350 (
            .O(N__26889),
            .I(N__26881));
    CascadeMux I__5349 (
            .O(N__26888),
            .I(N__26877));
    InMux I__5348 (
            .O(N__26887),
            .I(N__26870));
    InMux I__5347 (
            .O(N__26884),
            .I(N__26870));
    InMux I__5346 (
            .O(N__26881),
            .I(N__26867));
    InMux I__5345 (
            .O(N__26880),
            .I(N__26860));
    InMux I__5344 (
            .O(N__26877),
            .I(N__26860));
    InMux I__5343 (
            .O(N__26876),
            .I(N__26860));
    InMux I__5342 (
            .O(N__26875),
            .I(N__26857));
    LocalMux I__5341 (
            .O(N__26870),
            .I(N__26854));
    LocalMux I__5340 (
            .O(N__26867),
            .I(M_this_oam_address_qZ0Z_1));
    LocalMux I__5339 (
            .O(N__26860),
            .I(M_this_oam_address_qZ0Z_1));
    LocalMux I__5338 (
            .O(N__26857),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__5337 (
            .O(N__26854),
            .I(M_this_oam_address_qZ0Z_1));
    InMux I__5336 (
            .O(N__26845),
            .I(N__26835));
    InMux I__5335 (
            .O(N__26844),
            .I(N__26830));
    InMux I__5334 (
            .O(N__26843),
            .I(N__26830));
    InMux I__5333 (
            .O(N__26842),
            .I(N__26827));
    InMux I__5332 (
            .O(N__26841),
            .I(N__26824));
    InMux I__5331 (
            .O(N__26840),
            .I(N__26819));
    InMux I__5330 (
            .O(N__26839),
            .I(N__26819));
    InMux I__5329 (
            .O(N__26838),
            .I(N__26816));
    LocalMux I__5328 (
            .O(N__26835),
            .I(N__26813));
    LocalMux I__5327 (
            .O(N__26830),
            .I(N__26810));
    LocalMux I__5326 (
            .O(N__26827),
            .I(M_this_oam_address_qZ0Z_0));
    LocalMux I__5325 (
            .O(N__26824),
            .I(M_this_oam_address_qZ0Z_0));
    LocalMux I__5324 (
            .O(N__26819),
            .I(M_this_oam_address_qZ0Z_0));
    LocalMux I__5323 (
            .O(N__26816),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__5322 (
            .O(N__26813),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__5321 (
            .O(N__26810),
            .I(M_this_oam_address_qZ0Z_0));
    CascadeMux I__5320 (
            .O(N__26797),
            .I(N__26793));
    InMux I__5319 (
            .O(N__26796),
            .I(N__26786));
    InMux I__5318 (
            .O(N__26793),
            .I(N__26779));
    InMux I__5317 (
            .O(N__26792),
            .I(N__26779));
    InMux I__5316 (
            .O(N__26791),
            .I(N__26779));
    InMux I__5315 (
            .O(N__26790),
            .I(N__26776));
    InMux I__5314 (
            .O(N__26789),
            .I(N__26773));
    LocalMux I__5313 (
            .O(N__26786),
            .I(N__26766));
    LocalMux I__5312 (
            .O(N__26779),
            .I(N__26766));
    LocalMux I__5311 (
            .O(N__26776),
            .I(N__26766));
    LocalMux I__5310 (
            .O(N__26773),
            .I(N_778_0));
    Odrv4 I__5309 (
            .O(N__26766),
            .I(N_778_0));
    InMux I__5308 (
            .O(N__26761),
            .I(N__26754));
    InMux I__5307 (
            .O(N__26760),
            .I(N__26749));
    InMux I__5306 (
            .O(N__26759),
            .I(N__26749));
    CEMux I__5305 (
            .O(N__26758),
            .I(N__26744));
    CEMux I__5304 (
            .O(N__26757),
            .I(N__26741));
    LocalMux I__5303 (
            .O(N__26754),
            .I(N__26713));
    LocalMux I__5302 (
            .O(N__26749),
            .I(N__26713));
    InMux I__5301 (
            .O(N__26748),
            .I(N__26708));
    InMux I__5300 (
            .O(N__26747),
            .I(N__26708));
    LocalMux I__5299 (
            .O(N__26744),
            .I(N__26703));
    LocalMux I__5298 (
            .O(N__26741),
            .I(N__26703));
    InMux I__5297 (
            .O(N__26740),
            .I(N__26698));
    InMux I__5296 (
            .O(N__26739),
            .I(N__26698));
    InMux I__5295 (
            .O(N__26738),
            .I(N__26689));
    InMux I__5294 (
            .O(N__26737),
            .I(N__26689));
    InMux I__5293 (
            .O(N__26736),
            .I(N__26689));
    InMux I__5292 (
            .O(N__26735),
            .I(N__26689));
    InMux I__5291 (
            .O(N__26734),
            .I(N__26680));
    InMux I__5290 (
            .O(N__26733),
            .I(N__26680));
    InMux I__5289 (
            .O(N__26732),
            .I(N__26680));
    InMux I__5288 (
            .O(N__26731),
            .I(N__26680));
    InMux I__5287 (
            .O(N__26730),
            .I(N__26675));
    InMux I__5286 (
            .O(N__26729),
            .I(N__26675));
    InMux I__5285 (
            .O(N__26728),
            .I(N__26667));
    InMux I__5284 (
            .O(N__26727),
            .I(N__26667));
    InMux I__5283 (
            .O(N__26726),
            .I(N__26667));
    InMux I__5282 (
            .O(N__26725),
            .I(N__26658));
    InMux I__5281 (
            .O(N__26724),
            .I(N__26658));
    InMux I__5280 (
            .O(N__26723),
            .I(N__26658));
    InMux I__5279 (
            .O(N__26722),
            .I(N__26658));
    InMux I__5278 (
            .O(N__26721),
            .I(N__26649));
    InMux I__5277 (
            .O(N__26720),
            .I(N__26649));
    InMux I__5276 (
            .O(N__26719),
            .I(N__26649));
    InMux I__5275 (
            .O(N__26718),
            .I(N__26649));
    Span4Mux_h I__5274 (
            .O(N__26713),
            .I(N__26644));
    LocalMux I__5273 (
            .O(N__26708),
            .I(N__26644));
    Span4Mux_v I__5272 (
            .O(N__26703),
            .I(N__26638));
    LocalMux I__5271 (
            .O(N__26698),
            .I(N__26633));
    LocalMux I__5270 (
            .O(N__26689),
            .I(N__26633));
    LocalMux I__5269 (
            .O(N__26680),
            .I(N__26628));
    LocalMux I__5268 (
            .O(N__26675),
            .I(N__26628));
    InMux I__5267 (
            .O(N__26674),
            .I(N__26625));
    LocalMux I__5266 (
            .O(N__26667),
            .I(N__26618));
    LocalMux I__5265 (
            .O(N__26658),
            .I(N__26618));
    LocalMux I__5264 (
            .O(N__26649),
            .I(N__26618));
    Span4Mux_v I__5263 (
            .O(N__26644),
            .I(N__26615));
    InMux I__5262 (
            .O(N__26643),
            .I(N__26612));
    InMux I__5261 (
            .O(N__26642),
            .I(N__26609));
    InMux I__5260 (
            .O(N__26641),
            .I(N__26606));
    Span4Mux_h I__5259 (
            .O(N__26638),
            .I(N__26599));
    Span4Mux_v I__5258 (
            .O(N__26633),
            .I(N__26599));
    Span4Mux_h I__5257 (
            .O(N__26628),
            .I(N__26599));
    LocalMux I__5256 (
            .O(N__26625),
            .I(N__26594));
    Span4Mux_h I__5255 (
            .O(N__26618),
            .I(N__26594));
    Sp12to4 I__5254 (
            .O(N__26615),
            .I(N__26585));
    LocalMux I__5253 (
            .O(N__26612),
            .I(N__26585));
    LocalMux I__5252 (
            .O(N__26609),
            .I(N__26585));
    LocalMux I__5251 (
            .O(N__26606),
            .I(N__26585));
    Span4Mux_h I__5250 (
            .O(N__26599),
            .I(N__26582));
    Span4Mux_h I__5249 (
            .O(N__26594),
            .I(N__26579));
    Odrv12 I__5248 (
            .O(N__26585),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    Odrv4 I__5247 (
            .O(N__26582),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    Odrv4 I__5246 (
            .O(N__26579),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    CascadeMux I__5245 (
            .O(N__26572),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_ ));
    CascadeMux I__5244 (
            .O(N__26569),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_0_1_cascade_ ));
    CascadeMux I__5243 (
            .O(N__26566),
            .I(N_778_0_cascade_));
    CEMux I__5242 (
            .O(N__26563),
            .I(N__26560));
    LocalMux I__5241 (
            .O(N__26560),
            .I(N__26555));
    CEMux I__5240 (
            .O(N__26559),
            .I(N__26552));
    CEMux I__5239 (
            .O(N__26558),
            .I(N__26549));
    Span4Mux_h I__5238 (
            .O(N__26555),
            .I(N__26544));
    LocalMux I__5237 (
            .O(N__26552),
            .I(N__26544));
    LocalMux I__5236 (
            .O(N__26549),
            .I(N__26541));
    Span4Mux_h I__5235 (
            .O(N__26544),
            .I(N__26538));
    Span4Mux_h I__5234 (
            .O(N__26541),
            .I(N__26535));
    Span4Mux_v I__5233 (
            .O(N__26538),
            .I(N__26532));
    Odrv4 I__5232 (
            .O(N__26535),
            .I(N_1701_0));
    Odrv4 I__5231 (
            .O(N__26532),
            .I(N_1701_0));
    InMux I__5230 (
            .O(N__26527),
            .I(N__26524));
    LocalMux I__5229 (
            .O(N__26524),
            .I(un1_M_this_oam_address_q_c5));
    CascadeMux I__5228 (
            .O(N__26521),
            .I(N__26518));
    CascadeBuf I__5227 (
            .O(N__26518),
            .I(N__26515));
    CascadeMux I__5226 (
            .O(N__26515),
            .I(N__26511));
    CascadeMux I__5225 (
            .O(N__26514),
            .I(N__26508));
    InMux I__5224 (
            .O(N__26511),
            .I(N__26505));
    InMux I__5223 (
            .O(N__26508),
            .I(N__26502));
    LocalMux I__5222 (
            .O(N__26505),
            .I(N__26499));
    LocalMux I__5221 (
            .O(N__26502),
            .I(N__26494));
    Sp12to4 I__5220 (
            .O(N__26499),
            .I(N__26491));
    InMux I__5219 (
            .O(N__26498),
            .I(N__26486));
    InMux I__5218 (
            .O(N__26497),
            .I(N__26486));
    Span4Mux_v I__5217 (
            .O(N__26494),
            .I(N__26483));
    Span12Mux_s7_v I__5216 (
            .O(N__26491),
            .I(N__26480));
    LocalMux I__5215 (
            .O(N__26486),
            .I(M_this_oam_address_qZ0Z_5));
    Odrv4 I__5214 (
            .O(N__26483),
            .I(M_this_oam_address_qZ0Z_5));
    Odrv12 I__5213 (
            .O(N__26480),
            .I(M_this_oam_address_qZ0Z_5));
    CascadeMux I__5212 (
            .O(N__26473),
            .I(un1_M_this_oam_address_q_c5_cascade_));
    CascadeMux I__5211 (
            .O(N__26470),
            .I(N__26467));
    CascadeBuf I__5210 (
            .O(N__26467),
            .I(N__26464));
    CascadeMux I__5209 (
            .O(N__26464),
            .I(N__26461));
    InMux I__5208 (
            .O(N__26461),
            .I(N__26458));
    LocalMux I__5207 (
            .O(N__26458),
            .I(N__26454));
    InMux I__5206 (
            .O(N__26457),
            .I(N__26451));
    Span4Mux_h I__5205 (
            .O(N__26454),
            .I(N__26448));
    LocalMux I__5204 (
            .O(N__26451),
            .I(N__26442));
    Span4Mux_h I__5203 (
            .O(N__26448),
            .I(N__26442));
    InMux I__5202 (
            .O(N__26447),
            .I(N__26439));
    Span4Mux_h I__5201 (
            .O(N__26442),
            .I(N__26436));
    LocalMux I__5200 (
            .O(N__26439),
            .I(M_this_oam_address_qZ0Z_6));
    Odrv4 I__5199 (
            .O(N__26436),
            .I(M_this_oam_address_qZ0Z_6));
    InMux I__5198 (
            .O(N__26431),
            .I(N__26428));
    LocalMux I__5197 (
            .O(N__26428),
            .I(N__26423));
    InMux I__5196 (
            .O(N__26427),
            .I(N__26418));
    InMux I__5195 (
            .O(N__26426),
            .I(N__26418));
    Odrv4 I__5194 (
            .O(N__26423),
            .I(un1_M_this_oam_address_q_c2));
    LocalMux I__5193 (
            .O(N__26418),
            .I(un1_M_this_oam_address_q_c2));
    CascadeMux I__5192 (
            .O(N__26413),
            .I(N__26410));
    CascadeBuf I__5191 (
            .O(N__26410),
            .I(N__26407));
    CascadeMux I__5190 (
            .O(N__26407),
            .I(N__26404));
    InMux I__5189 (
            .O(N__26404),
            .I(N__26400));
    CascadeMux I__5188 (
            .O(N__26403),
            .I(N__26394));
    LocalMux I__5187 (
            .O(N__26400),
            .I(N__26391));
    InMux I__5186 (
            .O(N__26399),
            .I(N__26388));
    InMux I__5185 (
            .O(N__26398),
            .I(N__26383));
    InMux I__5184 (
            .O(N__26397),
            .I(N__26383));
    InMux I__5183 (
            .O(N__26394),
            .I(N__26380));
    Span12Mux_s8_h I__5182 (
            .O(N__26391),
            .I(N__26377));
    LocalMux I__5181 (
            .O(N__26388),
            .I(M_this_oam_address_qZ0Z_2));
    LocalMux I__5180 (
            .O(N__26383),
            .I(M_this_oam_address_qZ0Z_2));
    LocalMux I__5179 (
            .O(N__26380),
            .I(M_this_oam_address_qZ0Z_2));
    Odrv12 I__5178 (
            .O(N__26377),
            .I(M_this_oam_address_qZ0Z_2));
    InMux I__5177 (
            .O(N__26368),
            .I(N__26364));
    InMux I__5176 (
            .O(N__26367),
            .I(N__26361));
    LocalMux I__5175 (
            .O(N__26364),
            .I(N__26358));
    LocalMux I__5174 (
            .O(N__26361),
            .I(N__26354));
    Span4Mux_h I__5173 (
            .O(N__26358),
            .I(N__26351));
    InMux I__5172 (
            .O(N__26357),
            .I(N__26348));
    Odrv12 I__5171 (
            .O(N__26354),
            .I(N_782_0));
    Odrv4 I__5170 (
            .O(N__26351),
            .I(N_782_0));
    LocalMux I__5169 (
            .O(N__26348),
            .I(N_782_0));
    CEMux I__5168 (
            .O(N__26341),
            .I(N__26338));
    LocalMux I__5167 (
            .O(N__26338),
            .I(N__26335));
    Span4Mux_h I__5166 (
            .O(N__26335),
            .I(N__26332));
    Span4Mux_h I__5165 (
            .O(N__26332),
            .I(N__26329));
    Odrv4 I__5164 (
            .O(N__26329),
            .I(N_1725_0));
    CEMux I__5163 (
            .O(N__26326),
            .I(N__26323));
    LocalMux I__5162 (
            .O(N__26323),
            .I(N__26320));
    Span4Mux_v I__5161 (
            .O(N__26320),
            .I(N__26317));
    Odrv4 I__5160 (
            .O(N__26317),
            .I(N_1717_0));
    InMux I__5159 (
            .O(N__26314),
            .I(N__26311));
    LocalMux I__5158 (
            .O(N__26311),
            .I(N__26308));
    Odrv4 I__5157 (
            .O(N__26308),
            .I(\this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_12 ));
    InMux I__5156 (
            .O(N__26305),
            .I(N__26302));
    LocalMux I__5155 (
            .O(N__26302),
            .I(N__26299));
    Span4Mux_h I__5154 (
            .O(N__26299),
            .I(N__26296));
    Span4Mux_h I__5153 (
            .O(N__26296),
            .I(N__26293));
    Odrv4 I__5152 (
            .O(N__26293),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    InMux I__5151 (
            .O(N__26290),
            .I(N__26287));
    LocalMux I__5150 (
            .O(N__26287),
            .I(N__26284));
    Span4Mux_h I__5149 (
            .O(N__26284),
            .I(N__26280));
    InMux I__5148 (
            .O(N__26283),
            .I(N__26277));
    Odrv4 I__5147 (
            .O(N__26280),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_16 ));
    LocalMux I__5146 (
            .O(N__26277),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_16 ));
    CascadeMux I__5145 (
            .O(N__26272),
            .I(N__26269));
    InMux I__5144 (
            .O(N__26269),
            .I(N__26266));
    LocalMux I__5143 (
            .O(N__26266),
            .I(N__26262));
    InMux I__5142 (
            .O(N__26265),
            .I(N__26259));
    Odrv4 I__5141 (
            .O(N__26262),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_16 ));
    LocalMux I__5140 (
            .O(N__26259),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_16 ));
    InMux I__5139 (
            .O(N__26254),
            .I(N__26250));
    InMux I__5138 (
            .O(N__26253),
            .I(N__26247));
    LocalMux I__5137 (
            .O(N__26250),
            .I(N__26244));
    LocalMux I__5136 (
            .O(N__26247),
            .I(N__26241));
    Odrv4 I__5135 (
            .O(N__26244),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_10Z0Z_16 ));
    Odrv4 I__5134 (
            .O(N__26241),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_10Z0Z_16 ));
    CascadeMux I__5133 (
            .O(N__26236),
            .I(N__26232));
    CascadeMux I__5132 (
            .O(N__26235),
            .I(N__26229));
    InMux I__5131 (
            .O(N__26232),
            .I(N__26225));
    InMux I__5130 (
            .O(N__26229),
            .I(N__26222));
    CascadeMux I__5129 (
            .O(N__26228),
            .I(N__26219));
    LocalMux I__5128 (
            .O(N__26225),
            .I(N__26216));
    LocalMux I__5127 (
            .O(N__26222),
            .I(N__26213));
    InMux I__5126 (
            .O(N__26219),
            .I(N__26210));
    Odrv12 I__5125 (
            .O(N__26216),
            .I(N_771_0));
    Odrv12 I__5124 (
            .O(N__26213),
            .I(N_771_0));
    LocalMux I__5123 (
            .O(N__26210),
            .I(N_771_0));
    CascadeMux I__5122 (
            .O(N__26203),
            .I(N_771_0_cascade_));
    InMux I__5121 (
            .O(N__26200),
            .I(N__26196));
    InMux I__5120 (
            .O(N__26199),
            .I(N__26193));
    LocalMux I__5119 (
            .O(N__26196),
            .I(N__26190));
    LocalMux I__5118 (
            .O(N__26193),
            .I(N__26187));
    Span4Mux_h I__5117 (
            .O(N__26190),
            .I(N__26184));
    Span4Mux_v I__5116 (
            .O(N__26187),
            .I(N__26181));
    Span4Mux_h I__5115 (
            .O(N__26184),
            .I(N__26178));
    Odrv4 I__5114 (
            .O(N__26181),
            .I(\this_ppu.N_774_0 ));
    Odrv4 I__5113 (
            .O(N__26178),
            .I(\this_ppu.N_774_0 ));
    CascadeMux I__5112 (
            .O(N__26173),
            .I(\this_vga_signals.g1_0_0_cascade_ ));
    InMux I__5111 (
            .O(N__26170),
            .I(N__26167));
    LocalMux I__5110 (
            .O(N__26167),
            .I(\this_vga_signals.if_N_6_0_0_0 ));
    CascadeMux I__5109 (
            .O(N__26164),
            .I(N__26161));
    InMux I__5108 (
            .O(N__26161),
            .I(N__26158));
    LocalMux I__5107 (
            .O(N__26158),
            .I(\this_vga_signals.g1_0_0 ));
    CascadeMux I__5106 (
            .O(N__26155),
            .I(\this_vga_signals.N_27_0_1_0_cascade_ ));
    InMux I__5105 (
            .O(N__26152),
            .I(N__26149));
    LocalMux I__5104 (
            .O(N__26149),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0 ));
    CascadeMux I__5103 (
            .O(N__26146),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_1_0_cascade_ ));
    CascadeMux I__5102 (
            .O(N__26143),
            .I(N__26138));
    CascadeMux I__5101 (
            .O(N__26142),
            .I(N__26132));
    CascadeMux I__5100 (
            .O(N__26141),
            .I(N__26125));
    InMux I__5099 (
            .O(N__26138),
            .I(N__26122));
    InMux I__5098 (
            .O(N__26137),
            .I(N__26119));
    InMux I__5097 (
            .O(N__26136),
            .I(N__26112));
    InMux I__5096 (
            .O(N__26135),
            .I(N__26109));
    InMux I__5095 (
            .O(N__26132),
            .I(N__26106));
    InMux I__5094 (
            .O(N__26131),
            .I(N__26103));
    InMux I__5093 (
            .O(N__26130),
            .I(N__26098));
    InMux I__5092 (
            .O(N__26129),
            .I(N__26098));
    InMux I__5091 (
            .O(N__26128),
            .I(N__26093));
    InMux I__5090 (
            .O(N__26125),
            .I(N__26093));
    LocalMux I__5089 (
            .O(N__26122),
            .I(N__26090));
    LocalMux I__5088 (
            .O(N__26119),
            .I(N__26087));
    InMux I__5087 (
            .O(N__26118),
            .I(N__26081));
    InMux I__5086 (
            .O(N__26117),
            .I(N__26081));
    IoInMux I__5085 (
            .O(N__26116),
            .I(N__26078));
    InMux I__5084 (
            .O(N__26115),
            .I(N__26070));
    LocalMux I__5083 (
            .O(N__26112),
            .I(N__26067));
    LocalMux I__5082 (
            .O(N__26109),
            .I(N__26064));
    LocalMux I__5081 (
            .O(N__26106),
            .I(N__26051));
    LocalMux I__5080 (
            .O(N__26103),
            .I(N__26051));
    LocalMux I__5079 (
            .O(N__26098),
            .I(N__26051));
    LocalMux I__5078 (
            .O(N__26093),
            .I(N__26051));
    Span4Mux_h I__5077 (
            .O(N__26090),
            .I(N__26051));
    Span4Mux_v I__5076 (
            .O(N__26087),
            .I(N__26051));
    InMux I__5075 (
            .O(N__26086),
            .I(N__26048));
    LocalMux I__5074 (
            .O(N__26081),
            .I(N__26045));
    LocalMux I__5073 (
            .O(N__26078),
            .I(N__26042));
    InMux I__5072 (
            .O(N__26077),
            .I(N__26039));
    InMux I__5071 (
            .O(N__26076),
            .I(N__26036));
    InMux I__5070 (
            .O(N__26075),
            .I(N__26033));
    InMux I__5069 (
            .O(N__26074),
            .I(N__26028));
    InMux I__5068 (
            .O(N__26073),
            .I(N__26028));
    LocalMux I__5067 (
            .O(N__26070),
            .I(N__26025));
    Span4Mux_v I__5066 (
            .O(N__26067),
            .I(N__26018));
    Span4Mux_v I__5065 (
            .O(N__26064),
            .I(N__26018));
    Span4Mux_v I__5064 (
            .O(N__26051),
            .I(N__26018));
    LocalMux I__5063 (
            .O(N__26048),
            .I(N__26013));
    Span4Mux_h I__5062 (
            .O(N__26045),
            .I(N__26013));
    Span12Mux_s6_h I__5061 (
            .O(N__26042),
            .I(N__26010));
    LocalMux I__5060 (
            .O(N__26039),
            .I(M_this_reset_cond_out_0));
    LocalMux I__5059 (
            .O(N__26036),
            .I(M_this_reset_cond_out_0));
    LocalMux I__5058 (
            .O(N__26033),
            .I(M_this_reset_cond_out_0));
    LocalMux I__5057 (
            .O(N__26028),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__5056 (
            .O(N__26025),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__5055 (
            .O(N__26018),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__5054 (
            .O(N__26013),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__5053 (
            .O(N__26010),
            .I(M_this_reset_cond_out_0));
    CascadeMux I__5052 (
            .O(N__25993),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_2_cascade_ ));
    CascadeMux I__5051 (
            .O(N__25990),
            .I(N__25987));
    InMux I__5050 (
            .O(N__25987),
            .I(N__25984));
    LocalMux I__5049 (
            .O(N__25984),
            .I(\this_vga_signals.N_4_0 ));
    InMux I__5048 (
            .O(N__25981),
            .I(N__25978));
    LocalMux I__5047 (
            .O(N__25978),
            .I(\this_vga_signals.if_m1_0_x2_1 ));
    InMux I__5046 (
            .O(N__25975),
            .I(N__25972));
    LocalMux I__5045 (
            .O(N__25972),
            .I(\this_vga_signals.r_N_2_i_0 ));
    CascadeMux I__5044 (
            .O(N__25969),
            .I(N__25965));
    InMux I__5043 (
            .O(N__25968),
            .I(N__25962));
    InMux I__5042 (
            .O(N__25965),
            .I(N__25958));
    LocalMux I__5041 (
            .O(N__25962),
            .I(N__25955));
    InMux I__5040 (
            .O(N__25961),
            .I(N__25952));
    LocalMux I__5039 (
            .O(N__25958),
            .I(N__25949));
    Odrv4 I__5038 (
            .O(N__25955),
            .I(\this_vga_signals.N_836_0 ));
    LocalMux I__5037 (
            .O(N__25952),
            .I(\this_vga_signals.N_836_0 ));
    Odrv12 I__5036 (
            .O(N__25949),
            .I(\this_vga_signals.N_836_0 ));
    CascadeMux I__5035 (
            .O(N__25942),
            .I(\this_vga_signals.N_1043_cascade_ ));
    InMux I__5034 (
            .O(N__25939),
            .I(N__25933));
    InMux I__5033 (
            .O(N__25938),
            .I(N__25933));
    LocalMux I__5032 (
            .O(N__25933),
            .I(N__25928));
    InMux I__5031 (
            .O(N__25932),
            .I(N__25923));
    InMux I__5030 (
            .O(N__25931),
            .I(N__25923));
    Odrv4 I__5029 (
            .O(N__25928),
            .I(this_vga_signals_M_lcounter_q_0));
    LocalMux I__5028 (
            .O(N__25923),
            .I(this_vga_signals_M_lcounter_q_0));
    InMux I__5027 (
            .O(N__25918),
            .I(N__25913));
    InMux I__5026 (
            .O(N__25917),
            .I(N__25910));
    InMux I__5025 (
            .O(N__25916),
            .I(N__25907));
    LocalMux I__5024 (
            .O(N__25913),
            .I(N__25899));
    LocalMux I__5023 (
            .O(N__25910),
            .I(N__25899));
    LocalMux I__5022 (
            .O(N__25907),
            .I(N__25899));
    InMux I__5021 (
            .O(N__25906),
            .I(N__25896));
    Odrv12 I__5020 (
            .O(N__25899),
            .I(N_792_0));
    LocalMux I__5019 (
            .O(N__25896),
            .I(N_792_0));
    CascadeMux I__5018 (
            .O(N__25891),
            .I(N__25888));
    InMux I__5017 (
            .O(N__25888),
            .I(N__25880));
    InMux I__5016 (
            .O(N__25887),
            .I(N__25880));
    CascadeMux I__5015 (
            .O(N__25886),
            .I(N__25876));
    CascadeMux I__5014 (
            .O(N__25885),
            .I(N__25873));
    LocalMux I__5013 (
            .O(N__25880),
            .I(N__25870));
    InMux I__5012 (
            .O(N__25879),
            .I(N__25863));
    InMux I__5011 (
            .O(N__25876),
            .I(N__25863));
    InMux I__5010 (
            .O(N__25873),
            .I(N__25863));
    Span4Mux_v I__5009 (
            .O(N__25870),
            .I(N__25860));
    LocalMux I__5008 (
            .O(N__25863),
            .I(this_vga_signals_M_lcounter_q_1));
    Odrv4 I__5007 (
            .O(N__25860),
            .I(this_vga_signals_M_lcounter_q_1));
    InMux I__5006 (
            .O(N__25855),
            .I(N__25852));
    LocalMux I__5005 (
            .O(N__25852),
            .I(N__25849));
    Odrv4 I__5004 (
            .O(N__25849),
            .I(\this_ppu.M_last_q_0 ));
    InMux I__5003 (
            .O(N__25846),
            .I(N__25843));
    LocalMux I__5002 (
            .O(N__25843),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x1 ));
    CascadeMux I__5001 (
            .O(N__25840),
            .I(N__25837));
    InMux I__5000 (
            .O(N__25837),
            .I(N__25834));
    LocalMux I__4999 (
            .O(N__25834),
            .I(M_this_scroll_qZ0Z_10));
    InMux I__4998 (
            .O(N__25831),
            .I(N__25828));
    LocalMux I__4997 (
            .O(N__25828),
            .I(N__25825));
    Odrv12 I__4996 (
            .O(N__25825),
            .I(M_this_scroll_qZ0Z_11));
    CascadeMux I__4995 (
            .O(N__25822),
            .I(N__25819));
    InMux I__4994 (
            .O(N__25819),
            .I(N__25816));
    LocalMux I__4993 (
            .O(N__25816),
            .I(N__25813));
    Span4Mux_v I__4992 (
            .O(N__25813),
            .I(N__25810));
    Span4Mux_h I__4991 (
            .O(N__25810),
            .I(N__25807));
    Odrv4 I__4990 (
            .O(N__25807),
            .I(M_this_scroll_qZ0Z_12));
    InMux I__4989 (
            .O(N__25804),
            .I(N__25801));
    LocalMux I__4988 (
            .O(N__25801),
            .I(N__25798));
    Odrv4 I__4987 (
            .O(N__25798),
            .I(M_this_scroll_qZ0Z_13));
    CascadeMux I__4986 (
            .O(N__25795),
            .I(N__25792));
    InMux I__4985 (
            .O(N__25792),
            .I(N__25789));
    LocalMux I__4984 (
            .O(N__25789),
            .I(N__25786));
    Span4Mux_h I__4983 (
            .O(N__25786),
            .I(N__25783));
    Odrv4 I__4982 (
            .O(N__25783),
            .I(M_this_scroll_qZ0Z_14));
    CascadeMux I__4981 (
            .O(N__25780),
            .I(N__25777));
    InMux I__4980 (
            .O(N__25777),
            .I(N__25774));
    LocalMux I__4979 (
            .O(N__25774),
            .I(N__25771));
    Span4Mux_h I__4978 (
            .O(N__25771),
            .I(N__25768));
    Odrv4 I__4977 (
            .O(N__25768),
            .I(M_this_scroll_qZ0Z_15));
    CascadeMux I__4976 (
            .O(N__25765),
            .I(N__25762));
    InMux I__4975 (
            .O(N__25762),
            .I(N__25759));
    LocalMux I__4974 (
            .O(N__25759),
            .I(N__25756));
    Odrv4 I__4973 (
            .O(N__25756),
            .I(M_this_scroll_qZ0Z_8));
    InMux I__4972 (
            .O(N__25753),
            .I(N__25750));
    LocalMux I__4971 (
            .O(N__25750),
            .I(N__25747));
    Span4Mux_h I__4970 (
            .O(N__25747),
            .I(N__25744));
    Odrv4 I__4969 (
            .O(N__25744),
            .I(M_this_scroll_qZ0Z_9));
    InMux I__4968 (
            .O(N__25741),
            .I(N__25738));
    LocalMux I__4967 (
            .O(N__25738),
            .I(N__25734));
    InMux I__4966 (
            .O(N__25737),
            .I(N__25730));
    Span4Mux_v I__4965 (
            .O(N__25734),
            .I(N__25727));
    InMux I__4964 (
            .O(N__25733),
            .I(N__25724));
    LocalMux I__4963 (
            .O(N__25730),
            .I(M_this_data_count_qZ0Z_7));
    Odrv4 I__4962 (
            .O(N__25727),
            .I(M_this_data_count_qZ0Z_7));
    LocalMux I__4961 (
            .O(N__25724),
            .I(M_this_data_count_qZ0Z_7));
    CascadeMux I__4960 (
            .O(N__25717),
            .I(N__25712));
    InMux I__4959 (
            .O(N__25716),
            .I(N__25709));
    InMux I__4958 (
            .O(N__25715),
            .I(N__25706));
    InMux I__4957 (
            .O(N__25712),
            .I(N__25703));
    LocalMux I__4956 (
            .O(N__25709),
            .I(N__25700));
    LocalMux I__4955 (
            .O(N__25706),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__4954 (
            .O(N__25703),
            .I(M_this_data_count_qZ0Z_6));
    Odrv4 I__4953 (
            .O(N__25700),
            .I(M_this_data_count_qZ0Z_6));
    InMux I__4952 (
            .O(N__25693),
            .I(N__25690));
    LocalMux I__4951 (
            .O(N__25690),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_16 ));
    CEMux I__4950 (
            .O(N__25687),
            .I(N__25682));
    CEMux I__4949 (
            .O(N__25686),
            .I(N__25678));
    CEMux I__4948 (
            .O(N__25685),
            .I(N__25675));
    LocalMux I__4947 (
            .O(N__25682),
            .I(N__25672));
    CEMux I__4946 (
            .O(N__25681),
            .I(N__25669));
    LocalMux I__4945 (
            .O(N__25678),
            .I(N__25665));
    LocalMux I__4944 (
            .O(N__25675),
            .I(N__25662));
    Span4Mux_v I__4943 (
            .O(N__25672),
            .I(N__25657));
    LocalMux I__4942 (
            .O(N__25669),
            .I(N__25657));
    CEMux I__4941 (
            .O(N__25668),
            .I(N__25654));
    Span4Mux_v I__4940 (
            .O(N__25665),
            .I(N__25651));
    Span4Mux_v I__4939 (
            .O(N__25662),
            .I(N__25644));
    Span4Mux_v I__4938 (
            .O(N__25657),
            .I(N__25644));
    LocalMux I__4937 (
            .O(N__25654),
            .I(N__25644));
    Span4Mux_h I__4936 (
            .O(N__25651),
            .I(N__25641));
    Span4Mux_h I__4935 (
            .O(N__25644),
            .I(N__25638));
    Odrv4 I__4934 (
            .O(N__25641),
            .I(N_1709_0));
    Odrv4 I__4933 (
            .O(N__25638),
            .I(N_1709_0));
    CEMux I__4932 (
            .O(N__25633),
            .I(N__25628));
    CEMux I__4931 (
            .O(N__25632),
            .I(N__25625));
    CEMux I__4930 (
            .O(N__25631),
            .I(N__25622));
    LocalMux I__4929 (
            .O(N__25628),
            .I(N__25619));
    LocalMux I__4928 (
            .O(N__25625),
            .I(N__25616));
    LocalMux I__4927 (
            .O(N__25622),
            .I(N__25613));
    Span4Mux_h I__4926 (
            .O(N__25619),
            .I(N__25610));
    Span4Mux_h I__4925 (
            .O(N__25616),
            .I(N__25605));
    Span4Mux_h I__4924 (
            .O(N__25613),
            .I(N__25605));
    Odrv4 I__4923 (
            .O(N__25610),
            .I(N_1693_0));
    Odrv4 I__4922 (
            .O(N__25605),
            .I(N_1693_0));
    IoInMux I__4921 (
            .O(N__25600),
            .I(N__25597));
    LocalMux I__4920 (
            .O(N__25597),
            .I(N__25594));
    Span12Mux_s5_v I__4919 (
            .O(N__25594),
            .I(N__25591));
    Odrv12 I__4918 (
            .O(N__25591),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI01JU6Z0Z_9 ));
    CascadeMux I__4917 (
            .O(N__25588),
            .I(\this_ppu.N_1269_cascade_ ));
    InMux I__4916 (
            .O(N__25585),
            .I(N__25582));
    LocalMux I__4915 (
            .O(N__25582),
            .I(N__25579));
    Span4Mux_v I__4914 (
            .O(N__25579),
            .I(N__25576));
    Odrv4 I__4913 (
            .O(N__25576),
            .I(\this_ppu.N_1006_0 ));
    CascadeMux I__4912 (
            .O(N__25573),
            .I(\this_vga_signals.N_1264_cascade_ ));
    InMux I__4911 (
            .O(N__25570),
            .I(N__25567));
    LocalMux I__4910 (
            .O(N__25567),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x0 ));
    CascadeMux I__4909 (
            .O(N__25564),
            .I(\this_ppu.N_1301_cascade_ ));
    InMux I__4908 (
            .O(N__25561),
            .I(N__25558));
    LocalMux I__4907 (
            .O(N__25558),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_CO ));
    CascadeMux I__4906 (
            .O(N__25555),
            .I(N__25552));
    InMux I__4905 (
            .O(N__25552),
            .I(N__25547));
    CascadeMux I__4904 (
            .O(N__25551),
            .I(N__25544));
    CascadeMux I__4903 (
            .O(N__25550),
            .I(N__25541));
    LocalMux I__4902 (
            .O(N__25547),
            .I(N__25538));
    InMux I__4901 (
            .O(N__25544),
            .I(N__25533));
    InMux I__4900 (
            .O(N__25541),
            .I(N__25533));
    Odrv4 I__4899 (
            .O(N__25538),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_6 ));
    LocalMux I__4898 (
            .O(N__25533),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_6 ));
    InMux I__4897 (
            .O(N__25528),
            .I(N__25520));
    InMux I__4896 (
            .O(N__25527),
            .I(N__25509));
    InMux I__4895 (
            .O(N__25526),
            .I(N__25509));
    InMux I__4894 (
            .O(N__25525),
            .I(N__25509));
    InMux I__4893 (
            .O(N__25524),
            .I(N__25509));
    InMux I__4892 (
            .O(N__25523),
            .I(N__25509));
    LocalMux I__4891 (
            .O(N__25520),
            .I(N__25505));
    LocalMux I__4890 (
            .O(N__25509),
            .I(N__25502));
    InMux I__4889 (
            .O(N__25508),
            .I(N__25499));
    Odrv4 I__4888 (
            .O(N__25505),
            .I(\this_ppu.N_1730_0 ));
    Odrv4 I__4887 (
            .O(N__25502),
            .I(\this_ppu.N_1730_0 ));
    LocalMux I__4886 (
            .O(N__25499),
            .I(\this_ppu.N_1730_0 ));
    InMux I__4885 (
            .O(N__25492),
            .I(N__25489));
    LocalMux I__4884 (
            .O(N__25489),
            .I(N__25486));
    Odrv4 I__4883 (
            .O(N__25486),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_CO ));
    InMux I__4882 (
            .O(N__25483),
            .I(N__25475));
    InMux I__4881 (
            .O(N__25482),
            .I(N__25464));
    InMux I__4880 (
            .O(N__25481),
            .I(N__25464));
    InMux I__4879 (
            .O(N__25480),
            .I(N__25464));
    InMux I__4878 (
            .O(N__25479),
            .I(N__25464));
    InMux I__4877 (
            .O(N__25478),
            .I(N__25464));
    LocalMux I__4876 (
            .O(N__25475),
            .I(N__25459));
    LocalMux I__4875 (
            .O(N__25464),
            .I(N__25456));
    InMux I__4874 (
            .O(N__25463),
            .I(N__25453));
    InMux I__4873 (
            .O(N__25462),
            .I(N__25450));
    Odrv12 I__4872 (
            .O(N__25459),
            .I(\this_ppu.N_677_0 ));
    Odrv4 I__4871 (
            .O(N__25456),
            .I(\this_ppu.N_677_0 ));
    LocalMux I__4870 (
            .O(N__25453),
            .I(\this_ppu.N_677_0 ));
    LocalMux I__4869 (
            .O(N__25450),
            .I(\this_ppu.N_677_0 ));
    CascadeMux I__4868 (
            .O(N__25441),
            .I(N__25436));
    CascadeMux I__4867 (
            .O(N__25440),
            .I(N__25433));
    CascadeMux I__4866 (
            .O(N__25439),
            .I(N__25430));
    InMux I__4865 (
            .O(N__25436),
            .I(N__25427));
    InMux I__4864 (
            .O(N__25433),
            .I(N__25424));
    InMux I__4863 (
            .O(N__25430),
            .I(N__25421));
    LocalMux I__4862 (
            .O(N__25427),
            .I(N__25418));
    LocalMux I__4861 (
            .O(N__25424),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_4 ));
    LocalMux I__4860 (
            .O(N__25421),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_4 ));
    Odrv12 I__4859 (
            .O(N__25418),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_4 ));
    InMux I__4858 (
            .O(N__25411),
            .I(N__25408));
    LocalMux I__4857 (
            .O(N__25408),
            .I(N__25405));
    Span4Mux_v I__4856 (
            .O(N__25405),
            .I(N__25402));
    Odrv4 I__4855 (
            .O(N__25402),
            .I(M_this_data_count_q_cry_6_THRU_CO));
    InMux I__4854 (
            .O(N__25399),
            .I(N__25396));
    LocalMux I__4853 (
            .O(N__25396),
            .I(N__25393));
    Odrv4 I__4852 (
            .O(N__25393),
            .I(M_this_data_count_q_cry_8_THRU_CO));
    InMux I__4851 (
            .O(N__25390),
            .I(N__25385));
    CascadeMux I__4850 (
            .O(N__25389),
            .I(N__25382));
    InMux I__4849 (
            .O(N__25388),
            .I(N__25379));
    LocalMux I__4848 (
            .O(N__25385),
            .I(N__25376));
    InMux I__4847 (
            .O(N__25382),
            .I(N__25373));
    LocalMux I__4846 (
            .O(N__25379),
            .I(M_this_data_count_qZ0Z_9));
    Odrv4 I__4845 (
            .O(N__25376),
            .I(M_this_data_count_qZ0Z_9));
    LocalMux I__4844 (
            .O(N__25373),
            .I(M_this_data_count_qZ0Z_9));
    CEMux I__4843 (
            .O(N__25366),
            .I(N__25362));
    CEMux I__4842 (
            .O(N__25365),
            .I(N__25359));
    LocalMux I__4841 (
            .O(N__25362),
            .I(N__25353));
    LocalMux I__4840 (
            .O(N__25359),
            .I(N__25353));
    CEMux I__4839 (
            .O(N__25358),
            .I(N__25350));
    Span4Mux_v I__4838 (
            .O(N__25353),
            .I(N__25347));
    LocalMux I__4837 (
            .O(N__25350),
            .I(N__25344));
    Odrv4 I__4836 (
            .O(N__25347),
            .I(N_231));
    Odrv4 I__4835 (
            .O(N__25344),
            .I(N_231));
    InMux I__4834 (
            .O(N__25339),
            .I(N__25336));
    LocalMux I__4833 (
            .O(N__25336),
            .I(N__25333));
    Span4Mux_h I__4832 (
            .O(N__25333),
            .I(N__25330));
    Odrv4 I__4831 (
            .O(N__25330),
            .I(M_this_data_tmp_qZ0Z_2));
    InMux I__4830 (
            .O(N__25327),
            .I(N__25324));
    LocalMux I__4829 (
            .O(N__25324),
            .I(N__25321));
    Span4Mux_h I__4828 (
            .O(N__25321),
            .I(N__25318));
    Span4Mux_h I__4827 (
            .O(N__25318),
            .I(N__25315));
    Odrv4 I__4826 (
            .O(N__25315),
            .I(M_this_oam_ram_write_data_2));
    InMux I__4825 (
            .O(N__25312),
            .I(N__25307));
    InMux I__4824 (
            .O(N__25311),
            .I(N__25304));
    InMux I__4823 (
            .O(N__25310),
            .I(N__25301));
    LocalMux I__4822 (
            .O(N__25307),
            .I(N__25298));
    LocalMux I__4821 (
            .O(N__25304),
            .I(N__25295));
    LocalMux I__4820 (
            .O(N__25301),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_3 ));
    Odrv12 I__4819 (
            .O(N__25298),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_3 ));
    Odrv4 I__4818 (
            .O(N__25295),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_3 ));
    CascadeMux I__4817 (
            .O(N__25288),
            .I(N__25285));
    InMux I__4816 (
            .O(N__25285),
            .I(N__25282));
    LocalMux I__4815 (
            .O(N__25282),
            .I(N__25279));
    Span4Mux_v I__4814 (
            .O(N__25279),
            .I(N__25276));
    Odrv4 I__4813 (
            .O(N__25276),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_CO ));
    InMux I__4812 (
            .O(N__25273),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1 ));
    InMux I__4811 (
            .O(N__25270),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1 ));
    InMux I__4810 (
            .O(N__25267),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1 ));
    SRMux I__4809 (
            .O(N__25264),
            .I(N__25256));
    SRMux I__4808 (
            .O(N__25263),
            .I(N__25252));
    SRMux I__4807 (
            .O(N__25262),
            .I(N__25248));
    SRMux I__4806 (
            .O(N__25261),
            .I(N__25244));
    IoInMux I__4805 (
            .O(N__25260),
            .I(N__25240));
    SRMux I__4804 (
            .O(N__25259),
            .I(N__25237));
    LocalMux I__4803 (
            .O(N__25256),
            .I(N__25232));
    SRMux I__4802 (
            .O(N__25255),
            .I(N__25229));
    LocalMux I__4801 (
            .O(N__25252),
            .I(N__25224));
    SRMux I__4800 (
            .O(N__25251),
            .I(N__25221));
    LocalMux I__4799 (
            .O(N__25248),
            .I(N__25216));
    SRMux I__4798 (
            .O(N__25247),
            .I(N__25213));
    LocalMux I__4797 (
            .O(N__25244),
            .I(N__25210));
    SRMux I__4796 (
            .O(N__25243),
            .I(N__25207));
    LocalMux I__4795 (
            .O(N__25240),
            .I(N__25200));
    LocalMux I__4794 (
            .O(N__25237),
            .I(N__25196));
    SRMux I__4793 (
            .O(N__25236),
            .I(N__25193));
    SRMux I__4792 (
            .O(N__25235),
            .I(N__25190));
    Span4Mux_s3_v I__4791 (
            .O(N__25232),
            .I(N__25187));
    LocalMux I__4790 (
            .O(N__25229),
            .I(N__25184));
    SRMux I__4789 (
            .O(N__25228),
            .I(N__25181));
    SRMux I__4788 (
            .O(N__25227),
            .I(N__25178));
    Span4Mux_v I__4787 (
            .O(N__25224),
            .I(N__25171));
    LocalMux I__4786 (
            .O(N__25221),
            .I(N__25171));
    SRMux I__4785 (
            .O(N__25220),
            .I(N__25168));
    SRMux I__4784 (
            .O(N__25219),
            .I(N__25165));
    Span4Mux_v I__4783 (
            .O(N__25216),
            .I(N__25155));
    LocalMux I__4782 (
            .O(N__25213),
            .I(N__25155));
    Span4Mux_h I__4781 (
            .O(N__25210),
            .I(N__25155));
    LocalMux I__4780 (
            .O(N__25207),
            .I(N__25155));
    SRMux I__4779 (
            .O(N__25206),
            .I(N__25152));
    SRMux I__4778 (
            .O(N__25205),
            .I(N__25149));
    SRMux I__4777 (
            .O(N__25204),
            .I(N__25146));
    SRMux I__4776 (
            .O(N__25203),
            .I(N__25143));
    IoSpan4Mux I__4775 (
            .O(N__25200),
            .I(N__25139));
    SRMux I__4774 (
            .O(N__25199),
            .I(N__25135));
    Span4Mux_s3_v I__4773 (
            .O(N__25196),
            .I(N__25126));
    LocalMux I__4772 (
            .O(N__25193),
            .I(N__25126));
    LocalMux I__4771 (
            .O(N__25190),
            .I(N__25126));
    Span4Mux_h I__4770 (
            .O(N__25187),
            .I(N__25117));
    Span4Mux_s3_v I__4769 (
            .O(N__25184),
            .I(N__25117));
    LocalMux I__4768 (
            .O(N__25181),
            .I(N__25117));
    LocalMux I__4767 (
            .O(N__25178),
            .I(N__25117));
    SRMux I__4766 (
            .O(N__25177),
            .I(N__25114));
    SRMux I__4765 (
            .O(N__25176),
            .I(N__25111));
    Span4Mux_v I__4764 (
            .O(N__25171),
            .I(N__25103));
    LocalMux I__4763 (
            .O(N__25168),
            .I(N__25103));
    LocalMux I__4762 (
            .O(N__25165),
            .I(N__25103));
    SRMux I__4761 (
            .O(N__25164),
            .I(N__25100));
    Span4Mux_v I__4760 (
            .O(N__25155),
            .I(N__25093));
    LocalMux I__4759 (
            .O(N__25152),
            .I(N__25093));
    LocalMux I__4758 (
            .O(N__25149),
            .I(N__25093));
    LocalMux I__4757 (
            .O(N__25146),
            .I(N__25088));
    LocalMux I__4756 (
            .O(N__25143),
            .I(N__25088));
    SRMux I__4755 (
            .O(N__25142),
            .I(N__25085));
    Span4Mux_s0_h I__4754 (
            .O(N__25139),
            .I(N__25080));
    SRMux I__4753 (
            .O(N__25138),
            .I(N__25077));
    LocalMux I__4752 (
            .O(N__25135),
            .I(N__25068));
    SRMux I__4751 (
            .O(N__25134),
            .I(N__25065));
    SRMux I__4750 (
            .O(N__25133),
            .I(N__25062));
    Span4Mux_v I__4749 (
            .O(N__25126),
            .I(N__25050));
    Span4Mux_v I__4748 (
            .O(N__25117),
            .I(N__25050));
    LocalMux I__4747 (
            .O(N__25114),
            .I(N__25050));
    LocalMux I__4746 (
            .O(N__25111),
            .I(N__25050));
    SRMux I__4745 (
            .O(N__25110),
            .I(N__25047));
    Span4Mux_v I__4744 (
            .O(N__25103),
            .I(N__25036));
    LocalMux I__4743 (
            .O(N__25100),
            .I(N__25036));
    Span4Mux_v I__4742 (
            .O(N__25093),
            .I(N__25036));
    Span4Mux_v I__4741 (
            .O(N__25088),
            .I(N__25036));
    LocalMux I__4740 (
            .O(N__25085),
            .I(N__25036));
    SRMux I__4739 (
            .O(N__25084),
            .I(N__25033));
    SRMux I__4738 (
            .O(N__25083),
            .I(N__25030));
    Span4Mux_h I__4737 (
            .O(N__25080),
            .I(N__25025));
    LocalMux I__4736 (
            .O(N__25077),
            .I(N__25025));
    SRMux I__4735 (
            .O(N__25076),
            .I(N__25022));
    CascadeMux I__4734 (
            .O(N__25075),
            .I(N__25014));
    CascadeMux I__4733 (
            .O(N__25074),
            .I(N__25010));
    CascadeMux I__4732 (
            .O(N__25073),
            .I(N__25006));
    SRMux I__4731 (
            .O(N__25072),
            .I(N__25003));
    SRMux I__4730 (
            .O(N__25071),
            .I(N__25000));
    Span4Mux_s3_v I__4729 (
            .O(N__25068),
            .I(N__24992));
    LocalMux I__4728 (
            .O(N__25065),
            .I(N__24992));
    LocalMux I__4727 (
            .O(N__25062),
            .I(N__24992));
    SRMux I__4726 (
            .O(N__25061),
            .I(N__24988));
    SRMux I__4725 (
            .O(N__25060),
            .I(N__24983));
    SRMux I__4724 (
            .O(N__25059),
            .I(N__24980));
    Span4Mux_v I__4723 (
            .O(N__25050),
            .I(N__24971));
    LocalMux I__4722 (
            .O(N__25047),
            .I(N__24971));
    Span4Mux_v I__4721 (
            .O(N__25036),
            .I(N__24971));
    LocalMux I__4720 (
            .O(N__25033),
            .I(N__24971));
    LocalMux I__4719 (
            .O(N__25030),
            .I(N__24968));
    Span4Mux_h I__4718 (
            .O(N__25025),
            .I(N__24965));
    LocalMux I__4717 (
            .O(N__25022),
            .I(N__24962));
    CascadeMux I__4716 (
            .O(N__25021),
            .I(N__24959));
    CascadeMux I__4715 (
            .O(N__25020),
            .I(N__24955));
    CascadeMux I__4714 (
            .O(N__25019),
            .I(N__24951));
    CascadeMux I__4713 (
            .O(N__25018),
            .I(N__24947));
    InMux I__4712 (
            .O(N__25017),
            .I(N__24934));
    InMux I__4711 (
            .O(N__25014),
            .I(N__24934));
    InMux I__4710 (
            .O(N__25013),
            .I(N__24934));
    InMux I__4709 (
            .O(N__25010),
            .I(N__24934));
    InMux I__4708 (
            .O(N__25009),
            .I(N__24934));
    InMux I__4707 (
            .O(N__25006),
            .I(N__24934));
    LocalMux I__4706 (
            .O(N__25003),
            .I(N__24930));
    LocalMux I__4705 (
            .O(N__25000),
            .I(N__24927));
    SRMux I__4704 (
            .O(N__24999),
            .I(N__24924));
    Span4Mux_v I__4703 (
            .O(N__24992),
            .I(N__24920));
    SRMux I__4702 (
            .O(N__24991),
            .I(N__24917));
    LocalMux I__4701 (
            .O(N__24988),
            .I(N__24914));
    SRMux I__4700 (
            .O(N__24987),
            .I(N__24911));
    SRMux I__4699 (
            .O(N__24986),
            .I(N__24908));
    LocalMux I__4698 (
            .O(N__24983),
            .I(N__24899));
    LocalMux I__4697 (
            .O(N__24980),
            .I(N__24899));
    Span4Mux_v I__4696 (
            .O(N__24971),
            .I(N__24899));
    Span4Mux_h I__4695 (
            .O(N__24968),
            .I(N__24896));
    Span4Mux_v I__4694 (
            .O(N__24965),
            .I(N__24891));
    Span4Mux_h I__4693 (
            .O(N__24962),
            .I(N__24891));
    InMux I__4692 (
            .O(N__24959),
            .I(N__24871));
    InMux I__4691 (
            .O(N__24958),
            .I(N__24871));
    InMux I__4690 (
            .O(N__24955),
            .I(N__24871));
    InMux I__4689 (
            .O(N__24954),
            .I(N__24871));
    InMux I__4688 (
            .O(N__24951),
            .I(N__24871));
    InMux I__4687 (
            .O(N__24950),
            .I(N__24871));
    InMux I__4686 (
            .O(N__24947),
            .I(N__24871));
    LocalMux I__4685 (
            .O(N__24934),
            .I(N__24866));
    InMux I__4684 (
            .O(N__24933),
            .I(N__24863));
    Span4Mux_v I__4683 (
            .O(N__24930),
            .I(N__24856));
    Span4Mux_v I__4682 (
            .O(N__24927),
            .I(N__24856));
    LocalMux I__4681 (
            .O(N__24924),
            .I(N__24856));
    SRMux I__4680 (
            .O(N__24923),
            .I(N__24853));
    Span4Mux_h I__4679 (
            .O(N__24920),
            .I(N__24847));
    LocalMux I__4678 (
            .O(N__24917),
            .I(N__24847));
    Span4Mux_v I__4677 (
            .O(N__24914),
            .I(N__24840));
    LocalMux I__4676 (
            .O(N__24911),
            .I(N__24840));
    LocalMux I__4675 (
            .O(N__24908),
            .I(N__24840));
    SRMux I__4674 (
            .O(N__24907),
            .I(N__24837));
    SRMux I__4673 (
            .O(N__24906),
            .I(N__24834));
    Span4Mux_v I__4672 (
            .O(N__24899),
            .I(N__24830));
    Sp12to4 I__4671 (
            .O(N__24896),
            .I(N__24825));
    Sp12to4 I__4670 (
            .O(N__24891),
            .I(N__24825));
    CascadeMux I__4669 (
            .O(N__24890),
            .I(N__24822));
    CascadeMux I__4668 (
            .O(N__24889),
            .I(N__24819));
    CascadeMux I__4667 (
            .O(N__24888),
            .I(N__24816));
    CascadeMux I__4666 (
            .O(N__24887),
            .I(N__24813));
    CascadeMux I__4665 (
            .O(N__24886),
            .I(N__24810));
    LocalMux I__4664 (
            .O(N__24871),
            .I(N__24807));
    SRMux I__4663 (
            .O(N__24870),
            .I(N__24804));
    IoInMux I__4662 (
            .O(N__24869),
            .I(N__24801));
    Span4Mux_v I__4661 (
            .O(N__24866),
            .I(N__24796));
    LocalMux I__4660 (
            .O(N__24863),
            .I(N__24796));
    Span4Mux_v I__4659 (
            .O(N__24856),
            .I(N__24791));
    LocalMux I__4658 (
            .O(N__24853),
            .I(N__24791));
    SRMux I__4657 (
            .O(N__24852),
            .I(N__24788));
    Span4Mux_v I__4656 (
            .O(N__24847),
            .I(N__24779));
    Span4Mux_v I__4655 (
            .O(N__24840),
            .I(N__24779));
    LocalMux I__4654 (
            .O(N__24837),
            .I(N__24779));
    LocalMux I__4653 (
            .O(N__24834),
            .I(N__24779));
    SRMux I__4652 (
            .O(N__24833),
            .I(N__24776));
    Sp12to4 I__4651 (
            .O(N__24830),
            .I(N__24771));
    Span12Mux_v I__4650 (
            .O(N__24825),
            .I(N__24771));
    InMux I__4649 (
            .O(N__24822),
            .I(N__24766));
    InMux I__4648 (
            .O(N__24819),
            .I(N__24766));
    InMux I__4647 (
            .O(N__24816),
            .I(N__24759));
    InMux I__4646 (
            .O(N__24813),
            .I(N__24759));
    InMux I__4645 (
            .O(N__24810),
            .I(N__24759));
    Span4Mux_v I__4644 (
            .O(N__24807),
            .I(N__24756));
    LocalMux I__4643 (
            .O(N__24804),
            .I(N__24753));
    LocalMux I__4642 (
            .O(N__24801),
            .I(N__24750));
    Span4Mux_h I__4641 (
            .O(N__24796),
            .I(N__24743));
    Span4Mux_v I__4640 (
            .O(N__24791),
            .I(N__24743));
    LocalMux I__4639 (
            .O(N__24788),
            .I(N__24743));
    Span4Mux_v I__4638 (
            .O(N__24779),
            .I(N__24738));
    LocalMux I__4637 (
            .O(N__24776),
            .I(N__24738));
    Span12Mux_h I__4636 (
            .O(N__24771),
            .I(N__24729));
    LocalMux I__4635 (
            .O(N__24766),
            .I(N__24729));
    LocalMux I__4634 (
            .O(N__24759),
            .I(N__24729));
    Sp12to4 I__4633 (
            .O(N__24756),
            .I(N__24729));
    Span4Mux_v I__4632 (
            .O(N__24753),
            .I(N__24726));
    IoSpan4Mux I__4631 (
            .O(N__24750),
            .I(N__24723));
    Span4Mux_h I__4630 (
            .O(N__24743),
            .I(N__24720));
    Span4Mux_v I__4629 (
            .O(N__24738),
            .I(N__24717));
    Span12Mux_h I__4628 (
            .O(N__24729),
            .I(N__24714));
    Span4Mux_h I__4627 (
            .O(N__24726),
            .I(N__24707));
    Span4Mux_s3_h I__4626 (
            .O(N__24723),
            .I(N__24707));
    Span4Mux_h I__4625 (
            .O(N__24720),
            .I(N__24707));
    Span4Mux_h I__4624 (
            .O(N__24717),
            .I(N__24704));
    Odrv12 I__4623 (
            .O(N__24714),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4622 (
            .O(N__24707),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4621 (
            .O(N__24704),
            .I(CONSTANT_ONE_NET));
    InMux I__4620 (
            .O(N__24697),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1 ));
    InMux I__4619 (
            .O(N__24694),
            .I(N__24690));
    InMux I__4618 (
            .O(N__24693),
            .I(N__24687));
    LocalMux I__4617 (
            .O(N__24690),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_7 ));
    LocalMux I__4616 (
            .O(N__24687),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_7 ));
    CascadeMux I__4615 (
            .O(N__24682),
            .I(N__24671));
    InMux I__4614 (
            .O(N__24681),
            .I(N__24661));
    CascadeMux I__4613 (
            .O(N__24680),
            .I(N__24658));
    CascadeMux I__4612 (
            .O(N__24679),
            .I(N__24655));
    InMux I__4611 (
            .O(N__24678),
            .I(N__24652));
    InMux I__4610 (
            .O(N__24677),
            .I(N__24649));
    InMux I__4609 (
            .O(N__24676),
            .I(N__24644));
    InMux I__4608 (
            .O(N__24675),
            .I(N__24644));
    InMux I__4607 (
            .O(N__24674),
            .I(N__24631));
    InMux I__4606 (
            .O(N__24671),
            .I(N__24631));
    InMux I__4605 (
            .O(N__24670),
            .I(N__24631));
    InMux I__4604 (
            .O(N__24669),
            .I(N__24631));
    InMux I__4603 (
            .O(N__24668),
            .I(N__24631));
    InMux I__4602 (
            .O(N__24667),
            .I(N__24631));
    InMux I__4601 (
            .O(N__24666),
            .I(N__24628));
    InMux I__4600 (
            .O(N__24665),
            .I(N__24625));
    InMux I__4599 (
            .O(N__24664),
            .I(N__24622));
    LocalMux I__4598 (
            .O(N__24661),
            .I(N__24619));
    InMux I__4597 (
            .O(N__24658),
            .I(N__24616));
    InMux I__4596 (
            .O(N__24655),
            .I(N__24611));
    LocalMux I__4595 (
            .O(N__24652),
            .I(N__24608));
    LocalMux I__4594 (
            .O(N__24649),
            .I(N__24605));
    LocalMux I__4593 (
            .O(N__24644),
            .I(N__24600));
    LocalMux I__4592 (
            .O(N__24631),
            .I(N__24600));
    LocalMux I__4591 (
            .O(N__24628),
            .I(N__24597));
    LocalMux I__4590 (
            .O(N__24625),
            .I(N__24588));
    LocalMux I__4589 (
            .O(N__24622),
            .I(N__24588));
    Span4Mux_v I__4588 (
            .O(N__24619),
            .I(N__24588));
    LocalMux I__4587 (
            .O(N__24616),
            .I(N__24588));
    InMux I__4586 (
            .O(N__24615),
            .I(N__24583));
    InMux I__4585 (
            .O(N__24614),
            .I(N__24583));
    LocalMux I__4584 (
            .O(N__24611),
            .I(N__24577));
    Span4Mux_v I__4583 (
            .O(N__24608),
            .I(N__24570));
    Span4Mux_h I__4582 (
            .O(N__24605),
            .I(N__24570));
    Span4Mux_h I__4581 (
            .O(N__24600),
            .I(N__24570));
    Span4Mux_v I__4580 (
            .O(N__24597),
            .I(N__24562));
    Span4Mux_v I__4579 (
            .O(N__24588),
            .I(N__24562));
    LocalMux I__4578 (
            .O(N__24583),
            .I(N__24562));
    InMux I__4577 (
            .O(N__24582),
            .I(N__24557));
    InMux I__4576 (
            .O(N__24581),
            .I(N__24557));
    InMux I__4575 (
            .O(N__24580),
            .I(N__24554));
    Span4Mux_h I__4574 (
            .O(N__24577),
            .I(N__24551));
    Span4Mux_h I__4573 (
            .O(N__24570),
            .I(N__24548));
    InMux I__4572 (
            .O(N__24569),
            .I(N__24545));
    Span4Mux_h I__4571 (
            .O(N__24562),
            .I(N__24542));
    LocalMux I__4570 (
            .O(N__24557),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0 ));
    LocalMux I__4569 (
            .O(N__24554),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0 ));
    Odrv4 I__4568 (
            .O(N__24551),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0 ));
    Odrv4 I__4567 (
            .O(N__24548),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0 ));
    LocalMux I__4566 (
            .O(N__24545),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0 ));
    Odrv4 I__4565 (
            .O(N__24542),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0 ));
    InMux I__4564 (
            .O(N__24529),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_6_s1 ));
    InMux I__4563 (
            .O(N__24526),
            .I(N__24523));
    LocalMux I__4562 (
            .O(N__24523),
            .I(\this_ppu.N_1205 ));
    InMux I__4561 (
            .O(N__24520),
            .I(N__24517));
    LocalMux I__4560 (
            .O(N__24517),
            .I(N__24514));
    Odrv4 I__4559 (
            .O(N__24514),
            .I(\this_ppu.M_state_d30_i_i_o2_4 ));
    InMux I__4558 (
            .O(N__24511),
            .I(N__24508));
    LocalMux I__4557 (
            .O(N__24508),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_CO ));
    CascadeMux I__4556 (
            .O(N__24505),
            .I(N__24501));
    InMux I__4555 (
            .O(N__24504),
            .I(N__24497));
    InMux I__4554 (
            .O(N__24501),
            .I(N__24492));
    InMux I__4553 (
            .O(N__24500),
            .I(N__24492));
    LocalMux I__4552 (
            .O(N__24497),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_1 ));
    LocalMux I__4551 (
            .O(N__24492),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_1 ));
    CascadeMux I__4550 (
            .O(N__24487),
            .I(N__24484));
    InMux I__4549 (
            .O(N__24484),
            .I(N__24481));
    LocalMux I__4548 (
            .O(N__24481),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_CO ));
    CascadeMux I__4547 (
            .O(N__24478),
            .I(N__24475));
    InMux I__4546 (
            .O(N__24475),
            .I(N__24470));
    InMux I__4545 (
            .O(N__24474),
            .I(N__24465));
    InMux I__4544 (
            .O(N__24473),
            .I(N__24465));
    LocalMux I__4543 (
            .O(N__24470),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_2 ));
    LocalMux I__4542 (
            .O(N__24465),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_2 ));
    CascadeMux I__4541 (
            .O(N__24460),
            .I(N__24457));
    InMux I__4540 (
            .O(N__24457),
            .I(N__24454));
    LocalMux I__4539 (
            .O(N__24454),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_CO ));
    InMux I__4538 (
            .O(N__24451),
            .I(N__24446));
    InMux I__4537 (
            .O(N__24450),
            .I(N__24441));
    InMux I__4536 (
            .O(N__24449),
            .I(N__24441));
    LocalMux I__4535 (
            .O(N__24446),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_5 ));
    LocalMux I__4534 (
            .O(N__24441),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_5 ));
    InMux I__4533 (
            .O(N__24436),
            .I(N__24433));
    LocalMux I__4532 (
            .O(N__24433),
            .I(\this_ppu.M_state_d30_i_i_o2_3 ));
    InMux I__4531 (
            .O(N__24430),
            .I(N__24425));
    InMux I__4530 (
            .O(N__24429),
            .I(N__24417));
    InMux I__4529 (
            .O(N__24428),
            .I(N__24417));
    LocalMux I__4528 (
            .O(N__24425),
            .I(N__24414));
    InMux I__4527 (
            .O(N__24424),
            .I(N__24411));
    InMux I__4526 (
            .O(N__24423),
            .I(N__24408));
    InMux I__4525 (
            .O(N__24422),
            .I(N__24405));
    LocalMux I__4524 (
            .O(N__24417),
            .I(N__24402));
    Span4Mux_v I__4523 (
            .O(N__24414),
            .I(N__24398));
    LocalMux I__4522 (
            .O(N__24411),
            .I(N__24393));
    LocalMux I__4521 (
            .O(N__24408),
            .I(N__24393));
    LocalMux I__4520 (
            .O(N__24405),
            .I(N__24388));
    Span4Mux_h I__4519 (
            .O(N__24402),
            .I(N__24388));
    InMux I__4518 (
            .O(N__24401),
            .I(N__24385));
    Span4Mux_v I__4517 (
            .O(N__24398),
            .I(N__24382));
    Span4Mux_v I__4516 (
            .O(N__24393),
            .I(N__24377));
    Span4Mux_h I__4515 (
            .O(N__24388),
            .I(N__24377));
    LocalMux I__4514 (
            .O(N__24385),
            .I(N__24374));
    Odrv4 I__4513 (
            .O(N__24382),
            .I(\this_ppu.N_79_0 ));
    Odrv4 I__4512 (
            .O(N__24377),
            .I(\this_ppu.N_79_0 ));
    Odrv4 I__4511 (
            .O(N__24374),
            .I(\this_ppu.N_79_0 ));
    CascadeMux I__4510 (
            .O(N__24367),
            .I(\this_ppu.N_79_0_cascade_ ));
    InMux I__4509 (
            .O(N__24364),
            .I(N__24361));
    LocalMux I__4508 (
            .O(N__24361),
            .I(N__24358));
    Odrv4 I__4507 (
            .O(N__24358),
            .I(\this_ppu.M_pixel_cnt_q_600_1 ));
    CascadeMux I__4506 (
            .O(N__24355),
            .I(N__24352));
    InMux I__4505 (
            .O(N__24352),
            .I(N__24349));
    LocalMux I__4504 (
            .O(N__24349),
            .I(N__24346));
    Odrv4 I__4503 (
            .O(N__24346),
            .I(\this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_i_0_0 ));
    InMux I__4502 (
            .O(N__24343),
            .I(N__24336));
    InMux I__4501 (
            .O(N__24342),
            .I(N__24336));
    InMux I__4500 (
            .O(N__24341),
            .I(N__24333));
    LocalMux I__4499 (
            .O(N__24336),
            .I(N__24330));
    LocalMux I__4498 (
            .O(N__24333),
            .I(N__24327));
    Span4Mux_v I__4497 (
            .O(N__24330),
            .I(N__24324));
    Odrv4 I__4496 (
            .O(N__24327),
            .I(\this_ppu.N_999_0 ));
    Odrv4 I__4495 (
            .O(N__24324),
            .I(\this_ppu.N_999_0 ));
    InMux I__4494 (
            .O(N__24319),
            .I(N__24315));
    InMux I__4493 (
            .O(N__24318),
            .I(N__24312));
    LocalMux I__4492 (
            .O(N__24315),
            .I(N__24308));
    LocalMux I__4491 (
            .O(N__24312),
            .I(N__24305));
    InMux I__4490 (
            .O(N__24311),
            .I(N__24302));
    Span4Mux_v I__4489 (
            .O(N__24308),
            .I(N__24298));
    Span4Mux_v I__4488 (
            .O(N__24305),
            .I(N__24295));
    LocalMux I__4487 (
            .O(N__24302),
            .I(N__24292));
    InMux I__4486 (
            .O(N__24301),
            .I(N__24289));
    Span4Mux_h I__4485 (
            .O(N__24298),
            .I(N__24286));
    Span4Mux_h I__4484 (
            .O(N__24295),
            .I(N__24283));
    Sp12to4 I__4483 (
            .O(N__24292),
            .I(N__24278));
    LocalMux I__4482 (
            .O(N__24289),
            .I(N__24278));
    Odrv4 I__4481 (
            .O(N__24286),
            .I(\this_ppu.N_838_0 ));
    Odrv4 I__4480 (
            .O(N__24283),
            .I(\this_ppu.N_838_0 ));
    Odrv12 I__4479 (
            .O(N__24278),
            .I(\this_ppu.N_838_0 ));
    CascadeMux I__4478 (
            .O(N__24271),
            .I(N__24267));
    InMux I__4477 (
            .O(N__24270),
            .I(N__24264));
    InMux I__4476 (
            .O(N__24267),
            .I(N__24260));
    LocalMux I__4475 (
            .O(N__24264),
            .I(N__24257));
    CascadeMux I__4474 (
            .O(N__24263),
            .I(N__24254));
    LocalMux I__4473 (
            .O(N__24260),
            .I(N__24251));
    Span4Mux_v I__4472 (
            .O(N__24257),
            .I(N__24247));
    InMux I__4471 (
            .O(N__24254),
            .I(N__24244));
    Span4Mux_h I__4470 (
            .O(N__24251),
            .I(N__24241));
    InMux I__4469 (
            .O(N__24250),
            .I(N__24238));
    Odrv4 I__4468 (
            .O(N__24247),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__4467 (
            .O(N__24244),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    Odrv4 I__4466 (
            .O(N__24241),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__4465 (
            .O(N__24238),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    InMux I__4464 (
            .O(N__24229),
            .I(N__24226));
    LocalMux I__4463 (
            .O(N__24226),
            .I(\this_ppu.N_1042_0 ));
    CascadeMux I__4462 (
            .O(N__24223),
            .I(N__24215));
    InMux I__4461 (
            .O(N__24222),
            .I(N__24212));
    InMux I__4460 (
            .O(N__24221),
            .I(N__24209));
    InMux I__4459 (
            .O(N__24220),
            .I(N__24206));
    InMux I__4458 (
            .O(N__24219),
            .I(N__24201));
    InMux I__4457 (
            .O(N__24218),
            .I(N__24201));
    InMux I__4456 (
            .O(N__24215),
            .I(N__24198));
    LocalMux I__4455 (
            .O(N__24212),
            .I(N__24193));
    LocalMux I__4454 (
            .O(N__24209),
            .I(N__24193));
    LocalMux I__4453 (
            .O(N__24206),
            .I(\this_ppu.M_state_qZ0Z_11 ));
    LocalMux I__4452 (
            .O(N__24201),
            .I(\this_ppu.M_state_qZ0Z_11 ));
    LocalMux I__4451 (
            .O(N__24198),
            .I(\this_ppu.M_state_qZ0Z_11 ));
    Odrv12 I__4450 (
            .O(N__24193),
            .I(\this_ppu.M_state_qZ0Z_11 ));
    CEMux I__4449 (
            .O(N__24184),
            .I(N__24168));
    CascadeMux I__4448 (
            .O(N__24183),
            .I(N__24165));
    InMux I__4447 (
            .O(N__24182),
            .I(N__24160));
    InMux I__4446 (
            .O(N__24181),
            .I(N__24157));
    InMux I__4445 (
            .O(N__24180),
            .I(N__24154));
    InMux I__4444 (
            .O(N__24179),
            .I(N__24149));
    InMux I__4443 (
            .O(N__24178),
            .I(N__24149));
    InMux I__4442 (
            .O(N__24177),
            .I(N__24146));
    CascadeMux I__4441 (
            .O(N__24176),
            .I(N__24143));
    InMux I__4440 (
            .O(N__24175),
            .I(N__24125));
    InMux I__4439 (
            .O(N__24174),
            .I(N__24125));
    InMux I__4438 (
            .O(N__24173),
            .I(N__24125));
    InMux I__4437 (
            .O(N__24172),
            .I(N__24125));
    InMux I__4436 (
            .O(N__24171),
            .I(N__24122));
    LocalMux I__4435 (
            .O(N__24168),
            .I(N__24119));
    InMux I__4434 (
            .O(N__24165),
            .I(N__24116));
    CascadeMux I__4433 (
            .O(N__24164),
            .I(N__24110));
    InMux I__4432 (
            .O(N__24163),
            .I(N__24107));
    LocalMux I__4431 (
            .O(N__24160),
            .I(N__24102));
    LocalMux I__4430 (
            .O(N__24157),
            .I(N__24102));
    LocalMux I__4429 (
            .O(N__24154),
            .I(N__24097));
    LocalMux I__4428 (
            .O(N__24149),
            .I(N__24097));
    LocalMux I__4427 (
            .O(N__24146),
            .I(N__24091));
    InMux I__4426 (
            .O(N__24143),
            .I(N__24088));
    InMux I__4425 (
            .O(N__24142),
            .I(N__24085));
    CEMux I__4424 (
            .O(N__24141),
            .I(N__24082));
    InMux I__4423 (
            .O(N__24140),
            .I(N__24078));
    InMux I__4422 (
            .O(N__24139),
            .I(N__24075));
    InMux I__4421 (
            .O(N__24138),
            .I(N__24070));
    InMux I__4420 (
            .O(N__24137),
            .I(N__24070));
    InMux I__4419 (
            .O(N__24136),
            .I(N__24067));
    InMux I__4418 (
            .O(N__24135),
            .I(N__24064));
    InMux I__4417 (
            .O(N__24134),
            .I(N__24061));
    LocalMux I__4416 (
            .O(N__24125),
            .I(N__24056));
    LocalMux I__4415 (
            .O(N__24122),
            .I(N__24056));
    Span4Mux_h I__4414 (
            .O(N__24119),
            .I(N__24051));
    LocalMux I__4413 (
            .O(N__24116),
            .I(N__24051));
    InMux I__4412 (
            .O(N__24115),
            .I(N__24044));
    InMux I__4411 (
            .O(N__24114),
            .I(N__24044));
    InMux I__4410 (
            .O(N__24113),
            .I(N__24044));
    InMux I__4409 (
            .O(N__24110),
            .I(N__24041));
    LocalMux I__4408 (
            .O(N__24107),
            .I(N__24034));
    Span4Mux_v I__4407 (
            .O(N__24102),
            .I(N__24034));
    Span4Mux_h I__4406 (
            .O(N__24097),
            .I(N__24034));
    InMux I__4405 (
            .O(N__24096),
            .I(N__24031));
    InMux I__4404 (
            .O(N__24095),
            .I(N__24026));
    InMux I__4403 (
            .O(N__24094),
            .I(N__24026));
    Span4Mux_h I__4402 (
            .O(N__24091),
            .I(N__24023));
    LocalMux I__4401 (
            .O(N__24088),
            .I(N__24018));
    LocalMux I__4400 (
            .O(N__24085),
            .I(N__24018));
    LocalMux I__4399 (
            .O(N__24082),
            .I(N__24013));
    InMux I__4398 (
            .O(N__24081),
            .I(N__24004));
    LocalMux I__4397 (
            .O(N__24078),
            .I(N__24001));
    LocalMux I__4396 (
            .O(N__24075),
            .I(N__23994));
    LocalMux I__4395 (
            .O(N__24070),
            .I(N__23994));
    LocalMux I__4394 (
            .O(N__24067),
            .I(N__23994));
    LocalMux I__4393 (
            .O(N__24064),
            .I(N__23986));
    LocalMux I__4392 (
            .O(N__24061),
            .I(N__23986));
    Span4Mux_v I__4391 (
            .O(N__24056),
            .I(N__23986));
    Span4Mux_h I__4390 (
            .O(N__24051),
            .I(N__23977));
    LocalMux I__4389 (
            .O(N__24044),
            .I(N__23977));
    LocalMux I__4388 (
            .O(N__24041),
            .I(N__23977));
    Span4Mux_h I__4387 (
            .O(N__24034),
            .I(N__23977));
    LocalMux I__4386 (
            .O(N__24031),
            .I(N__23968));
    LocalMux I__4385 (
            .O(N__24026),
            .I(N__23968));
    Span4Mux_v I__4384 (
            .O(N__24023),
            .I(N__23968));
    Span4Mux_h I__4383 (
            .O(N__24018),
            .I(N__23968));
    InMux I__4382 (
            .O(N__24017),
            .I(N__23963));
    InMux I__4381 (
            .O(N__24016),
            .I(N__23963));
    Span4Mux_v I__4380 (
            .O(N__24013),
            .I(N__23960));
    InMux I__4379 (
            .O(N__24012),
            .I(N__23957));
    InMux I__4378 (
            .O(N__24011),
            .I(N__23946));
    InMux I__4377 (
            .O(N__24010),
            .I(N__23946));
    InMux I__4376 (
            .O(N__24009),
            .I(N__23946));
    InMux I__4375 (
            .O(N__24008),
            .I(N__23946));
    InMux I__4374 (
            .O(N__24007),
            .I(N__23946));
    LocalMux I__4373 (
            .O(N__24004),
            .I(N__23939));
    Span4Mux_v I__4372 (
            .O(N__24001),
            .I(N__23939));
    Span4Mux_v I__4371 (
            .O(N__23994),
            .I(N__23939));
    InMux I__4370 (
            .O(N__23993),
            .I(N__23936));
    Span4Mux_v I__4369 (
            .O(N__23986),
            .I(N__23933));
    Span4Mux_v I__4368 (
            .O(N__23977),
            .I(N__23930));
    Span4Mux_h I__4367 (
            .O(N__23968),
            .I(N__23927));
    LocalMux I__4366 (
            .O(N__23963),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__4365 (
            .O(N__23960),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    LocalMux I__4364 (
            .O(N__23957),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    LocalMux I__4363 (
            .O(N__23946),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__4362 (
            .O(N__23939),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    LocalMux I__4361 (
            .O(N__23936),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__4360 (
            .O(N__23933),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__4359 (
            .O(N__23930),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__4358 (
            .O(N__23927),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    CascadeMux I__4357 (
            .O(N__23908),
            .I(\this_ppu.N_1042_0_cascade_ ));
    InMux I__4356 (
            .O(N__23905),
            .I(N__23902));
    LocalMux I__4355 (
            .O(N__23902),
            .I(N__23899));
    Span4Mux_h I__4354 (
            .O(N__23899),
            .I(N__23896));
    Sp12to4 I__4353 (
            .O(N__23896),
            .I(N__23893));
    Odrv12 I__4352 (
            .O(N__23893),
            .I(\this_ppu.un30_0_a2_i_0 ));
    InMux I__4351 (
            .O(N__23890),
            .I(N__23887));
    LocalMux I__4350 (
            .O(N__23887),
            .I(N__23882));
    InMux I__4349 (
            .O(N__23886),
            .I(N__23877));
    InMux I__4348 (
            .O(N__23885),
            .I(N__23877));
    Odrv4 I__4347 (
            .O(N__23882),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_0 ));
    LocalMux I__4346 (
            .O(N__23877),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_0 ));
    InMux I__4345 (
            .O(N__23872),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1 ));
    InMux I__4344 (
            .O(N__23869),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1 ));
    InMux I__4343 (
            .O(N__23866),
            .I(N__23863));
    LocalMux I__4342 (
            .O(N__23863),
            .I(N__23860));
    Odrv12 I__4341 (
            .O(N__23860),
            .I(\this_vga_signals.g0_2 ));
    CascadeMux I__4340 (
            .O(N__23857),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_cascade_ ));
    CascadeMux I__4339 (
            .O(N__23854),
            .I(N__23851));
    InMux I__4338 (
            .O(N__23851),
            .I(N__23848));
    LocalMux I__4337 (
            .O(N__23848),
            .I(N__23845));
    Span4Mux_h I__4336 (
            .O(N__23845),
            .I(N__23842));
    Span4Mux_h I__4335 (
            .O(N__23842),
            .I(N__23839));
    Odrv4 I__4334 (
            .O(N__23839),
            .I(M_this_vga_signals_address_7));
    CascadeMux I__4333 (
            .O(N__23836),
            .I(N__23832));
    InMux I__4332 (
            .O(N__23835),
            .I(N__23829));
    InMux I__4331 (
            .O(N__23832),
            .I(N__23826));
    LocalMux I__4330 (
            .O(N__23829),
            .I(N__23823));
    LocalMux I__4329 (
            .O(N__23826),
            .I(N__23819));
    Span4Mux_v I__4328 (
            .O(N__23823),
            .I(N__23815));
    InMux I__4327 (
            .O(N__23822),
            .I(N__23812));
    Span4Mux_h I__4326 (
            .O(N__23819),
            .I(N__23809));
    InMux I__4325 (
            .O(N__23818),
            .I(N__23806));
    Odrv4 I__4324 (
            .O(N__23815),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    LocalMux I__4323 (
            .O(N__23812),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    Odrv4 I__4322 (
            .O(N__23809),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    LocalMux I__4321 (
            .O(N__23806),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    InMux I__4320 (
            .O(N__23797),
            .I(N__23794));
    LocalMux I__4319 (
            .O(N__23794),
            .I(N__23790));
    InMux I__4318 (
            .O(N__23793),
            .I(N__23787));
    Span4Mux_v I__4317 (
            .O(N__23790),
            .I(N__23781));
    LocalMux I__4316 (
            .O(N__23787),
            .I(N__23781));
    InMux I__4315 (
            .O(N__23786),
            .I(N__23778));
    Odrv4 I__4314 (
            .O(N__23781),
            .I(\this_ppu.N_82_0 ));
    LocalMux I__4313 (
            .O(N__23778),
            .I(\this_ppu.N_82_0 ));
    InMux I__4312 (
            .O(N__23773),
            .I(N__23766));
    InMux I__4311 (
            .O(N__23772),
            .I(N__23757));
    InMux I__4310 (
            .O(N__23771),
            .I(N__23757));
    InMux I__4309 (
            .O(N__23770),
            .I(N__23757));
    InMux I__4308 (
            .O(N__23769),
            .I(N__23757));
    LocalMux I__4307 (
            .O(N__23766),
            .I(\this_ppu.N_1659_0 ));
    LocalMux I__4306 (
            .O(N__23757),
            .I(\this_ppu.N_1659_0 ));
    InMux I__4305 (
            .O(N__23752),
            .I(N__23746));
    InMux I__4304 (
            .O(N__23751),
            .I(N__23743));
    InMux I__4303 (
            .O(N__23750),
            .I(N__23740));
    InMux I__4302 (
            .O(N__23749),
            .I(N__23737));
    LocalMux I__4301 (
            .O(N__23746),
            .I(N__23733));
    LocalMux I__4300 (
            .O(N__23743),
            .I(N__23730));
    LocalMux I__4299 (
            .O(N__23740),
            .I(N__23727));
    LocalMux I__4298 (
            .O(N__23737),
            .I(N__23724));
    InMux I__4297 (
            .O(N__23736),
            .I(N__23721));
    Span4Mux_v I__4296 (
            .O(N__23733),
            .I(N__23718));
    Span4Mux_h I__4295 (
            .O(N__23730),
            .I(N__23715));
    Span4Mux_h I__4294 (
            .O(N__23727),
            .I(N__23712));
    Span4Mux_h I__4293 (
            .O(N__23724),
            .I(N__23709));
    LocalMux I__4292 (
            .O(N__23721),
            .I(\this_ppu.M_screen_y_qZ0Z_3 ));
    Odrv4 I__4291 (
            .O(N__23718),
            .I(\this_ppu.M_screen_y_qZ0Z_3 ));
    Odrv4 I__4290 (
            .O(N__23715),
            .I(\this_ppu.M_screen_y_qZ0Z_3 ));
    Odrv4 I__4289 (
            .O(N__23712),
            .I(\this_ppu.M_screen_y_qZ0Z_3 ));
    Odrv4 I__4288 (
            .O(N__23709),
            .I(\this_ppu.M_screen_y_qZ0Z_3 ));
    CascadeMux I__4287 (
            .O(N__23698),
            .I(N__23694));
    CascadeMux I__4286 (
            .O(N__23697),
            .I(N__23691));
    InMux I__4285 (
            .O(N__23694),
            .I(N__23688));
    InMux I__4284 (
            .O(N__23691),
            .I(N__23685));
    LocalMux I__4283 (
            .O(N__23688),
            .I(M_this_scroll_qZ0Z_3));
    LocalMux I__4282 (
            .O(N__23685),
            .I(M_this_scroll_qZ0Z_3));
    InMux I__4281 (
            .O(N__23680),
            .I(N__23677));
    LocalMux I__4280 (
            .O(N__23677),
            .I(N__23674));
    Odrv4 I__4279 (
            .O(N__23674),
            .I(\this_ppu.M_screen_y_q_esr_RNIF77F7Z0Z_3 ));
    CascadeMux I__4278 (
            .O(N__23671),
            .I(N__23668));
    InMux I__4277 (
            .O(N__23668),
            .I(N__23662));
    InMux I__4276 (
            .O(N__23667),
            .I(N__23659));
    CascadeMux I__4275 (
            .O(N__23666),
            .I(N__23654));
    InMux I__4274 (
            .O(N__23665),
            .I(N__23650));
    LocalMux I__4273 (
            .O(N__23662),
            .I(N__23647));
    LocalMux I__4272 (
            .O(N__23659),
            .I(N__23644));
    InMux I__4271 (
            .O(N__23658),
            .I(N__23639));
    InMux I__4270 (
            .O(N__23657),
            .I(N__23639));
    InMux I__4269 (
            .O(N__23654),
            .I(N__23636));
    InMux I__4268 (
            .O(N__23653),
            .I(N__23633));
    LocalMux I__4267 (
            .O(N__23650),
            .I(N__23628));
    Span4Mux_h I__4266 (
            .O(N__23647),
            .I(N__23628));
    Span4Mux_v I__4265 (
            .O(N__23644),
            .I(N__23625));
    LocalMux I__4264 (
            .O(N__23639),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    LocalMux I__4263 (
            .O(N__23636),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    LocalMux I__4262 (
            .O(N__23633),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    Odrv4 I__4261 (
            .O(N__23628),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    Odrv4 I__4260 (
            .O(N__23625),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    InMux I__4259 (
            .O(N__23614),
            .I(N__23606));
    CascadeMux I__4258 (
            .O(N__23613),
            .I(N__23603));
    InMux I__4257 (
            .O(N__23612),
            .I(N__23597));
    InMux I__4256 (
            .O(N__23611),
            .I(N__23597));
    InMux I__4255 (
            .O(N__23610),
            .I(N__23593));
    InMux I__4254 (
            .O(N__23609),
            .I(N__23590));
    LocalMux I__4253 (
            .O(N__23606),
            .I(N__23587));
    InMux I__4252 (
            .O(N__23603),
            .I(N__23584));
    InMux I__4251 (
            .O(N__23602),
            .I(N__23581));
    LocalMux I__4250 (
            .O(N__23597),
            .I(N__23578));
    InMux I__4249 (
            .O(N__23596),
            .I(N__23575));
    LocalMux I__4248 (
            .O(N__23593),
            .I(N__23572));
    LocalMux I__4247 (
            .O(N__23590),
            .I(N__23567));
    Span4Mux_h I__4246 (
            .O(N__23587),
            .I(N__23567));
    LocalMux I__4245 (
            .O(N__23584),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    LocalMux I__4244 (
            .O(N__23581),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv4 I__4243 (
            .O(N__23578),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    LocalMux I__4242 (
            .O(N__23575),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv4 I__4241 (
            .O(N__23572),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv4 I__4240 (
            .O(N__23567),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    InMux I__4239 (
            .O(N__23554),
            .I(N__23548));
    InMux I__4238 (
            .O(N__23553),
            .I(N__23548));
    LocalMux I__4237 (
            .O(N__23548),
            .I(\this_ppu.N_61_0 ));
    CascadeMux I__4236 (
            .O(N__23545),
            .I(N__23542));
    InMux I__4235 (
            .O(N__23542),
            .I(N__23539));
    LocalMux I__4234 (
            .O(N__23539),
            .I(N__23536));
    Span4Mux_v I__4233 (
            .O(N__23536),
            .I(N__23532));
    CascadeMux I__4232 (
            .O(N__23535),
            .I(N__23529));
    Span4Mux_h I__4231 (
            .O(N__23532),
            .I(N__23525));
    InMux I__4230 (
            .O(N__23529),
            .I(N__23520));
    InMux I__4229 (
            .O(N__23528),
            .I(N__23520));
    Odrv4 I__4228 (
            .O(N__23525),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__4227 (
            .O(N__23520),
            .I(M_this_ppu_vram_addr_1));
    CascadeMux I__4226 (
            .O(N__23515),
            .I(\this_ppu.N_61_0_cascade_ ));
    CascadeMux I__4225 (
            .O(N__23512),
            .I(N__23509));
    InMux I__4224 (
            .O(N__23509),
            .I(N__23506));
    LocalMux I__4223 (
            .O(N__23506),
            .I(N__23503));
    Span4Mux_h I__4222 (
            .O(N__23503),
            .I(N__23500));
    Span4Mux_h I__4221 (
            .O(N__23500),
            .I(N__23494));
    InMux I__4220 (
            .O(N__23499),
            .I(N__23487));
    InMux I__4219 (
            .O(N__23498),
            .I(N__23487));
    InMux I__4218 (
            .O(N__23497),
            .I(N__23487));
    Odrv4 I__4217 (
            .O(N__23494),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__4216 (
            .O(N__23487),
            .I(M_this_ppu_vram_addr_0));
    InMux I__4215 (
            .O(N__23482),
            .I(N__23470));
    InMux I__4214 (
            .O(N__23481),
            .I(N__23470));
    InMux I__4213 (
            .O(N__23480),
            .I(N__23470));
    InMux I__4212 (
            .O(N__23479),
            .I(N__23470));
    LocalMux I__4211 (
            .O(N__23470),
            .I(\this_ppu.un1_M_screen_x_q_c2 ));
    CascadeMux I__4210 (
            .O(N__23467),
            .I(N__23462));
    InMux I__4209 (
            .O(N__23466),
            .I(N__23456));
    InMux I__4208 (
            .O(N__23465),
            .I(N__23456));
    InMux I__4207 (
            .O(N__23462),
            .I(N__23450));
    InMux I__4206 (
            .O(N__23461),
            .I(N__23447));
    LocalMux I__4205 (
            .O(N__23456),
            .I(N__23444));
    InMux I__4204 (
            .O(N__23455),
            .I(N__23437));
    InMux I__4203 (
            .O(N__23454),
            .I(N__23437));
    InMux I__4202 (
            .O(N__23453),
            .I(N__23437));
    LocalMux I__4201 (
            .O(N__23450),
            .I(N__23434));
    LocalMux I__4200 (
            .O(N__23447),
            .I(\this_ppu.offset_x ));
    Odrv4 I__4199 (
            .O(N__23444),
            .I(\this_ppu.offset_x ));
    LocalMux I__4198 (
            .O(N__23437),
            .I(\this_ppu.offset_x ));
    Odrv4 I__4197 (
            .O(N__23434),
            .I(\this_ppu.offset_x ));
    InMux I__4196 (
            .O(N__23425),
            .I(N__23422));
    LocalMux I__4195 (
            .O(N__23422),
            .I(N__23419));
    Odrv4 I__4194 (
            .O(N__23419),
            .I(\this_ppu.un1_M_surface_x_q_c1 ));
    CascadeMux I__4193 (
            .O(N__23416),
            .I(N__23413));
    CascadeBuf I__4192 (
            .O(N__23413),
            .I(N__23410));
    CascadeMux I__4191 (
            .O(N__23410),
            .I(N__23407));
    InMux I__4190 (
            .O(N__23407),
            .I(N__23404));
    LocalMux I__4189 (
            .O(N__23404),
            .I(N__23401));
    Sp12to4 I__4188 (
            .O(N__23401),
            .I(N__23394));
    CascadeMux I__4187 (
            .O(N__23400),
            .I(N__23391));
    InMux I__4186 (
            .O(N__23399),
            .I(N__23385));
    InMux I__4185 (
            .O(N__23398),
            .I(N__23385));
    CascadeMux I__4184 (
            .O(N__23397),
            .I(N__23382));
    Span12Mux_s7_v I__4183 (
            .O(N__23394),
            .I(N__23379));
    InMux I__4182 (
            .O(N__23391),
            .I(N__23376));
    InMux I__4181 (
            .O(N__23390),
            .I(N__23373));
    LocalMux I__4180 (
            .O(N__23385),
            .I(N__23370));
    InMux I__4179 (
            .O(N__23382),
            .I(N__23367));
    Span12Mux_h I__4178 (
            .O(N__23379),
            .I(N__23364));
    LocalMux I__4177 (
            .O(N__23376),
            .I(M_this_ppu_map_addr_0));
    LocalMux I__4176 (
            .O(N__23373),
            .I(M_this_ppu_map_addr_0));
    Odrv4 I__4175 (
            .O(N__23370),
            .I(M_this_ppu_map_addr_0));
    LocalMux I__4174 (
            .O(N__23367),
            .I(M_this_ppu_map_addr_0));
    Odrv12 I__4173 (
            .O(N__23364),
            .I(M_this_ppu_map_addr_0));
    CascadeMux I__4172 (
            .O(N__23353),
            .I(N__23350));
    InMux I__4171 (
            .O(N__23350),
            .I(N__23347));
    LocalMux I__4170 (
            .O(N__23347),
            .I(N__23340));
    InMux I__4169 (
            .O(N__23346),
            .I(N__23337));
    InMux I__4168 (
            .O(N__23345),
            .I(N__23330));
    InMux I__4167 (
            .O(N__23344),
            .I(N__23330));
    InMux I__4166 (
            .O(N__23343),
            .I(N__23330));
    Span4Mux_v I__4165 (
            .O(N__23340),
            .I(N__23327));
    LocalMux I__4164 (
            .O(N__23337),
            .I(\this_ppu.M_surface_x_qZ0Z_2 ));
    LocalMux I__4163 (
            .O(N__23330),
            .I(\this_ppu.M_surface_x_qZ0Z_2 ));
    Odrv4 I__4162 (
            .O(N__23327),
            .I(\this_ppu.M_surface_x_qZ0Z_2 ));
    CascadeMux I__4161 (
            .O(N__23320),
            .I(\this_ppu.un1_M_surface_x_q_c1_cascade_ ));
    CascadeMux I__4160 (
            .O(N__23317),
            .I(N__23313));
    CascadeMux I__4159 (
            .O(N__23316),
            .I(N__23307));
    InMux I__4158 (
            .O(N__23313),
            .I(N__23304));
    InMux I__4157 (
            .O(N__23312),
            .I(N__23301));
    InMux I__4156 (
            .O(N__23311),
            .I(N__23296));
    InMux I__4155 (
            .O(N__23310),
            .I(N__23296));
    InMux I__4154 (
            .O(N__23307),
            .I(N__23293));
    LocalMux I__4153 (
            .O(N__23304),
            .I(N__23290));
    LocalMux I__4152 (
            .O(N__23301),
            .I(N__23285));
    LocalMux I__4151 (
            .O(N__23296),
            .I(N__23285));
    LocalMux I__4150 (
            .O(N__23293),
            .I(N__23282));
    Odrv4 I__4149 (
            .O(N__23290),
            .I(\this_ppu.M_surface_x_qZ0Z_1 ));
    Odrv4 I__4148 (
            .O(N__23285),
            .I(\this_ppu.M_surface_x_qZ0Z_1 ));
    Odrv4 I__4147 (
            .O(N__23282),
            .I(\this_ppu.M_surface_x_qZ0Z_1 ));
    InMux I__4146 (
            .O(N__23275),
            .I(N__23272));
    LocalMux I__4145 (
            .O(N__23272),
            .I(N__23268));
    InMux I__4144 (
            .O(N__23271),
            .I(N__23265));
    Span4Mux_v I__4143 (
            .O(N__23268),
            .I(N__23262));
    LocalMux I__4142 (
            .O(N__23265),
            .I(N__23259));
    Odrv4 I__4141 (
            .O(N__23262),
            .I(\this_ppu.un1_M_surface_x_q_c4 ));
    Odrv12 I__4140 (
            .O(N__23259),
            .I(\this_ppu.un1_M_surface_x_q_c4 ));
    InMux I__4139 (
            .O(N__23254),
            .I(N__23251));
    LocalMux I__4138 (
            .O(N__23251),
            .I(N__23246));
    InMux I__4137 (
            .O(N__23250),
            .I(N__23243));
    CascadeMux I__4136 (
            .O(N__23249),
            .I(N__23239));
    Span4Mux_v I__4135 (
            .O(N__23246),
            .I(N__23234));
    LocalMux I__4134 (
            .O(N__23243),
            .I(N__23234));
    InMux I__4133 (
            .O(N__23242),
            .I(N__23231));
    InMux I__4132 (
            .O(N__23239),
            .I(N__23228));
    Span4Mux_h I__4131 (
            .O(N__23234),
            .I(N__23223));
    LocalMux I__4130 (
            .O(N__23231),
            .I(N__23223));
    LocalMux I__4129 (
            .O(N__23228),
            .I(N__23219));
    Span4Mux_h I__4128 (
            .O(N__23223),
            .I(N__23216));
    InMux I__4127 (
            .O(N__23222),
            .I(N__23213));
    Span4Mux_h I__4126 (
            .O(N__23219),
            .I(N__23210));
    Odrv4 I__4125 (
            .O(N__23216),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    LocalMux I__4124 (
            .O(N__23213),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    Odrv4 I__4123 (
            .O(N__23210),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    InMux I__4122 (
            .O(N__23203),
            .I(N__23197));
    InMux I__4121 (
            .O(N__23202),
            .I(N__23194));
    InMux I__4120 (
            .O(N__23201),
            .I(N__23191));
    InMux I__4119 (
            .O(N__23200),
            .I(N__23188));
    LocalMux I__4118 (
            .O(N__23197),
            .I(\this_ppu.M_state_qZ0Z_10 ));
    LocalMux I__4117 (
            .O(N__23194),
            .I(\this_ppu.M_state_qZ0Z_10 ));
    LocalMux I__4116 (
            .O(N__23191),
            .I(\this_ppu.M_state_qZ0Z_10 ));
    LocalMux I__4115 (
            .O(N__23188),
            .I(\this_ppu.M_state_qZ0Z_10 ));
    CascadeMux I__4114 (
            .O(N__23179),
            .I(N__23176));
    InMux I__4113 (
            .O(N__23176),
            .I(N__23173));
    LocalMux I__4112 (
            .O(N__23173),
            .I(N__23167));
    InMux I__4111 (
            .O(N__23172),
            .I(N__23163));
    CascadeMux I__4110 (
            .O(N__23171),
            .I(N__23160));
    CascadeMux I__4109 (
            .O(N__23170),
            .I(N__23157));
    Span4Mux_h I__4108 (
            .O(N__23167),
            .I(N__23153));
    InMux I__4107 (
            .O(N__23166),
            .I(N__23150));
    LocalMux I__4106 (
            .O(N__23163),
            .I(N__23147));
    InMux I__4105 (
            .O(N__23160),
            .I(N__23140));
    InMux I__4104 (
            .O(N__23157),
            .I(N__23140));
    InMux I__4103 (
            .O(N__23156),
            .I(N__23140));
    Span4Mux_h I__4102 (
            .O(N__23153),
            .I(N__23133));
    LocalMux I__4101 (
            .O(N__23150),
            .I(N__23133));
    Span4Mux_h I__4100 (
            .O(N__23147),
            .I(N__23133));
    LocalMux I__4099 (
            .O(N__23140),
            .I(M_this_ppu_vram_addr_3));
    Odrv4 I__4098 (
            .O(N__23133),
            .I(M_this_ppu_vram_addr_3));
    CascadeMux I__4097 (
            .O(N__23128),
            .I(\this_ppu.N_798_0_cascade_ ));
    InMux I__4096 (
            .O(N__23125),
            .I(N__23122));
    LocalMux I__4095 (
            .O(N__23122),
            .I(N__23119));
    Span12Mux_h I__4094 (
            .O(N__23119),
            .I(N__23116));
    Odrv12 I__4093 (
            .O(N__23116),
            .I(M_this_ppu_vram_data_0));
    InMux I__4092 (
            .O(N__23113),
            .I(N__23108));
    InMux I__4091 (
            .O(N__23112),
            .I(N__23105));
    InMux I__4090 (
            .O(N__23111),
            .I(N__23102));
    LocalMux I__4089 (
            .O(N__23108),
            .I(N__23099));
    LocalMux I__4088 (
            .O(N__23105),
            .I(N__23096));
    LocalMux I__4087 (
            .O(N__23102),
            .I(N__23093));
    Span4Mux_v I__4086 (
            .O(N__23099),
            .I(N__23088));
    Span4Mux_h I__4085 (
            .O(N__23096),
            .I(N__23088));
    Odrv4 I__4084 (
            .O(N__23093),
            .I(\this_ppu.N_1182_1 ));
    Odrv4 I__4083 (
            .O(N__23088),
            .I(\this_ppu.N_1182_1 ));
    CascadeMux I__4082 (
            .O(N__23083),
            .I(N__23078));
    CascadeMux I__4081 (
            .O(N__23082),
            .I(N__23075));
    InMux I__4080 (
            .O(N__23081),
            .I(N__23068));
    InMux I__4079 (
            .O(N__23078),
            .I(N__23068));
    InMux I__4078 (
            .O(N__23075),
            .I(N__23065));
    InMux I__4077 (
            .O(N__23074),
            .I(N__23061));
    InMux I__4076 (
            .O(N__23073),
            .I(N__23058));
    LocalMux I__4075 (
            .O(N__23068),
            .I(N__23055));
    LocalMux I__4074 (
            .O(N__23065),
            .I(N__23052));
    InMux I__4073 (
            .O(N__23064),
            .I(N__23049));
    LocalMux I__4072 (
            .O(N__23061),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    LocalMux I__4071 (
            .O(N__23058),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    Odrv4 I__4070 (
            .O(N__23055),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    Odrv4 I__4069 (
            .O(N__23052),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    LocalMux I__4068 (
            .O(N__23049),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    CascadeMux I__4067 (
            .O(N__23038),
            .I(\this_vga_signals.M_lcounter_q_e_1_0_cascade_ ));
    CEMux I__4066 (
            .O(N__23035),
            .I(N__23032));
    LocalMux I__4065 (
            .O(N__23032),
            .I(N__23029));
    Span4Mux_h I__4064 (
            .O(N__23029),
            .I(N__23026));
    Span4Mux_h I__4063 (
            .O(N__23026),
            .I(N__23023));
    Span4Mux_v I__4062 (
            .O(N__23023),
            .I(N__23020));
    Odrv4 I__4061 (
            .O(N__23020),
            .I(N_26));
    InMux I__4060 (
            .O(N__23017),
            .I(N__23014));
    LocalMux I__4059 (
            .O(N__23014),
            .I(\this_ppu.N_1198 ));
    CascadeMux I__4058 (
            .O(N__23011),
            .I(\this_ppu.N_1198_cascade_ ));
    CascadeMux I__4057 (
            .O(N__23008),
            .I(N__23005));
    CascadeBuf I__4056 (
            .O(N__23005),
            .I(N__23001));
    CascadeMux I__4055 (
            .O(N__23004),
            .I(N__22998));
    CascadeMux I__4054 (
            .O(N__23001),
            .I(N__22994));
    InMux I__4053 (
            .O(N__22998),
            .I(N__22991));
    CascadeMux I__4052 (
            .O(N__22997),
            .I(N__22988));
    InMux I__4051 (
            .O(N__22994),
            .I(N__22983));
    LocalMux I__4050 (
            .O(N__22991),
            .I(N__22980));
    InMux I__4049 (
            .O(N__22988),
            .I(N__22977));
    InMux I__4048 (
            .O(N__22987),
            .I(N__22974));
    InMux I__4047 (
            .O(N__22986),
            .I(N__22971));
    LocalMux I__4046 (
            .O(N__22983),
            .I(N__22968));
    Span4Mux_h I__4045 (
            .O(N__22980),
            .I(N__22964));
    LocalMux I__4044 (
            .O(N__22977),
            .I(N__22961));
    LocalMux I__4043 (
            .O(N__22974),
            .I(N__22956));
    LocalMux I__4042 (
            .O(N__22971),
            .I(N__22956));
    Span12Mux_s2_v I__4041 (
            .O(N__22968),
            .I(N__22953));
    InMux I__4040 (
            .O(N__22967),
            .I(N__22950));
    Span4Mux_v I__4039 (
            .O(N__22964),
            .I(N__22947));
    Span4Mux_h I__4038 (
            .O(N__22961),
            .I(N__22944));
    Span12Mux_h I__4037 (
            .O(N__22956),
            .I(N__22939));
    Span12Mux_h I__4036 (
            .O(N__22953),
            .I(N__22939));
    LocalMux I__4035 (
            .O(N__22950),
            .I(M_this_ppu_map_addr_1));
    Odrv4 I__4034 (
            .O(N__22947),
            .I(M_this_ppu_map_addr_1));
    Odrv4 I__4033 (
            .O(N__22944),
            .I(M_this_ppu_map_addr_1));
    Odrv12 I__4032 (
            .O(N__22939),
            .I(M_this_ppu_map_addr_1));
    CascadeMux I__4031 (
            .O(N__22930),
            .I(\this_ppu.un1_M_surface_x_q_c2_cascade_ ));
    CascadeMux I__4030 (
            .O(N__22927),
            .I(\this_ppu.un1_M_surface_x_q_c5_cascade_ ));
    CascadeMux I__4029 (
            .O(N__22924),
            .I(N__22921));
    CascadeBuf I__4028 (
            .O(N__22921),
            .I(N__22918));
    CascadeMux I__4027 (
            .O(N__22918),
            .I(N__22915));
    InMux I__4026 (
            .O(N__22915),
            .I(N__22911));
    CascadeMux I__4025 (
            .O(N__22914),
            .I(N__22908));
    LocalMux I__4024 (
            .O(N__22911),
            .I(N__22905));
    InMux I__4023 (
            .O(N__22908),
            .I(N__22901));
    Span4Mux_s2_v I__4022 (
            .O(N__22905),
            .I(N__22898));
    InMux I__4021 (
            .O(N__22904),
            .I(N__22895));
    LocalMux I__4020 (
            .O(N__22901),
            .I(N__22892));
    Sp12to4 I__4019 (
            .O(N__22898),
            .I(N__22889));
    LocalMux I__4018 (
            .O(N__22895),
            .I(N__22882));
    Span4Mux_v I__4017 (
            .O(N__22892),
            .I(N__22882));
    Span12Mux_h I__4016 (
            .O(N__22889),
            .I(N__22879));
    InMux I__4015 (
            .O(N__22888),
            .I(N__22876));
    InMux I__4014 (
            .O(N__22887),
            .I(N__22873));
    Span4Mux_h I__4013 (
            .O(N__22882),
            .I(N__22870));
    Span12Mux_v I__4012 (
            .O(N__22879),
            .I(N__22867));
    LocalMux I__4011 (
            .O(N__22876),
            .I(M_this_ppu_map_addr_2));
    LocalMux I__4010 (
            .O(N__22873),
            .I(M_this_ppu_map_addr_2));
    Odrv4 I__4009 (
            .O(N__22870),
            .I(M_this_ppu_map_addr_2));
    Odrv12 I__4008 (
            .O(N__22867),
            .I(M_this_ppu_map_addr_2));
    InMux I__4007 (
            .O(N__22858),
            .I(N__22855));
    LocalMux I__4006 (
            .O(N__22855),
            .I(\this_ppu.un1_M_surface_x_q_c2 ));
    InMux I__4005 (
            .O(N__22852),
            .I(N__22849));
    LocalMux I__4004 (
            .O(N__22849),
            .I(N__22846));
    Odrv4 I__4003 (
            .O(N__22846),
            .I(M_this_data_count_q_s_13));
    CascadeMux I__4002 (
            .O(N__22843),
            .I(N__22839));
    InMux I__4001 (
            .O(N__22842),
            .I(N__22835));
    InMux I__4000 (
            .O(N__22839),
            .I(N__22830));
    InMux I__3999 (
            .O(N__22838),
            .I(N__22830));
    LocalMux I__3998 (
            .O(N__22835),
            .I(M_this_data_count_qZ0Z_12));
    LocalMux I__3997 (
            .O(N__22830),
            .I(M_this_data_count_qZ0Z_12));
    InMux I__3996 (
            .O(N__22825),
            .I(N__22820));
    InMux I__3995 (
            .O(N__22824),
            .I(N__22815));
    InMux I__3994 (
            .O(N__22823),
            .I(N__22815));
    LocalMux I__3993 (
            .O(N__22820),
            .I(M_this_data_count_qZ0Z_11));
    LocalMux I__3992 (
            .O(N__22815),
            .I(M_this_data_count_qZ0Z_11));
    CascadeMux I__3991 (
            .O(N__22810),
            .I(N__22806));
    InMux I__3990 (
            .O(N__22809),
            .I(N__22803));
    InMux I__3989 (
            .O(N__22806),
            .I(N__22800));
    LocalMux I__3988 (
            .O(N__22803),
            .I(M_this_data_count_qZ0Z_13));
    LocalMux I__3987 (
            .O(N__22800),
            .I(M_this_data_count_qZ0Z_13));
    InMux I__3986 (
            .O(N__22795),
            .I(N__22791));
    InMux I__3985 (
            .O(N__22794),
            .I(N__22788));
    LocalMux I__3984 (
            .O(N__22791),
            .I(M_this_data_count_qZ0Z_10));
    LocalMux I__3983 (
            .O(N__22788),
            .I(M_this_data_count_qZ0Z_10));
    InMux I__3982 (
            .O(N__22783),
            .I(N__22780));
    LocalMux I__3981 (
            .O(N__22780),
            .I(M_this_data_count_q_s_8));
    InMux I__3980 (
            .O(N__22777),
            .I(N__22773));
    InMux I__3979 (
            .O(N__22776),
            .I(N__22770));
    LocalMux I__3978 (
            .O(N__22773),
            .I(M_this_data_count_qZ0Z_8));
    LocalMux I__3977 (
            .O(N__22770),
            .I(M_this_data_count_qZ0Z_8));
    InMux I__3976 (
            .O(N__22765),
            .I(N__22760));
    InMux I__3975 (
            .O(N__22764),
            .I(N__22757));
    InMux I__3974 (
            .O(N__22763),
            .I(N__22754));
    LocalMux I__3973 (
            .O(N__22760),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__3972 (
            .O(N__22757),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__3971 (
            .O(N__22754),
            .I(M_this_data_count_qZ0Z_5));
    CascadeMux I__3970 (
            .O(N__22747),
            .I(N__22743));
    InMux I__3969 (
            .O(N__22746),
            .I(N__22739));
    InMux I__3968 (
            .O(N__22743),
            .I(N__22736));
    InMux I__3967 (
            .O(N__22742),
            .I(N__22733));
    LocalMux I__3966 (
            .O(N__22739),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__3965 (
            .O(N__22736),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__3964 (
            .O(N__22733),
            .I(M_this_data_count_qZ0Z_4));
    InMux I__3963 (
            .O(N__22726),
            .I(N__22723));
    LocalMux I__3962 (
            .O(N__22723),
            .I(un1_M_this_oam_address_q_c6));
    InMux I__3961 (
            .O(N__22720),
            .I(N__22717));
    LocalMux I__3960 (
            .O(N__22717),
            .I(N__22714));
    Span12Mux_h I__3959 (
            .O(N__22714),
            .I(N__22711));
    Odrv12 I__3958 (
            .O(N__22711),
            .I(\this_vga_signals.g0_1 ));
    InMux I__3957 (
            .O(N__22708),
            .I(N__22704));
    InMux I__3956 (
            .O(N__22707),
            .I(N__22701));
    LocalMux I__3955 (
            .O(N__22704),
            .I(N__22698));
    LocalMux I__3954 (
            .O(N__22701),
            .I(\this_vga_signals.N_3_0 ));
    Odrv4 I__3953 (
            .O(N__22698),
            .I(\this_vga_signals.N_3_0 ));
    InMux I__3952 (
            .O(N__22693),
            .I(N__22690));
    LocalMux I__3951 (
            .O(N__22690),
            .I(N__22687));
    Span4Mux_h I__3950 (
            .O(N__22687),
            .I(N__22683));
    InMux I__3949 (
            .O(N__22686),
            .I(N__22680));
    Span4Mux_v I__3948 (
            .O(N__22683),
            .I(N__22677));
    LocalMux I__3947 (
            .O(N__22680),
            .I(N__22674));
    Odrv4 I__3946 (
            .O(N__22677),
            .I(\this_vga_signals.M_pcounter_q_i_2_1 ));
    Odrv12 I__3945 (
            .O(N__22674),
            .I(\this_vga_signals.M_pcounter_q_i_2_1 ));
    InMux I__3944 (
            .O(N__22669),
            .I(N__22666));
    LocalMux I__3943 (
            .O(N__22666),
            .I(N__22663));
    Span12Mux_v I__3942 (
            .O(N__22663),
            .I(N__22660));
    Odrv12 I__3941 (
            .O(N__22660),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO ));
    CascadeMux I__3940 (
            .O(N__22657),
            .I(N__22654));
    CascadeBuf I__3939 (
            .O(N__22654),
            .I(N__22650));
    CascadeMux I__3938 (
            .O(N__22653),
            .I(N__22647));
    CascadeMux I__3937 (
            .O(N__22650),
            .I(N__22644));
    InMux I__3936 (
            .O(N__22647),
            .I(N__22640));
    InMux I__3935 (
            .O(N__22644),
            .I(N__22637));
    CascadeMux I__3934 (
            .O(N__22643),
            .I(N__22633));
    LocalMux I__3933 (
            .O(N__22640),
            .I(N__22630));
    LocalMux I__3932 (
            .O(N__22637),
            .I(N__22627));
    CascadeMux I__3931 (
            .O(N__22636),
            .I(N__22624));
    InMux I__3930 (
            .O(N__22633),
            .I(N__22621));
    Span4Mux_h I__3929 (
            .O(N__22630),
            .I(N__22618));
    Span4Mux_h I__3928 (
            .O(N__22627),
            .I(N__22615));
    InMux I__3927 (
            .O(N__22624),
            .I(N__22612));
    LocalMux I__3926 (
            .O(N__22621),
            .I(N__22609));
    Span4Mux_h I__3925 (
            .O(N__22618),
            .I(N__22606));
    Span4Mux_h I__3924 (
            .O(N__22615),
            .I(N__22603));
    LocalMux I__3923 (
            .O(N__22612),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_2 ));
    Odrv12 I__3922 (
            .O(N__22609),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_2 ));
    Odrv4 I__3921 (
            .O(N__22606),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_2 ));
    Odrv4 I__3920 (
            .O(N__22603),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_2 ));
    InMux I__3919 (
            .O(N__22594),
            .I(N__22591));
    LocalMux I__3918 (
            .O(N__22591),
            .I(M_this_data_count_q_cry_0_THRU_CO));
    InMux I__3917 (
            .O(N__22588),
            .I(N__22583));
    InMux I__3916 (
            .O(N__22587),
            .I(N__22578));
    InMux I__3915 (
            .O(N__22586),
            .I(N__22578));
    LocalMux I__3914 (
            .O(N__22583),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__3913 (
            .O(N__22578),
            .I(M_this_data_count_qZ0Z_1));
    InMux I__3912 (
            .O(N__22573),
            .I(N__22570));
    LocalMux I__3911 (
            .O(N__22570),
            .I(M_this_data_count_q_cry_1_THRU_CO));
    CascadeMux I__3910 (
            .O(N__22567),
            .I(N__22564));
    InMux I__3909 (
            .O(N__22564),
            .I(N__22559));
    InMux I__3908 (
            .O(N__22563),
            .I(N__22554));
    InMux I__3907 (
            .O(N__22562),
            .I(N__22554));
    LocalMux I__3906 (
            .O(N__22559),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__3905 (
            .O(N__22554),
            .I(M_this_data_count_qZ0Z_2));
    InMux I__3904 (
            .O(N__22549),
            .I(N__22546));
    LocalMux I__3903 (
            .O(N__22546),
            .I(M_this_data_count_q_cry_2_THRU_CO));
    CascadeMux I__3902 (
            .O(N__22543),
            .I(N__22538));
    CascadeMux I__3901 (
            .O(N__22542),
            .I(N__22535));
    InMux I__3900 (
            .O(N__22541),
            .I(N__22532));
    InMux I__3899 (
            .O(N__22538),
            .I(N__22527));
    InMux I__3898 (
            .O(N__22535),
            .I(N__22527));
    LocalMux I__3897 (
            .O(N__22532),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__3896 (
            .O(N__22527),
            .I(M_this_data_count_qZ0Z_3));
    InMux I__3895 (
            .O(N__22522),
            .I(N__22519));
    LocalMux I__3894 (
            .O(N__22519),
            .I(M_this_data_count_q_cry_3_THRU_CO));
    InMux I__3893 (
            .O(N__22516),
            .I(N__22513));
    LocalMux I__3892 (
            .O(N__22513),
            .I(M_this_data_count_q_cry_4_THRU_CO));
    InMux I__3891 (
            .O(N__22510),
            .I(N__22507));
    LocalMux I__3890 (
            .O(N__22507),
            .I(M_this_data_count_q_cry_5_THRU_CO));
    InMux I__3889 (
            .O(N__22504),
            .I(N__22501));
    LocalMux I__3888 (
            .O(N__22501),
            .I(M_this_data_count_q_cry_10_THRU_CO));
    InMux I__3887 (
            .O(N__22498),
            .I(N__22495));
    LocalMux I__3886 (
            .O(N__22495),
            .I(N__22492));
    Odrv4 I__3885 (
            .O(N__22492),
            .I(M_this_data_count_q_s_10));
    InMux I__3884 (
            .O(N__22489),
            .I(N__22486));
    LocalMux I__3883 (
            .O(N__22486),
            .I(M_this_data_count_q_cry_11_THRU_CO));
    CascadeMux I__3882 (
            .O(N__22483),
            .I(N__22480));
    InMux I__3881 (
            .O(N__22480),
            .I(N__22477));
    LocalMux I__3880 (
            .O(N__22477),
            .I(M_this_scroll_qZ0Z_2));
    CascadeMux I__3879 (
            .O(N__22474),
            .I(N__22471));
    InMux I__3878 (
            .O(N__22471),
            .I(N__22467));
    CascadeMux I__3877 (
            .O(N__22470),
            .I(N__22464));
    LocalMux I__3876 (
            .O(N__22467),
            .I(N__22461));
    InMux I__3875 (
            .O(N__22464),
            .I(N__22458));
    Span4Mux_h I__3874 (
            .O(N__22461),
            .I(N__22455));
    LocalMux I__3873 (
            .O(N__22458),
            .I(N__22452));
    Odrv4 I__3872 (
            .O(N__22455),
            .I(M_this_scroll_qZ0Z_4));
    Odrv4 I__3871 (
            .O(N__22452),
            .I(M_this_scroll_qZ0Z_4));
    InMux I__3870 (
            .O(N__22447),
            .I(N__22444));
    LocalMux I__3869 (
            .O(N__22444),
            .I(M_this_scroll_qZ0Z_7));
    IoInMux I__3868 (
            .O(N__22441),
            .I(N__22438));
    LocalMux I__3867 (
            .O(N__22438),
            .I(N__22435));
    Span12Mux_s1_v I__3866 (
            .O(N__22435),
            .I(N__22432));
    Span12Mux_h I__3865 (
            .O(N__22432),
            .I(N__22429));
    Odrv12 I__3864 (
            .O(N__22429),
            .I(this_vga_signals_vsync_1_i));
    InMux I__3863 (
            .O(N__22426),
            .I(N__22421));
    InMux I__3862 (
            .O(N__22425),
            .I(N__22416));
    InMux I__3861 (
            .O(N__22424),
            .I(N__22416));
    LocalMux I__3860 (
            .O(N__22421),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__3859 (
            .O(N__22416),
            .I(M_this_data_count_qZ0Z_0));
    CascadeMux I__3858 (
            .O(N__22411),
            .I(N__22408));
    InMux I__3857 (
            .O(N__22408),
            .I(N__22405));
    LocalMux I__3856 (
            .O(N__22405),
            .I(N__22398));
    InMux I__3855 (
            .O(N__22404),
            .I(N__22395));
    InMux I__3854 (
            .O(N__22403),
            .I(N__22391));
    InMux I__3853 (
            .O(N__22402),
            .I(N__22388));
    CascadeMux I__3852 (
            .O(N__22401),
            .I(N__22385));
    Span4Mux_v I__3851 (
            .O(N__22398),
            .I(N__22381));
    LocalMux I__3850 (
            .O(N__22395),
            .I(N__22378));
    InMux I__3849 (
            .O(N__22394),
            .I(N__22375));
    LocalMux I__3848 (
            .O(N__22391),
            .I(N__22370));
    LocalMux I__3847 (
            .O(N__22388),
            .I(N__22370));
    InMux I__3846 (
            .O(N__22385),
            .I(N__22367));
    InMux I__3845 (
            .O(N__22384),
            .I(N__22364));
    Span4Mux_h I__3844 (
            .O(N__22381),
            .I(N__22361));
    Span4Mux_v I__3843 (
            .O(N__22378),
            .I(N__22354));
    LocalMux I__3842 (
            .O(N__22375),
            .I(N__22354));
    Span4Mux_v I__3841 (
            .O(N__22370),
            .I(N__22354));
    LocalMux I__3840 (
            .O(N__22367),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__3839 (
            .O(N__22364),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__3838 (
            .O(N__22361),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__3837 (
            .O(N__22354),
            .I(M_this_ppu_vram_addr_7));
    InMux I__3836 (
            .O(N__22345),
            .I(N__22342));
    LocalMux I__3835 (
            .O(N__22342),
            .I(\this_ppu.M_screen_y_q_RNIQ9FQ6Z0Z_0 ));
    CascadeMux I__3834 (
            .O(N__22339),
            .I(\this_ppu.un1_M_screen_x_q_c4_cascade_ ));
    InMux I__3833 (
            .O(N__22336),
            .I(N__22333));
    LocalMux I__3832 (
            .O(N__22333),
            .I(\this_ppu.un1_M_screen_x_q_c4 ));
    CascadeMux I__3831 (
            .O(N__22330),
            .I(N__22327));
    InMux I__3830 (
            .O(N__22327),
            .I(N__22324));
    LocalMux I__3829 (
            .O(N__22324),
            .I(N__22321));
    Span4Mux_h I__3828 (
            .O(N__22321),
            .I(N__22317));
    CascadeMux I__3827 (
            .O(N__22320),
            .I(N__22314));
    Span4Mux_h I__3826 (
            .O(N__22317),
            .I(N__22309));
    InMux I__3825 (
            .O(N__22314),
            .I(N__22302));
    InMux I__3824 (
            .O(N__22313),
            .I(N__22302));
    InMux I__3823 (
            .O(N__22312),
            .I(N__22302));
    Odrv4 I__3822 (
            .O(N__22309),
            .I(M_this_ppu_vram_addr_4));
    LocalMux I__3821 (
            .O(N__22302),
            .I(M_this_ppu_vram_addr_4));
    CascadeMux I__3820 (
            .O(N__22297),
            .I(\this_ppu.un1_M_screen_x_q_c5_cascade_ ));
    CascadeMux I__3819 (
            .O(N__22294),
            .I(N__22291));
    InMux I__3818 (
            .O(N__22291),
            .I(N__22288));
    LocalMux I__3817 (
            .O(N__22288),
            .I(N__22285));
    Span4Mux_v I__3816 (
            .O(N__22285),
            .I(N__22282));
    Span4Mux_h I__3815 (
            .O(N__22282),
            .I(N__22277));
    InMux I__3814 (
            .O(N__22281),
            .I(N__22272));
    InMux I__3813 (
            .O(N__22280),
            .I(N__22272));
    Odrv4 I__3812 (
            .O(N__22277),
            .I(M_this_ppu_vram_addr_5));
    LocalMux I__3811 (
            .O(N__22272),
            .I(M_this_ppu_vram_addr_5));
    CascadeMux I__3810 (
            .O(N__22267),
            .I(N__22264));
    InMux I__3809 (
            .O(N__22264),
            .I(N__22261));
    LocalMux I__3808 (
            .O(N__22261),
            .I(N__22258));
    Span4Mux_v I__3807 (
            .O(N__22258),
            .I(N__22255));
    Span4Mux_h I__3806 (
            .O(N__22255),
            .I(N__22251));
    InMux I__3805 (
            .O(N__22254),
            .I(N__22248));
    Odrv4 I__3804 (
            .O(N__22251),
            .I(M_this_ppu_vram_addr_6));
    LocalMux I__3803 (
            .O(N__22248),
            .I(M_this_ppu_vram_addr_6));
    CascadeMux I__3802 (
            .O(N__22243),
            .I(N__22240));
    InMux I__3801 (
            .O(N__22240),
            .I(N__22237));
    LocalMux I__3800 (
            .O(N__22237),
            .I(N__22234));
    Span4Mux_v I__3799 (
            .O(N__22234),
            .I(N__22230));
    CascadeMux I__3798 (
            .O(N__22233),
            .I(N__22226));
    Span4Mux_h I__3797 (
            .O(N__22230),
            .I(N__22221));
    InMux I__3796 (
            .O(N__22229),
            .I(N__22212));
    InMux I__3795 (
            .O(N__22226),
            .I(N__22212));
    InMux I__3794 (
            .O(N__22225),
            .I(N__22212));
    InMux I__3793 (
            .O(N__22224),
            .I(N__22212));
    Odrv4 I__3792 (
            .O(N__22221),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__3791 (
            .O(N__22212),
            .I(M_this_ppu_vram_addr_2));
    CascadeMux I__3790 (
            .O(N__22207),
            .I(N__22204));
    InMux I__3789 (
            .O(N__22204),
            .I(N__22201));
    LocalMux I__3788 (
            .O(N__22201),
            .I(M_this_scroll_qZ0Z_0));
    CascadeMux I__3787 (
            .O(N__22198),
            .I(N__22195));
    InMux I__3786 (
            .O(N__22195),
            .I(N__22192));
    LocalMux I__3785 (
            .O(N__22192),
            .I(N__22189));
    Odrv4 I__3784 (
            .O(N__22189),
            .I(M_this_scroll_qZ0Z_1));
    CascadeMux I__3783 (
            .O(N__22186),
            .I(N__22182));
    InMux I__3782 (
            .O(N__22185),
            .I(N__22175));
    InMux I__3781 (
            .O(N__22182),
            .I(N__22175));
    InMux I__3780 (
            .O(N__22181),
            .I(N__22172));
    InMux I__3779 (
            .O(N__22180),
            .I(N__22169));
    LocalMux I__3778 (
            .O(N__22175),
            .I(N__22166));
    LocalMux I__3777 (
            .O(N__22172),
            .I(N__22161));
    LocalMux I__3776 (
            .O(N__22169),
            .I(N__22157));
    Span4Mux_v I__3775 (
            .O(N__22166),
            .I(N__22154));
    InMux I__3774 (
            .O(N__22165),
            .I(N__22149));
    InMux I__3773 (
            .O(N__22164),
            .I(N__22149));
    Span4Mux_h I__3772 (
            .O(N__22161),
            .I(N__22146));
    InMux I__3771 (
            .O(N__22160),
            .I(N__22143));
    Span4Mux_h I__3770 (
            .O(N__22157),
            .I(N__22136));
    Span4Mux_h I__3769 (
            .O(N__22154),
            .I(N__22136));
    LocalMux I__3768 (
            .O(N__22149),
            .I(N__22136));
    Odrv4 I__3767 (
            .O(N__22146),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    LocalMux I__3766 (
            .O(N__22143),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    Odrv4 I__3765 (
            .O(N__22136),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    InMux I__3764 (
            .O(N__22129),
            .I(N__22126));
    LocalMux I__3763 (
            .O(N__22126),
            .I(N__22123));
    Span4Mux_h I__3762 (
            .O(N__22123),
            .I(N__22120));
    Odrv4 I__3761 (
            .O(N__22120),
            .I(\this_ppu.M_state_q_srsts_1_8 ));
    InMux I__3760 (
            .O(N__22117),
            .I(N__22113));
    InMux I__3759 (
            .O(N__22116),
            .I(N__22110));
    LocalMux I__3758 (
            .O(N__22113),
            .I(N__22107));
    LocalMux I__3757 (
            .O(N__22110),
            .I(\this_ppu.N_1145 ));
    Odrv12 I__3756 (
            .O(N__22107),
            .I(\this_ppu.N_1145 ));
    CascadeMux I__3755 (
            .O(N__22102),
            .I(N__22099));
    InMux I__3754 (
            .O(N__22099),
            .I(N__22095));
    CascadeMux I__3753 (
            .O(N__22098),
            .I(N__22092));
    LocalMux I__3752 (
            .O(N__22095),
            .I(N__22089));
    InMux I__3751 (
            .O(N__22092),
            .I(N__22086));
    Odrv4 I__3750 (
            .O(N__22089),
            .I(\this_ppu.M_screen_y_qZ0Z_7 ));
    LocalMux I__3749 (
            .O(N__22086),
            .I(\this_ppu.M_screen_y_qZ0Z_7 ));
    InMux I__3748 (
            .O(N__22081),
            .I(N__22073));
    InMux I__3747 (
            .O(N__22080),
            .I(N__22073));
    InMux I__3746 (
            .O(N__22079),
            .I(N__22070));
    InMux I__3745 (
            .O(N__22078),
            .I(N__22067));
    LocalMux I__3744 (
            .O(N__22073),
            .I(N__22060));
    LocalMux I__3743 (
            .O(N__22070),
            .I(N__22060));
    LocalMux I__3742 (
            .O(N__22067),
            .I(N__22060));
    Span4Mux_v I__3741 (
            .O(N__22060),
            .I(N__22057));
    Odrv4 I__3740 (
            .O(N__22057),
            .I(\this_ppu.M_screen_y_qZ0Z_1 ));
    InMux I__3739 (
            .O(N__22054),
            .I(N__22051));
    LocalMux I__3738 (
            .O(N__22051),
            .I(N__22048));
    Odrv4 I__3737 (
            .O(N__22048),
            .I(\this_ppu.un3_M_screen_y_d_0_c2 ));
    CascadeMux I__3736 (
            .O(N__22045),
            .I(\this_ppu.un3_M_screen_y_d_0_c2_cascade_ ));
    CascadeMux I__3735 (
            .O(N__22042),
            .I(\this_ppu.un3_M_screen_y_d_0_c4_cascade_ ));
    InMux I__3734 (
            .O(N__22039),
            .I(N__22036));
    LocalMux I__3733 (
            .O(N__22036),
            .I(\this_ppu.un3_M_screen_y_d_0_c6 ));
    CascadeMux I__3732 (
            .O(N__22033),
            .I(N_861_0_cascade_));
    CascadeMux I__3731 (
            .O(N__22030),
            .I(N__22026));
    InMux I__3730 (
            .O(N__22029),
            .I(N__22022));
    InMux I__3729 (
            .O(N__22026),
            .I(N__22017));
    InMux I__3728 (
            .O(N__22025),
            .I(N__22017));
    LocalMux I__3727 (
            .O(N__22022),
            .I(N__22014));
    LocalMux I__3726 (
            .O(N__22017),
            .I(\this_ppu.M_screen_y_qZ0Z_2 ));
    Odrv4 I__3725 (
            .O(N__22014),
            .I(\this_ppu.M_screen_y_qZ0Z_2 ));
    CascadeMux I__3724 (
            .O(N__22009),
            .I(N__22006));
    InMux I__3723 (
            .O(N__22006),
            .I(N__22003));
    LocalMux I__3722 (
            .O(N__22003),
            .I(N__21999));
    InMux I__3721 (
            .O(N__22002),
            .I(N__21996));
    Odrv4 I__3720 (
            .O(N__21999),
            .I(\this_ppu.un3_M_screen_y_d_a_2 ));
    LocalMux I__3719 (
            .O(N__21996),
            .I(\this_ppu.un3_M_screen_y_d_a_2 ));
    CascadeMux I__3718 (
            .O(N__21991),
            .I(N__21988));
    InMux I__3717 (
            .O(N__21988),
            .I(N__21984));
    InMux I__3716 (
            .O(N__21987),
            .I(N__21981));
    LocalMux I__3715 (
            .O(N__21984),
            .I(N__21978));
    LocalMux I__3714 (
            .O(N__21981),
            .I(N__21975));
    Span4Mux_v I__3713 (
            .O(N__21978),
            .I(N__21970));
    Span4Mux_h I__3712 (
            .O(N__21975),
            .I(N__21970));
    Odrv4 I__3711 (
            .O(N__21970),
            .I(\this_ppu.N_762_0 ));
    InMux I__3710 (
            .O(N__21967),
            .I(N__21964));
    LocalMux I__3709 (
            .O(N__21964),
            .I(N__21960));
    InMux I__3708 (
            .O(N__21963),
            .I(N__21957));
    Odrv12 I__3707 (
            .O(N__21960),
            .I(\this_ppu.N_91_0 ));
    LocalMux I__3706 (
            .O(N__21957),
            .I(\this_ppu.N_91_0 ));
    CascadeMux I__3705 (
            .O(N__21952),
            .I(\this_ppu.N_91_0_cascade_ ));
    InMux I__3704 (
            .O(N__21949),
            .I(N__21946));
    LocalMux I__3703 (
            .O(N__21946),
            .I(\this_ppu.un1_M_surface_x_q_c3 ));
    CascadeMux I__3702 (
            .O(N__21943),
            .I(\this_ppu.un1_M_surface_x_q_c3_cascade_ ));
    InMux I__3701 (
            .O(N__21940),
            .I(N__21937));
    LocalMux I__3700 (
            .O(N__21937),
            .I(\this_ppu.un1_M_surface_x_q_c6 ));
    CascadeMux I__3699 (
            .O(N__21934),
            .I(N__21931));
    InMux I__3698 (
            .O(N__21931),
            .I(N__21928));
    LocalMux I__3697 (
            .O(N__21928),
            .I(N__21925));
    Odrv4 I__3696 (
            .O(N__21925),
            .I(\this_ppu.N_1202 ));
    InMux I__3695 (
            .O(N__21922),
            .I(N__21919));
    LocalMux I__3694 (
            .O(N__21919),
            .I(N__21913));
    InMux I__3693 (
            .O(N__21918),
            .I(N__21910));
    InMux I__3692 (
            .O(N__21917),
            .I(N__21905));
    InMux I__3691 (
            .O(N__21916),
            .I(N__21905));
    Span4Mux_v I__3690 (
            .O(N__21913),
            .I(N__21900));
    LocalMux I__3689 (
            .O(N__21910),
            .I(N__21900));
    LocalMux I__3688 (
            .O(N__21905),
            .I(N__21897));
    Span4Mux_h I__3687 (
            .O(N__21900),
            .I(N__21894));
    Odrv4 I__3686 (
            .O(N__21897),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    Odrv4 I__3685 (
            .O(N__21894),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    CascadeMux I__3684 (
            .O(N__21889),
            .I(N__21886));
    InMux I__3683 (
            .O(N__21886),
            .I(N__21882));
    CascadeMux I__3682 (
            .O(N__21885),
            .I(N__21879));
    LocalMux I__3681 (
            .O(N__21882),
            .I(N__21875));
    InMux I__3680 (
            .O(N__21879),
            .I(N__21872));
    InMux I__3679 (
            .O(N__21878),
            .I(N__21869));
    Span4Mux_v I__3678 (
            .O(N__21875),
            .I(N__21866));
    LocalMux I__3677 (
            .O(N__21872),
            .I(N__21863));
    LocalMux I__3676 (
            .O(N__21869),
            .I(N__21860));
    Span4Mux_v I__3675 (
            .O(N__21866),
            .I(N__21857));
    Span4Mux_h I__3674 (
            .O(N__21863),
            .I(N__21853));
    Span12Mux_s7_v I__3673 (
            .O(N__21860),
            .I(N__21850));
    Span4Mux_h I__3672 (
            .O(N__21857),
            .I(N__21847));
    InMux I__3671 (
            .O(N__21856),
            .I(N__21844));
    Span4Mux_v I__3670 (
            .O(N__21853),
            .I(N__21841));
    Odrv12 I__3669 (
            .O(N__21850),
            .I(M_this_status_flags_qZ0Z_0));
    Odrv4 I__3668 (
            .O(N__21847),
            .I(M_this_status_flags_qZ0Z_0));
    LocalMux I__3667 (
            .O(N__21844),
            .I(M_this_status_flags_qZ0Z_0));
    Odrv4 I__3666 (
            .O(N__21841),
            .I(M_this_status_flags_qZ0Z_0));
    InMux I__3665 (
            .O(N__21832),
            .I(N__21829));
    LocalMux I__3664 (
            .O(N__21829),
            .I(\this_ppu.N_1201 ));
    InMux I__3663 (
            .O(N__21826),
            .I(M_this_data_count_q_cry_9));
    InMux I__3662 (
            .O(N__21823),
            .I(M_this_data_count_q_cry_10));
    InMux I__3661 (
            .O(N__21820),
            .I(M_this_data_count_q_cry_11));
    InMux I__3660 (
            .O(N__21817),
            .I(M_this_data_count_q_cry_12));
    CascadeMux I__3659 (
            .O(N__21814),
            .I(N__21811));
    CascadeBuf I__3658 (
            .O(N__21811),
            .I(N__21808));
    CascadeMux I__3657 (
            .O(N__21808),
            .I(N__21804));
    CascadeMux I__3656 (
            .O(N__21807),
            .I(N__21801));
    InMux I__3655 (
            .O(N__21804),
            .I(N__21798));
    InMux I__3654 (
            .O(N__21801),
            .I(N__21795));
    LocalMux I__3653 (
            .O(N__21798),
            .I(N__21792));
    LocalMux I__3652 (
            .O(N__21795),
            .I(M_this_oam_address_qZ0Z_7));
    Odrv12 I__3651 (
            .O(N__21792),
            .I(M_this_oam_address_qZ0Z_7));
    IoInMux I__3650 (
            .O(N__21787),
            .I(N__21784));
    LocalMux I__3649 (
            .O(N__21784),
            .I(N__21781));
    Odrv12 I__3648 (
            .O(N__21781),
            .I(IO_port_data_write_i_m2_i_m2_0));
    IoInMux I__3647 (
            .O(N__21778),
            .I(N__21775));
    LocalMux I__3646 (
            .O(N__21775),
            .I(N__21772));
    IoSpan4Mux I__3645 (
            .O(N__21772),
            .I(N__21769));
    Sp12to4 I__3644 (
            .O(N__21769),
            .I(N__21766));
    Span12Mux_v I__3643 (
            .O(N__21766),
            .I(N__21763));
    Odrv12 I__3642 (
            .O(N__21763),
            .I(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO));
    InMux I__3641 (
            .O(N__21760),
            .I(N__21757));
    LocalMux I__3640 (
            .O(N__21757),
            .I(\this_ppu.M_state_qZ0Z_8 ));
    InMux I__3639 (
            .O(N__21754),
            .I(M_this_data_count_q_cry_0));
    InMux I__3638 (
            .O(N__21751),
            .I(M_this_data_count_q_cry_1));
    InMux I__3637 (
            .O(N__21748),
            .I(M_this_data_count_q_cry_2));
    InMux I__3636 (
            .O(N__21745),
            .I(M_this_data_count_q_cry_3));
    InMux I__3635 (
            .O(N__21742),
            .I(M_this_data_count_q_cry_4));
    InMux I__3634 (
            .O(N__21739),
            .I(M_this_data_count_q_cry_5));
    InMux I__3633 (
            .O(N__21736),
            .I(M_this_data_count_q_cry_6));
    InMux I__3632 (
            .O(N__21733),
            .I(bfn_14_25_0_));
    InMux I__3631 (
            .O(N__21730),
            .I(M_this_data_count_q_cry_8));
    InMux I__3630 (
            .O(N__21727),
            .I(bfn_14_22_0_));
    CascadeMux I__3629 (
            .O(N__21724),
            .I(N__21721));
    CascadeBuf I__3628 (
            .O(N__21721),
            .I(N__21718));
    CascadeMux I__3627 (
            .O(N__21718),
            .I(N__21715));
    InMux I__3626 (
            .O(N__21715),
            .I(N__21712));
    LocalMux I__3625 (
            .O(N__21712),
            .I(N__21709));
    Span4Mux_s2_v I__3624 (
            .O(N__21709),
            .I(N__21706));
    Sp12to4 I__3623 (
            .O(N__21706),
            .I(N__21702));
    InMux I__3622 (
            .O(N__21705),
            .I(N__21699));
    Span12Mux_s6_h I__3621 (
            .O(N__21702),
            .I(N__21696));
    LocalMux I__3620 (
            .O(N__21699),
            .I(N__21693));
    Span12Mux_h I__3619 (
            .O(N__21696),
            .I(N__21690));
    Odrv12 I__3618 (
            .O(N__21693),
            .I(M_this_ppu_map_addr_9));
    Odrv12 I__3617 (
            .O(N__21690),
            .I(M_this_ppu_map_addr_9));
    InMux I__3616 (
            .O(N__21685),
            .I(N__21682));
    LocalMux I__3615 (
            .O(N__21682),
            .I(N__21679));
    Odrv4 I__3614 (
            .O(N__21679),
            .I(\this_ppu.M_screen_y_q_esr_RNI563Q6Z0Z_2 ));
    InMux I__3613 (
            .O(N__21676),
            .I(N__21673));
    LocalMux I__3612 (
            .O(N__21673),
            .I(N__21669));
    InMux I__3611 (
            .O(N__21672),
            .I(N__21666));
    Span4Mux_h I__3610 (
            .O(N__21669),
            .I(N__21661));
    LocalMux I__3609 (
            .O(N__21666),
            .I(N__21661));
    Span4Mux_h I__3608 (
            .O(N__21661),
            .I(N__21658));
    Odrv4 I__3607 (
            .O(N__21658),
            .I(M_this_oam_ram_read_data_23));
    InMux I__3606 (
            .O(N__21655),
            .I(N__21652));
    LocalMux I__3605 (
            .O(N__21652),
            .I(N__21649));
    Span4Mux_h I__3604 (
            .O(N__21649),
            .I(N__21646));
    Span4Mux_h I__3603 (
            .O(N__21646),
            .I(N__21643));
    Odrv4 I__3602 (
            .O(N__21643),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_23 ));
    InMux I__3601 (
            .O(N__21640),
            .I(N__21637));
    LocalMux I__3600 (
            .O(N__21637),
            .I(N__21633));
    InMux I__3599 (
            .O(N__21636),
            .I(N__21630));
    Span4Mux_h I__3598 (
            .O(N__21633),
            .I(N__21627));
    LocalMux I__3597 (
            .O(N__21630),
            .I(N__21624));
    Span4Mux_h I__3596 (
            .O(N__21627),
            .I(N__21621));
    Span4Mux_h I__3595 (
            .O(N__21624),
            .I(N__21618));
    Odrv4 I__3594 (
            .O(N__21621),
            .I(M_this_oam_ram_read_data_1));
    Odrv4 I__3593 (
            .O(N__21618),
            .I(M_this_oam_ram_read_data_1));
    InMux I__3592 (
            .O(N__21613),
            .I(N__21610));
    LocalMux I__3591 (
            .O(N__21610),
            .I(N__21607));
    Span4Mux_h I__3590 (
            .O(N__21607),
            .I(N__21604));
    Span4Mux_v I__3589 (
            .O(N__21604),
            .I(N__21601));
    Odrv4 I__3588 (
            .O(N__21601),
            .I(\this_ppu.oam_cache.N_581_0 ));
    InMux I__3587 (
            .O(N__21598),
            .I(N__21595));
    LocalMux I__3586 (
            .O(N__21595),
            .I(M_this_data_tmp_qZ0Z_13));
    InMux I__3585 (
            .O(N__21592),
            .I(N__21589));
    LocalMux I__3584 (
            .O(N__21589),
            .I(\this_ppu.m13_0_i_1 ));
    InMux I__3583 (
            .O(N__21586),
            .I(N__21582));
    CascadeMux I__3582 (
            .O(N__21585),
            .I(N__21579));
    LocalMux I__3581 (
            .O(N__21582),
            .I(N__21576));
    InMux I__3580 (
            .O(N__21579),
            .I(N__21573));
    Span4Mux_h I__3579 (
            .O(N__21576),
            .I(N__21569));
    LocalMux I__3578 (
            .O(N__21573),
            .I(N__21566));
    InMux I__3577 (
            .O(N__21572),
            .I(N__21563));
    Span4Mux_h I__3576 (
            .O(N__21569),
            .I(N__21560));
    Span4Mux_h I__3575 (
            .O(N__21566),
            .I(N__21557));
    LocalMux I__3574 (
            .O(N__21563),
            .I(\this_ppu.offset_y ));
    Odrv4 I__3573 (
            .O(N__21560),
            .I(\this_ppu.offset_y ));
    Odrv4 I__3572 (
            .O(N__21557),
            .I(\this_ppu.offset_y ));
    InMux I__3571 (
            .O(N__21550),
            .I(\this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO ));
    InMux I__3570 (
            .O(N__21547),
            .I(N__21544));
    LocalMux I__3569 (
            .O(N__21544),
            .I(\this_ppu.M_screen_y_q_esr_RNI453Q6Z0Z_1 ));
    CascadeMux I__3568 (
            .O(N__21541),
            .I(N__21537));
    CascadeMux I__3567 (
            .O(N__21540),
            .I(N__21534));
    InMux I__3566 (
            .O(N__21537),
            .I(N__21531));
    InMux I__3565 (
            .O(N__21534),
            .I(N__21528));
    LocalMux I__3564 (
            .O(N__21531),
            .I(N__21525));
    LocalMux I__3563 (
            .O(N__21528),
            .I(N__21522));
    Span12Mux_h I__3562 (
            .O(N__21525),
            .I(N__21519));
    Span4Mux_h I__3561 (
            .O(N__21522),
            .I(N__21516));
    Odrv12 I__3560 (
            .O(N__21519),
            .I(\this_ppu.M_surface_y_qZ0Z_1 ));
    Odrv4 I__3559 (
            .O(N__21516),
            .I(\this_ppu.M_surface_y_qZ0Z_1 ));
    InMux I__3558 (
            .O(N__21511),
            .I(\this_ppu.un1_M_surface_y_d_cry_0 ));
    CascadeMux I__3557 (
            .O(N__21508),
            .I(N__21505));
    InMux I__3556 (
            .O(N__21505),
            .I(N__21501));
    CascadeMux I__3555 (
            .O(N__21504),
            .I(N__21498));
    LocalMux I__3554 (
            .O(N__21501),
            .I(N__21495));
    InMux I__3553 (
            .O(N__21498),
            .I(N__21492));
    Span4Mux_v I__3552 (
            .O(N__21495),
            .I(N__21489));
    LocalMux I__3551 (
            .O(N__21492),
            .I(N__21486));
    Span4Mux_h I__3550 (
            .O(N__21489),
            .I(N__21481));
    Span4Mux_v I__3549 (
            .O(N__21486),
            .I(N__21481));
    Odrv4 I__3548 (
            .O(N__21481),
            .I(\this_ppu.M_surface_y_qZ0Z_2 ));
    InMux I__3547 (
            .O(N__21478),
            .I(\this_ppu.un1_M_surface_y_d_cry_1 ));
    CascadeMux I__3546 (
            .O(N__21475),
            .I(N__21472));
    CascadeBuf I__3545 (
            .O(N__21472),
            .I(N__21469));
    CascadeMux I__3544 (
            .O(N__21469),
            .I(N__21465));
    CascadeMux I__3543 (
            .O(N__21468),
            .I(N__21462));
    InMux I__3542 (
            .O(N__21465),
            .I(N__21459));
    InMux I__3541 (
            .O(N__21462),
            .I(N__21456));
    LocalMux I__3540 (
            .O(N__21459),
            .I(N__21453));
    LocalMux I__3539 (
            .O(N__21456),
            .I(N__21450));
    Sp12to4 I__3538 (
            .O(N__21453),
            .I(N__21447));
    Span4Mux_v I__3537 (
            .O(N__21450),
            .I(N__21444));
    Span12Mux_s11_v I__3536 (
            .O(N__21447),
            .I(N__21441));
    Odrv4 I__3535 (
            .O(N__21444),
            .I(M_this_ppu_map_addr_5));
    Odrv12 I__3534 (
            .O(N__21441),
            .I(M_this_ppu_map_addr_5));
    InMux I__3533 (
            .O(N__21436),
            .I(\this_ppu.un1_M_surface_y_d_cry_2 ));
    InMux I__3532 (
            .O(N__21433),
            .I(N__21430));
    LocalMux I__3531 (
            .O(N__21430),
            .I(\this_ppu.M_screen_y_q_RNI8FJF7Z0Z_4 ));
    CascadeMux I__3530 (
            .O(N__21427),
            .I(N__21424));
    CascadeBuf I__3529 (
            .O(N__21424),
            .I(N__21420));
    CascadeMux I__3528 (
            .O(N__21423),
            .I(N__21417));
    CascadeMux I__3527 (
            .O(N__21420),
            .I(N__21414));
    InMux I__3526 (
            .O(N__21417),
            .I(N__21411));
    InMux I__3525 (
            .O(N__21414),
            .I(N__21408));
    LocalMux I__3524 (
            .O(N__21411),
            .I(N__21405));
    LocalMux I__3523 (
            .O(N__21408),
            .I(N__21402));
    Span4Mux_v I__3522 (
            .O(N__21405),
            .I(N__21399));
    Span12Mux_s11_v I__3521 (
            .O(N__21402),
            .I(N__21396));
    Odrv4 I__3520 (
            .O(N__21399),
            .I(M_this_ppu_map_addr_6));
    Odrv12 I__3519 (
            .O(N__21396),
            .I(M_this_ppu_map_addr_6));
    InMux I__3518 (
            .O(N__21391),
            .I(\this_ppu.un1_M_surface_y_d_cry_3 ));
    CascadeMux I__3517 (
            .O(N__21388),
            .I(N__21385));
    CascadeBuf I__3516 (
            .O(N__21385),
            .I(N__21382));
    CascadeMux I__3515 (
            .O(N__21382),
            .I(N__21379));
    InMux I__3514 (
            .O(N__21379),
            .I(N__21375));
    InMux I__3513 (
            .O(N__21378),
            .I(N__21372));
    LocalMux I__3512 (
            .O(N__21375),
            .I(N__21369));
    LocalMux I__3511 (
            .O(N__21372),
            .I(N__21366));
    Span4Mux_h I__3510 (
            .O(N__21369),
            .I(N__21363));
    Span4Mux_h I__3509 (
            .O(N__21366),
            .I(N__21360));
    Sp12to4 I__3508 (
            .O(N__21363),
            .I(N__21357));
    Span4Mux_h I__3507 (
            .O(N__21360),
            .I(N__21354));
    Span12Mux_s11_v I__3506 (
            .O(N__21357),
            .I(N__21351));
    Odrv4 I__3505 (
            .O(N__21354),
            .I(M_this_ppu_map_addr_7));
    Odrv12 I__3504 (
            .O(N__21351),
            .I(M_this_ppu_map_addr_7));
    InMux I__3503 (
            .O(N__21346),
            .I(\this_ppu.un1_M_surface_y_d_cry_4 ));
    CascadeMux I__3502 (
            .O(N__21343),
            .I(N__21340));
    CascadeBuf I__3501 (
            .O(N__21340),
            .I(N__21337));
    CascadeMux I__3500 (
            .O(N__21337),
            .I(N__21334));
    InMux I__3499 (
            .O(N__21334),
            .I(N__21331));
    LocalMux I__3498 (
            .O(N__21331),
            .I(N__21327));
    InMux I__3497 (
            .O(N__21330),
            .I(N__21324));
    Sp12to4 I__3496 (
            .O(N__21327),
            .I(N__21321));
    LocalMux I__3495 (
            .O(N__21324),
            .I(N__21318));
    Span12Mux_s4_v I__3494 (
            .O(N__21321),
            .I(N__21315));
    Span4Mux_h I__3493 (
            .O(N__21318),
            .I(N__21312));
    Span12Mux_h I__3492 (
            .O(N__21315),
            .I(N__21309));
    Odrv4 I__3491 (
            .O(N__21312),
            .I(M_this_ppu_map_addr_8));
    Odrv12 I__3490 (
            .O(N__21309),
            .I(M_this_ppu_map_addr_8));
    InMux I__3489 (
            .O(N__21304),
            .I(\this_ppu.un1_M_surface_y_d_cry_5 ));
    InMux I__3488 (
            .O(N__21301),
            .I(N__21298));
    LocalMux I__3487 (
            .O(N__21298),
            .I(N__21295));
    Odrv4 I__3486 (
            .O(N__21295),
            .I(\this_ppu.M_oam_cache_read_data_i_12 ));
    InMux I__3485 (
            .O(N__21292),
            .I(N__21289));
    LocalMux I__3484 (
            .O(N__21289),
            .I(\this_ppu.offset_x_4 ));
    InMux I__3483 (
            .O(N__21286),
            .I(\this_ppu.offset_x_cry_3 ));
    InMux I__3482 (
            .O(N__21283),
            .I(N__21280));
    LocalMux I__3481 (
            .O(N__21280),
            .I(\this_ppu.M_oam_cache_read_data_i_13 ));
    CascadeMux I__3480 (
            .O(N__21277),
            .I(N__21274));
    InMux I__3479 (
            .O(N__21274),
            .I(N__21271));
    LocalMux I__3478 (
            .O(N__21271),
            .I(\this_ppu.offset_x_5 ));
    InMux I__3477 (
            .O(N__21268),
            .I(\this_ppu.offset_x_cry_4 ));
    InMux I__3476 (
            .O(N__21265),
            .I(N__21262));
    LocalMux I__3475 (
            .O(N__21262),
            .I(\this_ppu.M_oam_cache_read_data_i_14 ));
    CascadeMux I__3474 (
            .O(N__21259),
            .I(N__21256));
    CascadeBuf I__3473 (
            .O(N__21256),
            .I(N__21253));
    CascadeMux I__3472 (
            .O(N__21253),
            .I(N__21250));
    InMux I__3471 (
            .O(N__21250),
            .I(N__21247));
    LocalMux I__3470 (
            .O(N__21247),
            .I(N__21244));
    Span4Mux_s2_v I__3469 (
            .O(N__21244),
            .I(N__21239));
    InMux I__3468 (
            .O(N__21243),
            .I(N__21235));
    CascadeMux I__3467 (
            .O(N__21242),
            .I(N__21232));
    Sp12to4 I__3466 (
            .O(N__21239),
            .I(N__21229));
    InMux I__3465 (
            .O(N__21238),
            .I(N__21226));
    LocalMux I__3464 (
            .O(N__21235),
            .I(N__21223));
    InMux I__3463 (
            .O(N__21232),
            .I(N__21220));
    Span12Mux_v I__3462 (
            .O(N__21229),
            .I(N__21217));
    LocalMux I__3461 (
            .O(N__21226),
            .I(M_this_ppu_map_addr_3));
    Odrv12 I__3460 (
            .O(N__21223),
            .I(M_this_ppu_map_addr_3));
    LocalMux I__3459 (
            .O(N__21220),
            .I(M_this_ppu_map_addr_3));
    Odrv12 I__3458 (
            .O(N__21217),
            .I(M_this_ppu_map_addr_3));
    InMux I__3457 (
            .O(N__21208),
            .I(N__21205));
    LocalMux I__3456 (
            .O(N__21205),
            .I(\this_ppu.offset_x_6 ));
    InMux I__3455 (
            .O(N__21202),
            .I(\this_ppu.offset_x_cry_5 ));
    InMux I__3454 (
            .O(N__21199),
            .I(N__21196));
    LocalMux I__3453 (
            .O(N__21196),
            .I(N__21193));
    Span4Mux_v I__3452 (
            .O(N__21193),
            .I(N__21190));
    Odrv4 I__3451 (
            .O(N__21190),
            .I(\this_ppu.M_oam_cache_read_data_15 ));
    CascadeMux I__3450 (
            .O(N__21187),
            .I(N__21184));
    CascadeBuf I__3449 (
            .O(N__21184),
            .I(N__21181));
    CascadeMux I__3448 (
            .O(N__21181),
            .I(N__21178));
    InMux I__3447 (
            .O(N__21178),
            .I(N__21175));
    LocalMux I__3446 (
            .O(N__21175),
            .I(N__21172));
    Span4Mux_v I__3445 (
            .O(N__21172),
            .I(N__21168));
    InMux I__3444 (
            .O(N__21171),
            .I(N__21164));
    Sp12to4 I__3443 (
            .O(N__21168),
            .I(N__21161));
    InMux I__3442 (
            .O(N__21167),
            .I(N__21158));
    LocalMux I__3441 (
            .O(N__21164),
            .I(N__21153));
    Span12Mux_h I__3440 (
            .O(N__21161),
            .I(N__21153));
    LocalMux I__3439 (
            .O(N__21158),
            .I(M_this_ppu_map_addr_4));
    Odrv12 I__3438 (
            .O(N__21153),
            .I(M_this_ppu_map_addr_4));
    InMux I__3437 (
            .O(N__21148),
            .I(bfn_14_20_0_));
    InMux I__3436 (
            .O(N__21145),
            .I(N__21142));
    LocalMux I__3435 (
            .O(N__21142),
            .I(\this_ppu.offset_x_7 ));
    CascadeMux I__3434 (
            .O(N__21139),
            .I(N__21136));
    InMux I__3433 (
            .O(N__21136),
            .I(N__21129));
    CascadeMux I__3432 (
            .O(N__21135),
            .I(N__21123));
    CascadeMux I__3431 (
            .O(N__21134),
            .I(N__21120));
    CascadeMux I__3430 (
            .O(N__21133),
            .I(N__21117));
    CascadeMux I__3429 (
            .O(N__21132),
            .I(N__21113));
    LocalMux I__3428 (
            .O(N__21129),
            .I(N__21108));
    CascadeMux I__3427 (
            .O(N__21128),
            .I(N__21105));
    CascadeMux I__3426 (
            .O(N__21127),
            .I(N__21100));
    CascadeMux I__3425 (
            .O(N__21126),
            .I(N__21097));
    InMux I__3424 (
            .O(N__21123),
            .I(N__21094));
    InMux I__3423 (
            .O(N__21120),
            .I(N__21091));
    InMux I__3422 (
            .O(N__21117),
            .I(N__21088));
    CascadeMux I__3421 (
            .O(N__21116),
            .I(N__21085));
    InMux I__3420 (
            .O(N__21113),
            .I(N__21079));
    CascadeMux I__3419 (
            .O(N__21112),
            .I(N__21076));
    CascadeMux I__3418 (
            .O(N__21111),
            .I(N__21073));
    Span4Mux_h I__3417 (
            .O(N__21108),
            .I(N__21070));
    InMux I__3416 (
            .O(N__21105),
            .I(N__21067));
    CascadeMux I__3415 (
            .O(N__21104),
            .I(N__21064));
    CascadeMux I__3414 (
            .O(N__21103),
            .I(N__21061));
    InMux I__3413 (
            .O(N__21100),
            .I(N__21058));
    InMux I__3412 (
            .O(N__21097),
            .I(N__21055));
    LocalMux I__3411 (
            .O(N__21094),
            .I(N__21052));
    LocalMux I__3410 (
            .O(N__21091),
            .I(N__21047));
    LocalMux I__3409 (
            .O(N__21088),
            .I(N__21047));
    InMux I__3408 (
            .O(N__21085),
            .I(N__21044));
    CascadeMux I__3407 (
            .O(N__21084),
            .I(N__21041));
    CascadeMux I__3406 (
            .O(N__21083),
            .I(N__21038));
    CascadeMux I__3405 (
            .O(N__21082),
            .I(N__21035));
    LocalMux I__3404 (
            .O(N__21079),
            .I(N__21032));
    InMux I__3403 (
            .O(N__21076),
            .I(N__21029));
    InMux I__3402 (
            .O(N__21073),
            .I(N__21026));
    IoSpan4Mux I__3401 (
            .O(N__21070),
            .I(N__21023));
    LocalMux I__3400 (
            .O(N__21067),
            .I(N__21020));
    InMux I__3399 (
            .O(N__21064),
            .I(N__21017));
    InMux I__3398 (
            .O(N__21061),
            .I(N__21014));
    LocalMux I__3397 (
            .O(N__21058),
            .I(N__21011));
    LocalMux I__3396 (
            .O(N__21055),
            .I(N__21002));
    Span4Mux_v I__3395 (
            .O(N__21052),
            .I(N__21002));
    Span4Mux_v I__3394 (
            .O(N__21047),
            .I(N__21002));
    LocalMux I__3393 (
            .O(N__21044),
            .I(N__21002));
    InMux I__3392 (
            .O(N__21041),
            .I(N__20999));
    InMux I__3391 (
            .O(N__21038),
            .I(N__20996));
    InMux I__3390 (
            .O(N__21035),
            .I(N__20993));
    Span4Mux_v I__3389 (
            .O(N__21032),
            .I(N__20990));
    LocalMux I__3388 (
            .O(N__21029),
            .I(N__20985));
    LocalMux I__3387 (
            .O(N__21026),
            .I(N__20985));
    IoSpan4Mux I__3386 (
            .O(N__21023),
            .I(N__20982));
    Span4Mux_h I__3385 (
            .O(N__21020),
            .I(N__20979));
    LocalMux I__3384 (
            .O(N__21017),
            .I(N__20974));
    LocalMux I__3383 (
            .O(N__21014),
            .I(N__20974));
    Span4Mux_v I__3382 (
            .O(N__21011),
            .I(N__20971));
    Span4Mux_v I__3381 (
            .O(N__21002),
            .I(N__20966));
    LocalMux I__3380 (
            .O(N__20999),
            .I(N__20966));
    LocalMux I__3379 (
            .O(N__20996),
            .I(N__20961));
    LocalMux I__3378 (
            .O(N__20993),
            .I(N__20961));
    Span4Mux_h I__3377 (
            .O(N__20990),
            .I(N__20956));
    Span4Mux_v I__3376 (
            .O(N__20985),
            .I(N__20956));
    Span4Mux_s3_v I__3375 (
            .O(N__20982),
            .I(N__20951));
    Span4Mux_h I__3374 (
            .O(N__20979),
            .I(N__20951));
    Span4Mux_v I__3373 (
            .O(N__20974),
            .I(N__20948));
    Span4Mux_h I__3372 (
            .O(N__20971),
            .I(N__20945));
    Span4Mux_v I__3371 (
            .O(N__20966),
            .I(N__20940));
    Span4Mux_v I__3370 (
            .O(N__20961),
            .I(N__20940));
    Sp12to4 I__3369 (
            .O(N__20956),
            .I(N__20937));
    Span4Mux_v I__3368 (
            .O(N__20951),
            .I(N__20934));
    Sp12to4 I__3367 (
            .O(N__20948),
            .I(N__20931));
    Sp12to4 I__3366 (
            .O(N__20945),
            .I(N__20926));
    Sp12to4 I__3365 (
            .O(N__20940),
            .I(N__20926));
    Span12Mux_h I__3364 (
            .O(N__20937),
            .I(N__20923));
    Span4Mux_v I__3363 (
            .O(N__20934),
            .I(N__20920));
    Span12Mux_h I__3362 (
            .O(N__20931),
            .I(N__20915));
    Span12Mux_h I__3361 (
            .O(N__20926),
            .I(N__20915));
    Span12Mux_v I__3360 (
            .O(N__20923),
            .I(N__20912));
    Odrv4 I__3359 (
            .O(N__20920),
            .I(M_this_ppu_spr_addr_0));
    Odrv12 I__3358 (
            .O(N__20915),
            .I(M_this_ppu_spr_addr_0));
    Odrv12 I__3357 (
            .O(N__20912),
            .I(M_this_ppu_spr_addr_0));
    CascadeMux I__3356 (
            .O(N__20905),
            .I(N__20902));
    InMux I__3355 (
            .O(N__20902),
            .I(N__20898));
    InMux I__3354 (
            .O(N__20901),
            .I(N__20895));
    LocalMux I__3353 (
            .O(N__20898),
            .I(\this_ppu.M_oam_cache_read_data_8 ));
    LocalMux I__3352 (
            .O(N__20895),
            .I(\this_ppu.M_oam_cache_read_data_8 ));
    InMux I__3351 (
            .O(N__20890),
            .I(N__20887));
    LocalMux I__3350 (
            .O(N__20887),
            .I(\this_ppu.M_oam_cache_read_data_i_8 ));
    InMux I__3349 (
            .O(N__20884),
            .I(N__20881));
    LocalMux I__3348 (
            .O(N__20881),
            .I(\this_ppu.M_oam_cache_read_data_i_9 ));
    CascadeMux I__3347 (
            .O(N__20878),
            .I(N__20875));
    InMux I__3346 (
            .O(N__20875),
            .I(N__20871));
    CascadeMux I__3345 (
            .O(N__20874),
            .I(N__20868));
    LocalMux I__3344 (
            .O(N__20871),
            .I(N__20864));
    InMux I__3343 (
            .O(N__20868),
            .I(N__20861));
    CascadeMux I__3342 (
            .O(N__20867),
            .I(N__20858));
    Span4Mux_s2_v I__3341 (
            .O(N__20864),
            .I(N__20852));
    LocalMux I__3340 (
            .O(N__20861),
            .I(N__20852));
    InMux I__3339 (
            .O(N__20858),
            .I(N__20849));
    CascadeMux I__3338 (
            .O(N__20857),
            .I(N__20846));
    Span4Mux_v I__3337 (
            .O(N__20852),
            .I(N__20840));
    LocalMux I__3336 (
            .O(N__20849),
            .I(N__20840));
    InMux I__3335 (
            .O(N__20846),
            .I(N__20837));
    CascadeMux I__3334 (
            .O(N__20845),
            .I(N__20834));
    Span4Mux_h I__3333 (
            .O(N__20840),
            .I(N__20824));
    LocalMux I__3332 (
            .O(N__20837),
            .I(N__20824));
    InMux I__3331 (
            .O(N__20834),
            .I(N__20821));
    CascadeMux I__3330 (
            .O(N__20833),
            .I(N__20818));
    CascadeMux I__3329 (
            .O(N__20832),
            .I(N__20814));
    CascadeMux I__3328 (
            .O(N__20831),
            .I(N__20811));
    CascadeMux I__3327 (
            .O(N__20830),
            .I(N__20807));
    CascadeMux I__3326 (
            .O(N__20829),
            .I(N__20804));
    Span4Mux_v I__3325 (
            .O(N__20824),
            .I(N__20797));
    LocalMux I__3324 (
            .O(N__20821),
            .I(N__20797));
    InMux I__3323 (
            .O(N__20818),
            .I(N__20794));
    CascadeMux I__3322 (
            .O(N__20817),
            .I(N__20791));
    InMux I__3321 (
            .O(N__20814),
            .I(N__20787));
    InMux I__3320 (
            .O(N__20811),
            .I(N__20784));
    CascadeMux I__3319 (
            .O(N__20810),
            .I(N__20781));
    InMux I__3318 (
            .O(N__20807),
            .I(N__20778));
    InMux I__3317 (
            .O(N__20804),
            .I(N__20775));
    CascadeMux I__3316 (
            .O(N__20803),
            .I(N__20772));
    CascadeMux I__3315 (
            .O(N__20802),
            .I(N__20769));
    Span4Mux_h I__3314 (
            .O(N__20797),
            .I(N__20764));
    LocalMux I__3313 (
            .O(N__20794),
            .I(N__20764));
    InMux I__3312 (
            .O(N__20791),
            .I(N__20761));
    CascadeMux I__3311 (
            .O(N__20790),
            .I(N__20758));
    LocalMux I__3310 (
            .O(N__20787),
            .I(N__20752));
    LocalMux I__3309 (
            .O(N__20784),
            .I(N__20752));
    InMux I__3308 (
            .O(N__20781),
            .I(N__20749));
    LocalMux I__3307 (
            .O(N__20778),
            .I(N__20744));
    LocalMux I__3306 (
            .O(N__20775),
            .I(N__20744));
    InMux I__3305 (
            .O(N__20772),
            .I(N__20741));
    InMux I__3304 (
            .O(N__20769),
            .I(N__20738));
    Span4Mux_v I__3303 (
            .O(N__20764),
            .I(N__20733));
    LocalMux I__3302 (
            .O(N__20761),
            .I(N__20733));
    InMux I__3301 (
            .O(N__20758),
            .I(N__20730));
    CascadeMux I__3300 (
            .O(N__20757),
            .I(N__20727));
    Span4Mux_v I__3299 (
            .O(N__20752),
            .I(N__20722));
    LocalMux I__3298 (
            .O(N__20749),
            .I(N__20722));
    Span4Mux_v I__3297 (
            .O(N__20744),
            .I(N__20715));
    LocalMux I__3296 (
            .O(N__20741),
            .I(N__20715));
    LocalMux I__3295 (
            .O(N__20738),
            .I(N__20715));
    Span4Mux_h I__3294 (
            .O(N__20733),
            .I(N__20710));
    LocalMux I__3293 (
            .O(N__20730),
            .I(N__20710));
    InMux I__3292 (
            .O(N__20727),
            .I(N__20707));
    Span4Mux_v I__3291 (
            .O(N__20722),
            .I(N__20704));
    Span4Mux_v I__3290 (
            .O(N__20715),
            .I(N__20697));
    Span4Mux_v I__3289 (
            .O(N__20710),
            .I(N__20697));
    LocalMux I__3288 (
            .O(N__20707),
            .I(N__20697));
    Span4Mux_h I__3287 (
            .O(N__20704),
            .I(N__20694));
    Span4Mux_h I__3286 (
            .O(N__20697),
            .I(N__20691));
    Span4Mux_v I__3285 (
            .O(N__20694),
            .I(N__20688));
    Span4Mux_h I__3284 (
            .O(N__20691),
            .I(N__20685));
    Odrv4 I__3283 (
            .O(N__20688),
            .I(M_this_ppu_spr_addr_1));
    Odrv4 I__3282 (
            .O(N__20685),
            .I(M_this_ppu_spr_addr_1));
    InMux I__3281 (
            .O(N__20680),
            .I(\this_ppu.offset_x_cry_0 ));
    InMux I__3280 (
            .O(N__20677),
            .I(N__20674));
    LocalMux I__3279 (
            .O(N__20674),
            .I(N__20671));
    Span4Mux_h I__3278 (
            .O(N__20671),
            .I(N__20668));
    Odrv4 I__3277 (
            .O(N__20668),
            .I(\this_ppu.M_oam_cache_read_data_i_10 ));
    CascadeMux I__3276 (
            .O(N__20665),
            .I(N__20662));
    InMux I__3275 (
            .O(N__20662),
            .I(N__20658));
    CascadeMux I__3274 (
            .O(N__20661),
            .I(N__20655));
    LocalMux I__3273 (
            .O(N__20658),
            .I(N__20649));
    InMux I__3272 (
            .O(N__20655),
            .I(N__20646));
    CascadeMux I__3271 (
            .O(N__20654),
            .I(N__20643));
    CascadeMux I__3270 (
            .O(N__20653),
            .I(N__20636));
    CascadeMux I__3269 (
            .O(N__20652),
            .I(N__20633));
    Span4Mux_h I__3268 (
            .O(N__20649),
            .I(N__20627));
    LocalMux I__3267 (
            .O(N__20646),
            .I(N__20627));
    InMux I__3266 (
            .O(N__20643),
            .I(N__20624));
    CascadeMux I__3265 (
            .O(N__20642),
            .I(N__20621));
    CascadeMux I__3264 (
            .O(N__20641),
            .I(N__20617));
    CascadeMux I__3263 (
            .O(N__20640),
            .I(N__20614));
    CascadeMux I__3262 (
            .O(N__20639),
            .I(N__20611));
    InMux I__3261 (
            .O(N__20636),
            .I(N__20606));
    InMux I__3260 (
            .O(N__20633),
            .I(N__20602));
    CascadeMux I__3259 (
            .O(N__20632),
            .I(N__20599));
    Span4Mux_v I__3258 (
            .O(N__20627),
            .I(N__20594));
    LocalMux I__3257 (
            .O(N__20624),
            .I(N__20594));
    InMux I__3256 (
            .O(N__20621),
            .I(N__20591));
    CascadeMux I__3255 (
            .O(N__20620),
            .I(N__20588));
    InMux I__3254 (
            .O(N__20617),
            .I(N__20585));
    InMux I__3253 (
            .O(N__20614),
            .I(N__20582));
    InMux I__3252 (
            .O(N__20611),
            .I(N__20579));
    CascadeMux I__3251 (
            .O(N__20610),
            .I(N__20576));
    CascadeMux I__3250 (
            .O(N__20609),
            .I(N__20573));
    LocalMux I__3249 (
            .O(N__20606),
            .I(N__20569));
    CascadeMux I__3248 (
            .O(N__20605),
            .I(N__20566));
    LocalMux I__3247 (
            .O(N__20602),
            .I(N__20562));
    InMux I__3246 (
            .O(N__20599),
            .I(N__20559));
    Span4Mux_h I__3245 (
            .O(N__20594),
            .I(N__20554));
    LocalMux I__3244 (
            .O(N__20591),
            .I(N__20554));
    InMux I__3243 (
            .O(N__20588),
            .I(N__20551));
    LocalMux I__3242 (
            .O(N__20585),
            .I(N__20548));
    LocalMux I__3241 (
            .O(N__20582),
            .I(N__20545));
    LocalMux I__3240 (
            .O(N__20579),
            .I(N__20542));
    InMux I__3239 (
            .O(N__20576),
            .I(N__20539));
    InMux I__3238 (
            .O(N__20573),
            .I(N__20536));
    CascadeMux I__3237 (
            .O(N__20572),
            .I(N__20533));
    Span4Mux_v I__3236 (
            .O(N__20569),
            .I(N__20530));
    InMux I__3235 (
            .O(N__20566),
            .I(N__20527));
    CascadeMux I__3234 (
            .O(N__20565),
            .I(N__20524));
    Span4Mux_h I__3233 (
            .O(N__20562),
            .I(N__20521));
    LocalMux I__3232 (
            .O(N__20559),
            .I(N__20518));
    Span4Mux_v I__3231 (
            .O(N__20554),
            .I(N__20513));
    LocalMux I__3230 (
            .O(N__20551),
            .I(N__20513));
    Span4Mux_v I__3229 (
            .O(N__20548),
            .I(N__20504));
    Span4Mux_v I__3228 (
            .O(N__20545),
            .I(N__20504));
    Span4Mux_h I__3227 (
            .O(N__20542),
            .I(N__20504));
    LocalMux I__3226 (
            .O(N__20539),
            .I(N__20504));
    LocalMux I__3225 (
            .O(N__20536),
            .I(N__20501));
    InMux I__3224 (
            .O(N__20533),
            .I(N__20498));
    Sp12to4 I__3223 (
            .O(N__20530),
            .I(N__20493));
    LocalMux I__3222 (
            .O(N__20527),
            .I(N__20493));
    InMux I__3221 (
            .O(N__20524),
            .I(N__20490));
    Span4Mux_v I__3220 (
            .O(N__20521),
            .I(N__20485));
    Span4Mux_h I__3219 (
            .O(N__20518),
            .I(N__20485));
    Span4Mux_h I__3218 (
            .O(N__20513),
            .I(N__20482));
    Span4Mux_v I__3217 (
            .O(N__20504),
            .I(N__20475));
    Span4Mux_v I__3216 (
            .O(N__20501),
            .I(N__20475));
    LocalMux I__3215 (
            .O(N__20498),
            .I(N__20475));
    Span12Mux_h I__3214 (
            .O(N__20493),
            .I(N__20472));
    LocalMux I__3213 (
            .O(N__20490),
            .I(N__20469));
    Span4Mux_h I__3212 (
            .O(N__20485),
            .I(N__20466));
    Span4Mux_v I__3211 (
            .O(N__20482),
            .I(N__20461));
    Span4Mux_h I__3210 (
            .O(N__20475),
            .I(N__20461));
    Span12Mux_v I__3209 (
            .O(N__20472),
            .I(N__20454));
    Span12Mux_h I__3208 (
            .O(N__20469),
            .I(N__20454));
    Sp12to4 I__3207 (
            .O(N__20466),
            .I(N__20454));
    Span4Mux_h I__3206 (
            .O(N__20461),
            .I(N__20451));
    Odrv12 I__3205 (
            .O(N__20454),
            .I(M_this_ppu_spr_addr_2));
    Odrv4 I__3204 (
            .O(N__20451),
            .I(M_this_ppu_spr_addr_2));
    InMux I__3203 (
            .O(N__20446),
            .I(\this_ppu.offset_x_cry_1 ));
    InMux I__3202 (
            .O(N__20443),
            .I(N__20440));
    LocalMux I__3201 (
            .O(N__20440),
            .I(\this_ppu.M_oam_cache_read_data_i_11 ));
    InMux I__3200 (
            .O(N__20437),
            .I(N__20434));
    LocalMux I__3199 (
            .O(N__20434),
            .I(\this_ppu.m68_0_o2_0 ));
    InMux I__3198 (
            .O(N__20431),
            .I(\this_ppu.offset_x_cry_2 ));
    InMux I__3197 (
            .O(N__20428),
            .I(N__20425));
    LocalMux I__3196 (
            .O(N__20425),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__3195 (
            .O(N__20422),
            .I(N__20413));
    InMux I__3194 (
            .O(N__20421),
            .I(N__20413));
    InMux I__3193 (
            .O(N__20420),
            .I(N__20413));
    LocalMux I__3192 (
            .O(N__20413),
            .I(N__20409));
    InMux I__3191 (
            .O(N__20412),
            .I(N__20406));
    Span4Mux_h I__3190 (
            .O(N__20409),
            .I(N__20403));
    LocalMux I__3189 (
            .O(N__20406),
            .I(N__20400));
    Span4Mux_v I__3188 (
            .O(N__20403),
            .I(N__20397));
    Span12Mux_h I__3187 (
            .O(N__20400),
            .I(N__20394));
    Span4Mux_v I__3186 (
            .O(N__20397),
            .I(N__20391));
    Span12Mux_v I__3185 (
            .O(N__20394),
            .I(N__20388));
    Span4Mux_v I__3184 (
            .O(N__20391),
            .I(N__20385));
    Odrv12 I__3183 (
            .O(N__20388),
            .I(rst_n_c));
    Odrv4 I__3182 (
            .O(N__20385),
            .I(rst_n_c));
    InMux I__3181 (
            .O(N__20380),
            .I(N__20377));
    LocalMux I__3180 (
            .O(N__20377),
            .I(N__20374));
    Odrv4 I__3179 (
            .O(N__20374),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    CascadeMux I__3178 (
            .O(N__20371),
            .I(N__20367));
    CascadeMux I__3177 (
            .O(N__20370),
            .I(N__20363));
    InMux I__3176 (
            .O(N__20367),
            .I(N__20360));
    InMux I__3175 (
            .O(N__20366),
            .I(N__20355));
    InMux I__3174 (
            .O(N__20363),
            .I(N__20355));
    LocalMux I__3173 (
            .O(N__20360),
            .I(\this_vga_signals.N_1417 ));
    LocalMux I__3172 (
            .O(N__20355),
            .I(\this_vga_signals.N_1417 ));
    InMux I__3171 (
            .O(N__20350),
            .I(N__20347));
    LocalMux I__3170 (
            .O(N__20347),
            .I(N__20343));
    InMux I__3169 (
            .O(N__20346),
            .I(N__20338));
    Span4Mux_v I__3168 (
            .O(N__20343),
            .I(N__20335));
    InMux I__3167 (
            .O(N__20342),
            .I(N__20332));
    InMux I__3166 (
            .O(N__20341),
            .I(N__20329));
    LocalMux I__3165 (
            .O(N__20338),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    Odrv4 I__3164 (
            .O(N__20335),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    LocalMux I__3163 (
            .O(N__20332),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    LocalMux I__3162 (
            .O(N__20329),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    InMux I__3161 (
            .O(N__20320),
            .I(N__20317));
    LocalMux I__3160 (
            .O(N__20317),
            .I(N__20314));
    Span12Mux_h I__3159 (
            .O(N__20314),
            .I(N__20311));
    Odrv12 I__3158 (
            .O(N__20311),
            .I(\this_vga_ramdac.i2_mux_0 ));
    InMux I__3157 (
            .O(N__20308),
            .I(N__20300));
    InMux I__3156 (
            .O(N__20307),
            .I(N__20297));
    InMux I__3155 (
            .O(N__20306),
            .I(N__20294));
    InMux I__3154 (
            .O(N__20305),
            .I(N__20291));
    InMux I__3153 (
            .O(N__20304),
            .I(N__20286));
    InMux I__3152 (
            .O(N__20303),
            .I(N__20286));
    LocalMux I__3151 (
            .O(N__20300),
            .I(N__20281));
    LocalMux I__3150 (
            .O(N__20297),
            .I(N__20281));
    LocalMux I__3149 (
            .O(N__20294),
            .I(M_pcounter_q_ret_1_RNIOILK7));
    LocalMux I__3148 (
            .O(N__20291),
            .I(M_pcounter_q_ret_1_RNIOILK7));
    LocalMux I__3147 (
            .O(N__20286),
            .I(M_pcounter_q_ret_1_RNIOILK7));
    Odrv4 I__3146 (
            .O(N__20281),
            .I(M_pcounter_q_ret_1_RNIOILK7));
    InMux I__3145 (
            .O(N__20272),
            .I(N__20269));
    LocalMux I__3144 (
            .O(N__20269),
            .I(N__20266));
    Span4Mux_h I__3143 (
            .O(N__20266),
            .I(N__20262));
    CascadeMux I__3142 (
            .O(N__20265),
            .I(N__20259));
    Span4Mux_h I__3141 (
            .O(N__20262),
            .I(N__20256));
    InMux I__3140 (
            .O(N__20259),
            .I(N__20253));
    Odrv4 I__3139 (
            .O(N__20256),
            .I(\this_vga_ramdac.N_3861_reto ));
    LocalMux I__3138 (
            .O(N__20253),
            .I(\this_vga_ramdac.N_3861_reto ));
    InMux I__3137 (
            .O(N__20248),
            .I(N__20245));
    LocalMux I__3136 (
            .O(N__20245),
            .I(N__20242));
    Odrv12 I__3135 (
            .O(N__20242),
            .I(\this_ppu.un1_M_surface_x_q_ac0_11 ));
    InMux I__3134 (
            .O(N__20239),
            .I(N__20236));
    LocalMux I__3133 (
            .O(N__20236),
            .I(M_this_data_tmp_qZ0Z_12));
    InMux I__3132 (
            .O(N__20233),
            .I(N__20230));
    LocalMux I__3131 (
            .O(N__20230),
            .I(M_this_data_tmp_qZ0Z_14));
    InMux I__3130 (
            .O(N__20227),
            .I(N__20224));
    LocalMux I__3129 (
            .O(N__20224),
            .I(M_this_data_tmp_qZ0Z_1));
    InMux I__3128 (
            .O(N__20221),
            .I(N__20218));
    LocalMux I__3127 (
            .O(N__20218),
            .I(N__20215));
    Span4Mux_v I__3126 (
            .O(N__20215),
            .I(N__20212));
    Span4Mux_h I__3125 (
            .O(N__20212),
            .I(N__20209));
    Odrv4 I__3124 (
            .O(N__20209),
            .I(M_this_oam_ram_write_data_22));
    InMux I__3123 (
            .O(N__20206),
            .I(N__20203));
    LocalMux I__3122 (
            .O(N__20203),
            .I(M_this_data_tmp_qZ0Z_22));
    InMux I__3121 (
            .O(N__20200),
            .I(N__20196));
    InMux I__3120 (
            .O(N__20199),
            .I(N__20193));
    LocalMux I__3119 (
            .O(N__20196),
            .I(N__20190));
    LocalMux I__3118 (
            .O(N__20193),
            .I(N__20187));
    Span12Mux_v I__3117 (
            .O(N__20190),
            .I(N__20184));
    Span12Mux_h I__3116 (
            .O(N__20187),
            .I(N__20181));
    Span12Mux_h I__3115 (
            .O(N__20184),
            .I(N__20178));
    Odrv12 I__3114 (
            .O(N__20181),
            .I(M_this_map_ram_read_data_1));
    Odrv12 I__3113 (
            .O(N__20178),
            .I(M_this_map_ram_read_data_1));
    IoInMux I__3112 (
            .O(N__20173),
            .I(N__20170));
    LocalMux I__3111 (
            .O(N__20170),
            .I(N__20167));
    Odrv4 I__3110 (
            .O(N__20167),
            .I(N_724_0));
    InMux I__3109 (
            .O(N__20164),
            .I(N__20161));
    LocalMux I__3108 (
            .O(N__20161),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__3107 (
            .O(N__20158),
            .I(N__20155));
    LocalMux I__3106 (
            .O(N__20155),
            .I(N__20152));
    Span12Mux_h I__3105 (
            .O(N__20152),
            .I(N__20148));
    InMux I__3104 (
            .O(N__20151),
            .I(N__20145));
    Odrv12 I__3103 (
            .O(N__20148),
            .I(\this_ppu.M_oam_cache_read_data_16 ));
    LocalMux I__3102 (
            .O(N__20145),
            .I(\this_ppu.M_oam_cache_read_data_16 ));
    CascadeMux I__3101 (
            .O(N__20140),
            .I(N__20136));
    CascadeMux I__3100 (
            .O(N__20139),
            .I(N__20133));
    InMux I__3099 (
            .O(N__20136),
            .I(N__20125));
    InMux I__3098 (
            .O(N__20133),
            .I(N__20122));
    CascadeMux I__3097 (
            .O(N__20132),
            .I(N__20119));
    CascadeMux I__3096 (
            .O(N__20131),
            .I(N__20108));
    CascadeMux I__3095 (
            .O(N__20130),
            .I(N__20105));
    CascadeMux I__3094 (
            .O(N__20129),
            .I(N__20101));
    CascadeMux I__3093 (
            .O(N__20128),
            .I(N__20098));
    LocalMux I__3092 (
            .O(N__20125),
            .I(N__20093));
    LocalMux I__3091 (
            .O(N__20122),
            .I(N__20093));
    InMux I__3090 (
            .O(N__20119),
            .I(N__20090));
    CascadeMux I__3089 (
            .O(N__20118),
            .I(N__20087));
    CascadeMux I__3088 (
            .O(N__20117),
            .I(N__20084));
    CascadeMux I__3087 (
            .O(N__20116),
            .I(N__20081));
    CascadeMux I__3086 (
            .O(N__20115),
            .I(N__20078));
    CascadeMux I__3085 (
            .O(N__20114),
            .I(N__20075));
    CascadeMux I__3084 (
            .O(N__20113),
            .I(N__20072));
    CascadeMux I__3083 (
            .O(N__20112),
            .I(N__20069));
    CascadeMux I__3082 (
            .O(N__20111),
            .I(N__20066));
    InMux I__3081 (
            .O(N__20108),
            .I(N__20063));
    InMux I__3080 (
            .O(N__20105),
            .I(N__20060));
    CascadeMux I__3079 (
            .O(N__20104),
            .I(N__20057));
    InMux I__3078 (
            .O(N__20101),
            .I(N__20054));
    InMux I__3077 (
            .O(N__20098),
            .I(N__20051));
    Span4Mux_v I__3076 (
            .O(N__20093),
            .I(N__20046));
    LocalMux I__3075 (
            .O(N__20090),
            .I(N__20046));
    InMux I__3074 (
            .O(N__20087),
            .I(N__20043));
    InMux I__3073 (
            .O(N__20084),
            .I(N__20040));
    InMux I__3072 (
            .O(N__20081),
            .I(N__20037));
    InMux I__3071 (
            .O(N__20078),
            .I(N__20034));
    InMux I__3070 (
            .O(N__20075),
            .I(N__20031));
    InMux I__3069 (
            .O(N__20072),
            .I(N__20028));
    InMux I__3068 (
            .O(N__20069),
            .I(N__20025));
    InMux I__3067 (
            .O(N__20066),
            .I(N__20022));
    LocalMux I__3066 (
            .O(N__20063),
            .I(N__20019));
    LocalMux I__3065 (
            .O(N__20060),
            .I(N__20016));
    InMux I__3064 (
            .O(N__20057),
            .I(N__20013));
    LocalMux I__3063 (
            .O(N__20054),
            .I(N__20008));
    LocalMux I__3062 (
            .O(N__20051),
            .I(N__20008));
    Sp12to4 I__3061 (
            .O(N__20046),
            .I(N__19997));
    LocalMux I__3060 (
            .O(N__20043),
            .I(N__19997));
    LocalMux I__3059 (
            .O(N__20040),
            .I(N__19997));
    LocalMux I__3058 (
            .O(N__20037),
            .I(N__19997));
    LocalMux I__3057 (
            .O(N__20034),
            .I(N__19997));
    LocalMux I__3056 (
            .O(N__20031),
            .I(N__19988));
    LocalMux I__3055 (
            .O(N__20028),
            .I(N__19988));
    LocalMux I__3054 (
            .O(N__20025),
            .I(N__19988));
    LocalMux I__3053 (
            .O(N__20022),
            .I(N__19988));
    Span4Mux_s3_v I__3052 (
            .O(N__20019),
            .I(N__19981));
    Span4Mux_h I__3051 (
            .O(N__20016),
            .I(N__19981));
    LocalMux I__3050 (
            .O(N__20013),
            .I(N__19981));
    Span12Mux_s11_v I__3049 (
            .O(N__20008),
            .I(N__19978));
    Span12Mux_v I__3048 (
            .O(N__19997),
            .I(N__19975));
    Span12Mux_v I__3047 (
            .O(N__19988),
            .I(N__19972));
    Span4Mux_v I__3046 (
            .O(N__19981),
            .I(N__19969));
    Span12Mux_h I__3045 (
            .O(N__19978),
            .I(N__19964));
    Span12Mux_h I__3044 (
            .O(N__19975),
            .I(N__19964));
    Span12Mux_h I__3043 (
            .O(N__19972),
            .I(N__19961));
    Span4Mux_h I__3042 (
            .O(N__19969),
            .I(N__19958));
    Odrv12 I__3041 (
            .O(N__19964),
            .I(M_this_ppu_spr_addr_3));
    Odrv12 I__3040 (
            .O(N__19961),
            .I(M_this_ppu_spr_addr_3));
    Odrv4 I__3039 (
            .O(N__19958),
            .I(M_this_ppu_spr_addr_3));
    InMux I__3038 (
            .O(N__19951),
            .I(N__19948));
    LocalMux I__3037 (
            .O(N__19948),
            .I(N__19945));
    Span4Mux_v I__3036 (
            .O(N__19945),
            .I(N__19942));
    Odrv4 I__3035 (
            .O(N__19942),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_2 ));
    CascadeMux I__3034 (
            .O(N__19939),
            .I(N__19933));
    CascadeMux I__3033 (
            .O(N__19938),
            .I(N__19930));
    CascadeMux I__3032 (
            .O(N__19937),
            .I(N__19925));
    CascadeMux I__3031 (
            .O(N__19936),
            .I(N__19919));
    InMux I__3030 (
            .O(N__19933),
            .I(N__19915));
    InMux I__3029 (
            .O(N__19930),
            .I(N__19912));
    CascadeMux I__3028 (
            .O(N__19929),
            .I(N__19909));
    CascadeMux I__3027 (
            .O(N__19928),
            .I(N__19906));
    InMux I__3026 (
            .O(N__19925),
            .I(N__19902));
    CascadeMux I__3025 (
            .O(N__19924),
            .I(N__19899));
    CascadeMux I__3024 (
            .O(N__19923),
            .I(N__19896));
    CascadeMux I__3023 (
            .O(N__19922),
            .I(N__19893));
    InMux I__3022 (
            .O(N__19919),
            .I(N__19890));
    CascadeMux I__3021 (
            .O(N__19918),
            .I(N__19887));
    LocalMux I__3020 (
            .O(N__19915),
            .I(N__19882));
    LocalMux I__3019 (
            .O(N__19912),
            .I(N__19879));
    InMux I__3018 (
            .O(N__19909),
            .I(N__19876));
    InMux I__3017 (
            .O(N__19906),
            .I(N__19873));
    CascadeMux I__3016 (
            .O(N__19905),
            .I(N__19870));
    LocalMux I__3015 (
            .O(N__19902),
            .I(N__19866));
    InMux I__3014 (
            .O(N__19899),
            .I(N__19863));
    InMux I__3013 (
            .O(N__19896),
            .I(N__19860));
    InMux I__3012 (
            .O(N__19893),
            .I(N__19857));
    LocalMux I__3011 (
            .O(N__19890),
            .I(N__19854));
    InMux I__3010 (
            .O(N__19887),
            .I(N__19851));
    CascadeMux I__3009 (
            .O(N__19886),
            .I(N__19848));
    CascadeMux I__3008 (
            .O(N__19885),
            .I(N__19845));
    Span4Mux_v I__3007 (
            .O(N__19882),
            .I(N__19836));
    Span4Mux_v I__3006 (
            .O(N__19879),
            .I(N__19836));
    LocalMux I__3005 (
            .O(N__19876),
            .I(N__19836));
    LocalMux I__3004 (
            .O(N__19873),
            .I(N__19833));
    InMux I__3003 (
            .O(N__19870),
            .I(N__19830));
    CascadeMux I__3002 (
            .O(N__19869),
            .I(N__19827));
    Span4Mux_v I__3001 (
            .O(N__19866),
            .I(N__19822));
    LocalMux I__3000 (
            .O(N__19863),
            .I(N__19822));
    LocalMux I__2999 (
            .O(N__19860),
            .I(N__19819));
    LocalMux I__2998 (
            .O(N__19857),
            .I(N__19816));
    Span4Mux_v I__2997 (
            .O(N__19854),
            .I(N__19811));
    LocalMux I__2996 (
            .O(N__19851),
            .I(N__19811));
    InMux I__2995 (
            .O(N__19848),
            .I(N__19808));
    InMux I__2994 (
            .O(N__19845),
            .I(N__19805));
    CascadeMux I__2993 (
            .O(N__19844),
            .I(N__19802));
    CascadeMux I__2992 (
            .O(N__19843),
            .I(N__19799));
    Span4Mux_v I__2991 (
            .O(N__19836),
            .I(N__19792));
    Span4Mux_h I__2990 (
            .O(N__19833),
            .I(N__19792));
    LocalMux I__2989 (
            .O(N__19830),
            .I(N__19792));
    InMux I__2988 (
            .O(N__19827),
            .I(N__19789));
    Span4Mux_h I__2987 (
            .O(N__19822),
            .I(N__19786));
    Span4Mux_v I__2986 (
            .O(N__19819),
            .I(N__19777));
    Span4Mux_v I__2985 (
            .O(N__19816),
            .I(N__19777));
    Span4Mux_v I__2984 (
            .O(N__19811),
            .I(N__19777));
    LocalMux I__2983 (
            .O(N__19808),
            .I(N__19777));
    LocalMux I__2982 (
            .O(N__19805),
            .I(N__19774));
    InMux I__2981 (
            .O(N__19802),
            .I(N__19771));
    InMux I__2980 (
            .O(N__19799),
            .I(N__19768));
    Span4Mux_v I__2979 (
            .O(N__19792),
            .I(N__19765));
    LocalMux I__2978 (
            .O(N__19789),
            .I(N__19762));
    Span4Mux_v I__2977 (
            .O(N__19786),
            .I(N__19757));
    Span4Mux_h I__2976 (
            .O(N__19777),
            .I(N__19757));
    Span4Mux_s3_v I__2975 (
            .O(N__19774),
            .I(N__19750));
    LocalMux I__2974 (
            .O(N__19771),
            .I(N__19750));
    LocalMux I__2973 (
            .O(N__19768),
            .I(N__19750));
    Sp12to4 I__2972 (
            .O(N__19765),
            .I(N__19745));
    Span12Mux_s7_h I__2971 (
            .O(N__19762),
            .I(N__19745));
    Span4Mux_h I__2970 (
            .O(N__19757),
            .I(N__19742));
    Span4Mux_v I__2969 (
            .O(N__19750),
            .I(N__19739));
    Span12Mux_h I__2968 (
            .O(N__19745),
            .I(N__19736));
    Span4Mux_h I__2967 (
            .O(N__19742),
            .I(N__19733));
    Span4Mux_h I__2966 (
            .O(N__19739),
            .I(N__19730));
    Odrv12 I__2965 (
            .O(N__19736),
            .I(read_data_RNI6RFJ1_2));
    Odrv4 I__2964 (
            .O(N__19733),
            .I(read_data_RNI6RFJ1_2));
    Odrv4 I__2963 (
            .O(N__19730),
            .I(read_data_RNI6RFJ1_2));
    InMux I__2962 (
            .O(N__19723),
            .I(N__19720));
    LocalMux I__2961 (
            .O(N__19720),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_3 ));
    CascadeMux I__2960 (
            .O(N__19717),
            .I(N__19710));
    CascadeMux I__2959 (
            .O(N__19716),
            .I(N__19706));
    CascadeMux I__2958 (
            .O(N__19715),
            .I(N__19701));
    CascadeMux I__2957 (
            .O(N__19714),
            .I(N__19698));
    CascadeMux I__2956 (
            .O(N__19713),
            .I(N__19695));
    InMux I__2955 (
            .O(N__19710),
            .I(N__19689));
    CascadeMux I__2954 (
            .O(N__19709),
            .I(N__19686));
    InMux I__2953 (
            .O(N__19706),
            .I(N__19678));
    CascadeMux I__2952 (
            .O(N__19705),
            .I(N__19675));
    CascadeMux I__2951 (
            .O(N__19704),
            .I(N__19672));
    InMux I__2950 (
            .O(N__19701),
            .I(N__19669));
    InMux I__2949 (
            .O(N__19698),
            .I(N__19666));
    InMux I__2948 (
            .O(N__19695),
            .I(N__19663));
    CascadeMux I__2947 (
            .O(N__19694),
            .I(N__19660));
    CascadeMux I__2946 (
            .O(N__19693),
            .I(N__19657));
    CascadeMux I__2945 (
            .O(N__19692),
            .I(N__19654));
    LocalMux I__2944 (
            .O(N__19689),
            .I(N__19651));
    InMux I__2943 (
            .O(N__19686),
            .I(N__19648));
    CascadeMux I__2942 (
            .O(N__19685),
            .I(N__19645));
    CascadeMux I__2941 (
            .O(N__19684),
            .I(N__19642));
    CascadeMux I__2940 (
            .O(N__19683),
            .I(N__19639));
    CascadeMux I__2939 (
            .O(N__19682),
            .I(N__19636));
    CascadeMux I__2938 (
            .O(N__19681),
            .I(N__19633));
    LocalMux I__2937 (
            .O(N__19678),
            .I(N__19630));
    InMux I__2936 (
            .O(N__19675),
            .I(N__19627));
    InMux I__2935 (
            .O(N__19672),
            .I(N__19624));
    LocalMux I__2934 (
            .O(N__19669),
            .I(N__19617));
    LocalMux I__2933 (
            .O(N__19666),
            .I(N__19617));
    LocalMux I__2932 (
            .O(N__19663),
            .I(N__19617));
    InMux I__2931 (
            .O(N__19660),
            .I(N__19614));
    InMux I__2930 (
            .O(N__19657),
            .I(N__19611));
    InMux I__2929 (
            .O(N__19654),
            .I(N__19608));
    Span4Mux_v I__2928 (
            .O(N__19651),
            .I(N__19603));
    LocalMux I__2927 (
            .O(N__19648),
            .I(N__19603));
    InMux I__2926 (
            .O(N__19645),
            .I(N__19600));
    InMux I__2925 (
            .O(N__19642),
            .I(N__19597));
    InMux I__2924 (
            .O(N__19639),
            .I(N__19594));
    InMux I__2923 (
            .O(N__19636),
            .I(N__19591));
    InMux I__2922 (
            .O(N__19633),
            .I(N__19588));
    Span4Mux_s3_v I__2921 (
            .O(N__19630),
            .I(N__19581));
    LocalMux I__2920 (
            .O(N__19627),
            .I(N__19581));
    LocalMux I__2919 (
            .O(N__19624),
            .I(N__19581));
    Span12Mux_v I__2918 (
            .O(N__19617),
            .I(N__19578));
    LocalMux I__2917 (
            .O(N__19614),
            .I(N__19571));
    LocalMux I__2916 (
            .O(N__19611),
            .I(N__19571));
    LocalMux I__2915 (
            .O(N__19608),
            .I(N__19571));
    Sp12to4 I__2914 (
            .O(N__19603),
            .I(N__19558));
    LocalMux I__2913 (
            .O(N__19600),
            .I(N__19558));
    LocalMux I__2912 (
            .O(N__19597),
            .I(N__19558));
    LocalMux I__2911 (
            .O(N__19594),
            .I(N__19558));
    LocalMux I__2910 (
            .O(N__19591),
            .I(N__19558));
    LocalMux I__2909 (
            .O(N__19588),
            .I(N__19558));
    Span4Mux_v I__2908 (
            .O(N__19581),
            .I(N__19555));
    Span12Mux_h I__2907 (
            .O(N__19578),
            .I(N__19552));
    Span12Mux_s10_v I__2906 (
            .O(N__19571),
            .I(N__19547));
    Span12Mux_v I__2905 (
            .O(N__19558),
            .I(N__19547));
    Span4Mux_h I__2904 (
            .O(N__19555),
            .I(N__19544));
    Odrv12 I__2903 (
            .O(N__19552),
            .I(read_data_RNI7SFJ1_3));
    Odrv12 I__2902 (
            .O(N__19547),
            .I(read_data_RNI7SFJ1_3));
    Odrv4 I__2901 (
            .O(N__19544),
            .I(read_data_RNI7SFJ1_3));
    InMux I__2900 (
            .O(N__19537),
            .I(N__19534));
    LocalMux I__2899 (
            .O(N__19534),
            .I(N__19531));
    Span4Mux_h I__2898 (
            .O(N__19531),
            .I(N__19528));
    Span4Mux_v I__2897 (
            .O(N__19528),
            .I(N__19525));
    Odrv4 I__2896 (
            .O(N__19525),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_4 ));
    CascadeMux I__2895 (
            .O(N__19522),
            .I(N__19519));
    InMux I__2894 (
            .O(N__19519),
            .I(N__19513));
    CascadeMux I__2893 (
            .O(N__19518),
            .I(N__19510));
    CascadeMux I__2892 (
            .O(N__19517),
            .I(N__19505));
    CascadeMux I__2891 (
            .O(N__19516),
            .I(N__19502));
    LocalMux I__2890 (
            .O(N__19513),
            .I(N__19493));
    InMux I__2889 (
            .O(N__19510),
            .I(N__19490));
    CascadeMux I__2888 (
            .O(N__19509),
            .I(N__19487));
    CascadeMux I__2887 (
            .O(N__19508),
            .I(N__19482));
    InMux I__2886 (
            .O(N__19505),
            .I(N__19477));
    InMux I__2885 (
            .O(N__19502),
            .I(N__19474));
    CascadeMux I__2884 (
            .O(N__19501),
            .I(N__19471));
    CascadeMux I__2883 (
            .O(N__19500),
            .I(N__19468));
    CascadeMux I__2882 (
            .O(N__19499),
            .I(N__19465));
    CascadeMux I__2881 (
            .O(N__19498),
            .I(N__19462));
    CascadeMux I__2880 (
            .O(N__19497),
            .I(N__19459));
    CascadeMux I__2879 (
            .O(N__19496),
            .I(N__19456));
    Span4Mux_v I__2878 (
            .O(N__19493),
            .I(N__19451));
    LocalMux I__2877 (
            .O(N__19490),
            .I(N__19451));
    InMux I__2876 (
            .O(N__19487),
            .I(N__19448));
    CascadeMux I__2875 (
            .O(N__19486),
            .I(N__19445));
    CascadeMux I__2874 (
            .O(N__19485),
            .I(N__19442));
    InMux I__2873 (
            .O(N__19482),
            .I(N__19439));
    CascadeMux I__2872 (
            .O(N__19481),
            .I(N__19436));
    CascadeMux I__2871 (
            .O(N__19480),
            .I(N__19433));
    LocalMux I__2870 (
            .O(N__19477),
            .I(N__19430));
    LocalMux I__2869 (
            .O(N__19474),
            .I(N__19427));
    InMux I__2868 (
            .O(N__19471),
            .I(N__19424));
    InMux I__2867 (
            .O(N__19468),
            .I(N__19421));
    InMux I__2866 (
            .O(N__19465),
            .I(N__19418));
    InMux I__2865 (
            .O(N__19462),
            .I(N__19415));
    InMux I__2864 (
            .O(N__19459),
            .I(N__19412));
    InMux I__2863 (
            .O(N__19456),
            .I(N__19409));
    Span4Mux_v I__2862 (
            .O(N__19451),
            .I(N__19404));
    LocalMux I__2861 (
            .O(N__19448),
            .I(N__19404));
    InMux I__2860 (
            .O(N__19445),
            .I(N__19401));
    InMux I__2859 (
            .O(N__19442),
            .I(N__19398));
    LocalMux I__2858 (
            .O(N__19439),
            .I(N__19395));
    InMux I__2857 (
            .O(N__19436),
            .I(N__19392));
    InMux I__2856 (
            .O(N__19433),
            .I(N__19389));
    Span12Mux_s4_v I__2855 (
            .O(N__19430),
            .I(N__19384));
    Span12Mux_s7_h I__2854 (
            .O(N__19427),
            .I(N__19384));
    LocalMux I__2853 (
            .O(N__19424),
            .I(N__19377));
    LocalMux I__2852 (
            .O(N__19421),
            .I(N__19377));
    LocalMux I__2851 (
            .O(N__19418),
            .I(N__19377));
    LocalMux I__2850 (
            .O(N__19415),
            .I(N__19374));
    LocalMux I__2849 (
            .O(N__19412),
            .I(N__19363));
    LocalMux I__2848 (
            .O(N__19409),
            .I(N__19363));
    Sp12to4 I__2847 (
            .O(N__19404),
            .I(N__19363));
    LocalMux I__2846 (
            .O(N__19401),
            .I(N__19363));
    LocalMux I__2845 (
            .O(N__19398),
            .I(N__19363));
    Span4Mux_s3_v I__2844 (
            .O(N__19395),
            .I(N__19358));
    LocalMux I__2843 (
            .O(N__19392),
            .I(N__19358));
    LocalMux I__2842 (
            .O(N__19389),
            .I(N__19355));
    Span12Mux_h I__2841 (
            .O(N__19384),
            .I(N__19352));
    Span12Mux_v I__2840 (
            .O(N__19377),
            .I(N__19345));
    Sp12to4 I__2839 (
            .O(N__19374),
            .I(N__19345));
    Span12Mux_v I__2838 (
            .O(N__19363),
            .I(N__19345));
    Span4Mux_v I__2837 (
            .O(N__19358),
            .I(N__19340));
    Span4Mux_v I__2836 (
            .O(N__19355),
            .I(N__19340));
    Span12Mux_v I__2835 (
            .O(N__19352),
            .I(N__19335));
    Span12Mux_h I__2834 (
            .O(N__19345),
            .I(N__19335));
    Span4Mux_h I__2833 (
            .O(N__19340),
            .I(N__19332));
    Odrv12 I__2832 (
            .O(N__19335),
            .I(read_data_RNI9TFJ1_4));
    Odrv4 I__2831 (
            .O(N__19332),
            .I(read_data_RNI9TFJ1_4));
    InMux I__2830 (
            .O(N__19327),
            .I(N__19324));
    LocalMux I__2829 (
            .O(N__19324),
            .I(N__19321));
    Span4Mux_v I__2828 (
            .O(N__19321),
            .I(N__19318));
    Odrv4 I__2827 (
            .O(N__19318),
            .I(\this_vga_signals.M_pcounter_q_0Z0Z_1 ));
    InMux I__2826 (
            .O(N__19315),
            .I(N__19312));
    LocalMux I__2825 (
            .O(N__19312),
            .I(N__19309));
    Span4Mux_v I__2824 (
            .O(N__19309),
            .I(N__19306));
    Odrv4 I__2823 (
            .O(N__19306),
            .I(M_this_data_tmp_qZ0Z_11));
    InMux I__2822 (
            .O(N__19303),
            .I(N__19300));
    LocalMux I__2821 (
            .O(N__19300),
            .I(N__19297));
    Odrv12 I__2820 (
            .O(N__19297),
            .I(M_this_oam_ram_write_data_11));
    InMux I__2819 (
            .O(N__19294),
            .I(N__19291));
    LocalMux I__2818 (
            .O(N__19291),
            .I(N__19288));
    Odrv12 I__2817 (
            .O(N__19288),
            .I(M_this_oam_ram_write_data_12));
    InMux I__2816 (
            .O(N__19285),
            .I(N__19282));
    LocalMux I__2815 (
            .O(N__19282),
            .I(N__19279));
    Odrv12 I__2814 (
            .O(N__19279),
            .I(M_this_oam_ram_write_data_13));
    InMux I__2813 (
            .O(N__19276),
            .I(N__19273));
    LocalMux I__2812 (
            .O(N__19273),
            .I(N__19270));
    Odrv12 I__2811 (
            .O(N__19270),
            .I(M_this_oam_ram_write_data_14));
    InMux I__2810 (
            .O(N__19267),
            .I(N__19264));
    LocalMux I__2809 (
            .O(N__19264),
            .I(N__19260));
    InMux I__2808 (
            .O(N__19263),
            .I(N__19257));
    Span4Mux_v I__2807 (
            .O(N__19260),
            .I(N__19251));
    LocalMux I__2806 (
            .O(N__19257),
            .I(N__19251));
    InMux I__2805 (
            .O(N__19256),
            .I(N__19248));
    Span4Mux_v I__2804 (
            .O(N__19251),
            .I(N__19245));
    LocalMux I__2803 (
            .O(N__19248),
            .I(this_pixel_clk_M_counter_q_0));
    Odrv4 I__2802 (
            .O(N__19245),
            .I(this_pixel_clk_M_counter_q_0));
    InMux I__2801 (
            .O(N__19240),
            .I(N__19236));
    InMux I__2800 (
            .O(N__19239),
            .I(N__19233));
    LocalMux I__2799 (
            .O(N__19236),
            .I(N__19230));
    LocalMux I__2798 (
            .O(N__19233),
            .I(this_pixel_clk_M_counter_q_i_1));
    Odrv12 I__2797 (
            .O(N__19230),
            .I(this_pixel_clk_M_counter_q_i_1));
    InMux I__2796 (
            .O(N__19225),
            .I(N__19217));
    CascadeMux I__2795 (
            .O(N__19224),
            .I(N__19212));
    InMux I__2794 (
            .O(N__19223),
            .I(N__19206));
    InMux I__2793 (
            .O(N__19222),
            .I(N__19201));
    InMux I__2792 (
            .O(N__19221),
            .I(N__19201));
    InMux I__2791 (
            .O(N__19220),
            .I(N__19198));
    LocalMux I__2790 (
            .O(N__19217),
            .I(N__19195));
    InMux I__2789 (
            .O(N__19216),
            .I(N__19192));
    InMux I__2788 (
            .O(N__19215),
            .I(N__19189));
    InMux I__2787 (
            .O(N__19212),
            .I(N__19186));
    InMux I__2786 (
            .O(N__19211),
            .I(N__19183));
    InMux I__2785 (
            .O(N__19210),
            .I(N__19178));
    InMux I__2784 (
            .O(N__19209),
            .I(N__19178));
    LocalMux I__2783 (
            .O(N__19206),
            .I(N__19171));
    LocalMux I__2782 (
            .O(N__19201),
            .I(N__19171));
    LocalMux I__2781 (
            .O(N__19198),
            .I(N__19171));
    Span4Mux_h I__2780 (
            .O(N__19195),
            .I(N__19164));
    LocalMux I__2779 (
            .O(N__19192),
            .I(N__19164));
    LocalMux I__2778 (
            .O(N__19189),
            .I(N__19164));
    LocalMux I__2777 (
            .O(N__19186),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2776 (
            .O(N__19183),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2775 (
            .O(N__19178),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__2774 (
            .O(N__19171),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__2773 (
            .O(N__19164),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__2772 (
            .O(N__19153),
            .I(N__19146));
    InMux I__2771 (
            .O(N__19152),
            .I(N__19143));
    InMux I__2770 (
            .O(N__19151),
            .I(N__19138));
    InMux I__2769 (
            .O(N__19150),
            .I(N__19138));
    InMux I__2768 (
            .O(N__19149),
            .I(N__19135));
    LocalMux I__2767 (
            .O(N__19146),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ));
    LocalMux I__2766 (
            .O(N__19143),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ));
    LocalMux I__2765 (
            .O(N__19138),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ));
    LocalMux I__2764 (
            .O(N__19135),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ));
    InMux I__2763 (
            .O(N__19126),
            .I(N__19115));
    CascadeMux I__2762 (
            .O(N__19125),
            .I(N__19112));
    CascadeMux I__2761 (
            .O(N__19124),
            .I(N__19109));
    InMux I__2760 (
            .O(N__19123),
            .I(N__19101));
    InMux I__2759 (
            .O(N__19122),
            .I(N__19101));
    InMux I__2758 (
            .O(N__19121),
            .I(N__19101));
    InMux I__2757 (
            .O(N__19120),
            .I(N__19098));
    InMux I__2756 (
            .O(N__19119),
            .I(N__19095));
    InMux I__2755 (
            .O(N__19118),
            .I(N__19092));
    LocalMux I__2754 (
            .O(N__19115),
            .I(N__19089));
    InMux I__2753 (
            .O(N__19112),
            .I(N__19086));
    InMux I__2752 (
            .O(N__19109),
            .I(N__19083));
    InMux I__2751 (
            .O(N__19108),
            .I(N__19080));
    LocalMux I__2750 (
            .O(N__19101),
            .I(N__19073));
    LocalMux I__2749 (
            .O(N__19098),
            .I(N__19073));
    LocalMux I__2748 (
            .O(N__19095),
            .I(N__19073));
    LocalMux I__2747 (
            .O(N__19092),
            .I(N__19067));
    Span4Mux_v I__2746 (
            .O(N__19089),
            .I(N__19067));
    LocalMux I__2745 (
            .O(N__19086),
            .I(N__19064));
    LocalMux I__2744 (
            .O(N__19083),
            .I(N__19059));
    LocalMux I__2743 (
            .O(N__19080),
            .I(N__19059));
    Span4Mux_h I__2742 (
            .O(N__19073),
            .I(N__19056));
    InMux I__2741 (
            .O(N__19072),
            .I(N__19053));
    Odrv4 I__2740 (
            .O(N__19067),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv12 I__2739 (
            .O(N__19064),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__2738 (
            .O(N__19059),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__2737 (
            .O(N__19056),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__2736 (
            .O(N__19053),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__2735 (
            .O(N__19042),
            .I(N__19038));
    InMux I__2734 (
            .O(N__19041),
            .I(N__19035));
    LocalMux I__2733 (
            .O(N__19038),
            .I(N__19031));
    LocalMux I__2732 (
            .O(N__19035),
            .I(N__19024));
    InMux I__2731 (
            .O(N__19034),
            .I(N__19021));
    Span4Mux_h I__2730 (
            .O(N__19031),
            .I(N__19018));
    InMux I__2729 (
            .O(N__19030),
            .I(N__19015));
    InMux I__2728 (
            .O(N__19029),
            .I(N__19008));
    InMux I__2727 (
            .O(N__19028),
            .I(N__19008));
    InMux I__2726 (
            .O(N__19027),
            .I(N__19008));
    Odrv4 I__2725 (
            .O(N__19024),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_3 ));
    LocalMux I__2724 (
            .O(N__19021),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_3 ));
    Odrv4 I__2723 (
            .O(N__19018),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_3 ));
    LocalMux I__2722 (
            .O(N__19015),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_3 ));
    LocalMux I__2721 (
            .O(N__19008),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_3 ));
    CascadeMux I__2720 (
            .O(N__18997),
            .I(N__18993));
    CascadeMux I__2719 (
            .O(N__18996),
            .I(N__18990));
    InMux I__2718 (
            .O(N__18993),
            .I(N__18985));
    InMux I__2717 (
            .O(N__18990),
            .I(N__18985));
    LocalMux I__2716 (
            .O(N__18985),
            .I(N__18982));
    Odrv4 I__2715 (
            .O(N__18982),
            .I(\this_vga_signals.M_hcounter_q_RNII1437Z0Z_3 ));
    InMux I__2714 (
            .O(N__18979),
            .I(N__18976));
    LocalMux I__2713 (
            .O(N__18976),
            .I(N__18973));
    Span4Mux_h I__2712 (
            .O(N__18973),
            .I(N__18970));
    Span4Mux_h I__2711 (
            .O(N__18970),
            .I(N__18967));
    Odrv4 I__2710 (
            .O(N__18967),
            .I(M_this_oam_ram_read_data_30));
    InMux I__2709 (
            .O(N__18964),
            .I(N__18961));
    LocalMux I__2708 (
            .O(N__18961),
            .I(N__18958));
    Span4Mux_h I__2707 (
            .O(N__18958),
            .I(N__18955));
    Span4Mux_h I__2706 (
            .O(N__18955),
            .I(N__18952));
    Odrv4 I__2705 (
            .O(N__18952),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_30 ));
    InMux I__2704 (
            .O(N__18949),
            .I(N__18946));
    LocalMux I__2703 (
            .O(N__18946),
            .I(N__18943));
    Span4Mux_h I__2702 (
            .O(N__18943),
            .I(N__18940));
    Span4Mux_h I__2701 (
            .O(N__18940),
            .I(N__18937));
    Odrv4 I__2700 (
            .O(N__18937),
            .I(\this_ppu.oam_cache.mem_3 ));
    InMux I__2699 (
            .O(N__18934),
            .I(N__18931));
    LocalMux I__2698 (
            .O(N__18931),
            .I(N__18928));
    Span4Mux_v I__2697 (
            .O(N__18928),
            .I(N__18925));
    Odrv4 I__2696 (
            .O(N__18925),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_1 ));
    CascadeMux I__2695 (
            .O(N__18922),
            .I(N__18918));
    CascadeMux I__2694 (
            .O(N__18921),
            .I(N__18913));
    InMux I__2693 (
            .O(N__18918),
            .I(N__18910));
    CascadeMux I__2692 (
            .O(N__18917),
            .I(N__18907));
    CascadeMux I__2691 (
            .O(N__18916),
            .I(N__18900));
    InMux I__2690 (
            .O(N__18913),
            .I(N__18891));
    LocalMux I__2689 (
            .O(N__18910),
            .I(N__18888));
    InMux I__2688 (
            .O(N__18907),
            .I(N__18885));
    CascadeMux I__2687 (
            .O(N__18906),
            .I(N__18882));
    CascadeMux I__2686 (
            .O(N__18905),
            .I(N__18879));
    CascadeMux I__2685 (
            .O(N__18904),
            .I(N__18876));
    CascadeMux I__2684 (
            .O(N__18903),
            .I(N__18873));
    InMux I__2683 (
            .O(N__18900),
            .I(N__18870));
    CascadeMux I__2682 (
            .O(N__18899),
            .I(N__18867));
    CascadeMux I__2681 (
            .O(N__18898),
            .I(N__18864));
    CascadeMux I__2680 (
            .O(N__18897),
            .I(N__18861));
    CascadeMux I__2679 (
            .O(N__18896),
            .I(N__18858));
    CascadeMux I__2678 (
            .O(N__18895),
            .I(N__18855));
    CascadeMux I__2677 (
            .O(N__18894),
            .I(N__18851));
    LocalMux I__2676 (
            .O(N__18891),
            .I(N__18847));
    Span4Mux_v I__2675 (
            .O(N__18888),
            .I(N__18844));
    LocalMux I__2674 (
            .O(N__18885),
            .I(N__18841));
    InMux I__2673 (
            .O(N__18882),
            .I(N__18838));
    InMux I__2672 (
            .O(N__18879),
            .I(N__18835));
    InMux I__2671 (
            .O(N__18876),
            .I(N__18832));
    InMux I__2670 (
            .O(N__18873),
            .I(N__18829));
    LocalMux I__2669 (
            .O(N__18870),
            .I(N__18826));
    InMux I__2668 (
            .O(N__18867),
            .I(N__18823));
    InMux I__2667 (
            .O(N__18864),
            .I(N__18820));
    InMux I__2666 (
            .O(N__18861),
            .I(N__18817));
    InMux I__2665 (
            .O(N__18858),
            .I(N__18814));
    InMux I__2664 (
            .O(N__18855),
            .I(N__18811));
    CascadeMux I__2663 (
            .O(N__18854),
            .I(N__18808));
    InMux I__2662 (
            .O(N__18851),
            .I(N__18805));
    CascadeMux I__2661 (
            .O(N__18850),
            .I(N__18802));
    Span12Mux_s6_v I__2660 (
            .O(N__18847),
            .I(N__18795));
    Sp12to4 I__2659 (
            .O(N__18844),
            .I(N__18795));
    Span12Mux_s7_h I__2658 (
            .O(N__18841),
            .I(N__18795));
    LocalMux I__2657 (
            .O(N__18838),
            .I(N__18786));
    LocalMux I__2656 (
            .O(N__18835),
            .I(N__18786));
    LocalMux I__2655 (
            .O(N__18832),
            .I(N__18786));
    LocalMux I__2654 (
            .O(N__18829),
            .I(N__18786));
    Span4Mux_v I__2653 (
            .O(N__18826),
            .I(N__18783));
    LocalMux I__2652 (
            .O(N__18823),
            .I(N__18780));
    LocalMux I__2651 (
            .O(N__18820),
            .I(N__18771));
    LocalMux I__2650 (
            .O(N__18817),
            .I(N__18771));
    LocalMux I__2649 (
            .O(N__18814),
            .I(N__18771));
    LocalMux I__2648 (
            .O(N__18811),
            .I(N__18771));
    InMux I__2647 (
            .O(N__18808),
            .I(N__18768));
    LocalMux I__2646 (
            .O(N__18805),
            .I(N__18765));
    InMux I__2645 (
            .O(N__18802),
            .I(N__18762));
    Span12Mux_h I__2644 (
            .O(N__18795),
            .I(N__18759));
    Span12Mux_v I__2643 (
            .O(N__18786),
            .I(N__18750));
    Sp12to4 I__2642 (
            .O(N__18783),
            .I(N__18750));
    Sp12to4 I__2641 (
            .O(N__18780),
            .I(N__18750));
    Span12Mux_v I__2640 (
            .O(N__18771),
            .I(N__18750));
    LocalMux I__2639 (
            .O(N__18768),
            .I(N__18743));
    Sp12to4 I__2638 (
            .O(N__18765),
            .I(N__18743));
    LocalMux I__2637 (
            .O(N__18762),
            .I(N__18743));
    Span12Mux_v I__2636 (
            .O(N__18759),
            .I(N__18738));
    Span12Mux_h I__2635 (
            .O(N__18750),
            .I(N__18738));
    Span12Mux_s10_v I__2634 (
            .O(N__18743),
            .I(N__18735));
    Odrv12 I__2633 (
            .O(N__18738),
            .I(read_data_RNI5QFJ1_1));
    Odrv12 I__2632 (
            .O(N__18735),
            .I(read_data_RNI5QFJ1_1));
    InMux I__2631 (
            .O(N__18730),
            .I(N__18726));
    InMux I__2630 (
            .O(N__18729),
            .I(N__18723));
    LocalMux I__2629 (
            .O(N__18726),
            .I(N__18718));
    LocalMux I__2628 (
            .O(N__18723),
            .I(N__18718));
    Odrv4 I__2627 (
            .O(N__18718),
            .I(\this_ppu.N_1196_1 ));
    InMux I__2626 (
            .O(N__18715),
            .I(N__18708));
    InMux I__2625 (
            .O(N__18714),
            .I(N__18708));
    CascadeMux I__2624 (
            .O(N__18713),
            .I(N__18705));
    LocalMux I__2623 (
            .O(N__18708),
            .I(N__18702));
    InMux I__2622 (
            .O(N__18705),
            .I(N__18699));
    Span4Mux_h I__2621 (
            .O(N__18702),
            .I(N__18696));
    LocalMux I__2620 (
            .O(N__18699),
            .I(\this_ppu.M_oam_curr_qZ0Z_6 ));
    Odrv4 I__2619 (
            .O(N__18696),
            .I(\this_ppu.M_oam_curr_qZ0Z_6 ));
    InMux I__2618 (
            .O(N__18691),
            .I(N__18688));
    LocalMux I__2617 (
            .O(N__18688),
            .I(N__18685));
    Odrv4 I__2616 (
            .O(N__18685),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_13 ));
    SRMux I__2615 (
            .O(N__18682),
            .I(N__18678));
    SRMux I__2614 (
            .O(N__18681),
            .I(N__18675));
    LocalMux I__2613 (
            .O(N__18678),
            .I(N__18671));
    LocalMux I__2612 (
            .O(N__18675),
            .I(N__18668));
    SRMux I__2611 (
            .O(N__18674),
            .I(N__18665));
    Span4Mux_v I__2610 (
            .O(N__18671),
            .I(N__18658));
    Span4Mux_h I__2609 (
            .O(N__18668),
            .I(N__18658));
    LocalMux I__2608 (
            .O(N__18665),
            .I(N__18658));
    Sp12to4 I__2607 (
            .O(N__18658),
            .I(N__18655));
    Odrv12 I__2606 (
            .O(N__18655),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9 ));
    CascadeMux I__2605 (
            .O(N__18652),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9_cascade_ ));
    CEMux I__2604 (
            .O(N__18649),
            .I(N__18646));
    LocalMux I__2603 (
            .O(N__18646),
            .I(\this_vga_signals.N_1307_1 ));
    InMux I__2602 (
            .O(N__18643),
            .I(N__18640));
    LocalMux I__2601 (
            .O(N__18640),
            .I(N__18637));
    Span4Mux_h I__2600 (
            .O(N__18637),
            .I(N__18634));
    Span4Mux_h I__2599 (
            .O(N__18634),
            .I(N__18631));
    Odrv4 I__2598 (
            .O(N__18631),
            .I(\this_ppu.oam_cache.mem_8 ));
    InMux I__2597 (
            .O(N__18628),
            .I(N__18625));
    LocalMux I__2596 (
            .O(N__18625),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_11 ));
    CascadeMux I__2595 (
            .O(N__18622),
            .I(N__18615));
    CascadeMux I__2594 (
            .O(N__18621),
            .I(N__18611));
    CascadeMux I__2593 (
            .O(N__18620),
            .I(N__18607));
    CascadeMux I__2592 (
            .O(N__18619),
            .I(N__18604));
    InMux I__2591 (
            .O(N__18618),
            .I(N__18600));
    InMux I__2590 (
            .O(N__18615),
            .I(N__18595));
    InMux I__2589 (
            .O(N__18614),
            .I(N__18595));
    InMux I__2588 (
            .O(N__18611),
            .I(N__18589));
    InMux I__2587 (
            .O(N__18610),
            .I(N__18589));
    InMux I__2586 (
            .O(N__18607),
            .I(N__18586));
    InMux I__2585 (
            .O(N__18604),
            .I(N__18583));
    InMux I__2584 (
            .O(N__18603),
            .I(N__18580));
    LocalMux I__2583 (
            .O(N__18600),
            .I(N__18577));
    LocalMux I__2582 (
            .O(N__18595),
            .I(N__18574));
    InMux I__2581 (
            .O(N__18594),
            .I(N__18571));
    LocalMux I__2580 (
            .O(N__18589),
            .I(N__18568));
    LocalMux I__2579 (
            .O(N__18586),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2578 (
            .O(N__18583),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2577 (
            .O(N__18580),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__2576 (
            .O(N__18577),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv12 I__2575 (
            .O(N__18574),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2574 (
            .O(N__18571),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__2573 (
            .O(N__18568),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    InMux I__2572 (
            .O(N__18553),
            .I(N__18550));
    LocalMux I__2571 (
            .O(N__18550),
            .I(N__18546));
    InMux I__2570 (
            .O(N__18549),
            .I(N__18543));
    Odrv4 I__2569 (
            .O(N__18546),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1_0 ));
    LocalMux I__2568 (
            .O(N__18543),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1_0 ));
    CascadeMux I__2567 (
            .O(N__18538),
            .I(\this_vga_signals.N_2_0_cascade_ ));
    InMux I__2566 (
            .O(N__18535),
            .I(N__18532));
    LocalMux I__2565 (
            .O(N__18532),
            .I(N__18529));
    Odrv4 I__2564 (
            .O(N__18529),
            .I(\this_vga_ramdac.m19 ));
    InMux I__2563 (
            .O(N__18526),
            .I(N__18522));
    CascadeMux I__2562 (
            .O(N__18525),
            .I(N__18519));
    LocalMux I__2561 (
            .O(N__18522),
            .I(N__18516));
    InMux I__2560 (
            .O(N__18519),
            .I(N__18513));
    Odrv12 I__2559 (
            .O(N__18516),
            .I(\this_vga_ramdac.N_3860_reto ));
    LocalMux I__2558 (
            .O(N__18513),
            .I(\this_vga_ramdac.N_3860_reto ));
    InMux I__2557 (
            .O(N__18508),
            .I(N__18505));
    LocalMux I__2556 (
            .O(N__18505),
            .I(N__18502));
    Span12Mux_h I__2555 (
            .O(N__18502),
            .I(N__18499));
    Odrv12 I__2554 (
            .O(N__18499),
            .I(\this_ppu.oam_cache.mem_14 ));
    CascadeMux I__2553 (
            .O(N__18496),
            .I(\this_ppu.m35_i_0_a3_0_cascade_ ));
    InMux I__2552 (
            .O(N__18493),
            .I(N__18490));
    LocalMux I__2551 (
            .O(N__18490),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_9 ));
    InMux I__2550 (
            .O(N__18487),
            .I(N__18484));
    LocalMux I__2549 (
            .O(N__18484),
            .I(N__18481));
    Span4Mux_v I__2548 (
            .O(N__18481),
            .I(N__18478));
    Span4Mux_h I__2547 (
            .O(N__18478),
            .I(N__18475));
    Odrv4 I__2546 (
            .O(N__18475),
            .I(\this_ppu.oam_cache.mem_11 ));
    InMux I__2545 (
            .O(N__18472),
            .I(N__18469));
    LocalMux I__2544 (
            .O(N__18469),
            .I(N__18466));
    Span4Mux_h I__2543 (
            .O(N__18466),
            .I(N__18463));
    Odrv4 I__2542 (
            .O(N__18463),
            .I(\this_ppu.oam_cache.mem_1 ));
    InMux I__2541 (
            .O(N__18460),
            .I(N__18457));
    LocalMux I__2540 (
            .O(N__18457),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_14 ));
    InMux I__2539 (
            .O(N__18454),
            .I(N__18451));
    LocalMux I__2538 (
            .O(N__18451),
            .I(\this_vga_ramdac.N_24_mux ));
    InMux I__2537 (
            .O(N__18448),
            .I(N__18439));
    InMux I__2536 (
            .O(N__18447),
            .I(N__18439));
    InMux I__2535 (
            .O(N__18446),
            .I(N__18439));
    LocalMux I__2534 (
            .O(N__18439),
            .I(N__18434));
    InMux I__2533 (
            .O(N__18438),
            .I(N__18429));
    InMux I__2532 (
            .O(N__18437),
            .I(N__18429));
    Span4Mux_v I__2531 (
            .O(N__18434),
            .I(N__18423));
    LocalMux I__2530 (
            .O(N__18429),
            .I(N__18423));
    InMux I__2529 (
            .O(N__18428),
            .I(N__18420));
    Span4Mux_h I__2528 (
            .O(N__18423),
            .I(N__18415));
    LocalMux I__2527 (
            .O(N__18420),
            .I(N__18415));
    Span4Mux_v I__2526 (
            .O(N__18415),
            .I(N__18412));
    Odrv4 I__2525 (
            .O(N__18412),
            .I(M_this_vram_read_data_0));
    CascadeMux I__2524 (
            .O(N__18409),
            .I(N__18405));
    InMux I__2523 (
            .O(N__18408),
            .I(N__18399));
    InMux I__2522 (
            .O(N__18405),
            .I(N__18399));
    CascadeMux I__2521 (
            .O(N__18404),
            .I(N__18395));
    LocalMux I__2520 (
            .O(N__18399),
            .I(N__18391));
    InMux I__2519 (
            .O(N__18398),
            .I(N__18386));
    InMux I__2518 (
            .O(N__18395),
            .I(N__18386));
    CascadeMux I__2517 (
            .O(N__18394),
            .I(N__18383));
    Span4Mux_h I__2516 (
            .O(N__18391),
            .I(N__18380));
    LocalMux I__2515 (
            .O(N__18386),
            .I(N__18377));
    InMux I__2514 (
            .O(N__18383),
            .I(N__18374));
    Span4Mux_h I__2513 (
            .O(N__18380),
            .I(N__18371));
    Span4Mux_v I__2512 (
            .O(N__18377),
            .I(N__18366));
    LocalMux I__2511 (
            .O(N__18374),
            .I(N__18366));
    Span4Mux_v I__2510 (
            .O(N__18371),
            .I(N__18363));
    Span4Mux_h I__2509 (
            .O(N__18366),
            .I(N__18360));
    Odrv4 I__2508 (
            .O(N__18363),
            .I(M_this_vram_read_data_2));
    Odrv4 I__2507 (
            .O(N__18360),
            .I(M_this_vram_read_data_2));
    CascadeMux I__2506 (
            .O(N__18355),
            .I(N__18350));
    InMux I__2505 (
            .O(N__18354),
            .I(N__18343));
    InMux I__2504 (
            .O(N__18353),
            .I(N__18343));
    InMux I__2503 (
            .O(N__18350),
            .I(N__18335));
    InMux I__2502 (
            .O(N__18349),
            .I(N__18335));
    InMux I__2501 (
            .O(N__18348),
            .I(N__18335));
    LocalMux I__2500 (
            .O(N__18343),
            .I(N__18332));
    InMux I__2499 (
            .O(N__18342),
            .I(N__18329));
    LocalMux I__2498 (
            .O(N__18335),
            .I(N__18326));
    Span4Mux_h I__2497 (
            .O(N__18332),
            .I(N__18323));
    LocalMux I__2496 (
            .O(N__18329),
            .I(N__18318));
    Span4Mux_v I__2495 (
            .O(N__18326),
            .I(N__18318));
    Span4Mux_v I__2494 (
            .O(N__18323),
            .I(N__18315));
    Span4Mux_h I__2493 (
            .O(N__18318),
            .I(N__18312));
    Odrv4 I__2492 (
            .O(N__18315),
            .I(M_this_vram_read_data_3));
    Odrv4 I__2491 (
            .O(N__18312),
            .I(M_this_vram_read_data_3));
    CascadeMux I__2490 (
            .O(N__18307),
            .I(N__18304));
    InMux I__2489 (
            .O(N__18304),
            .I(N__18295));
    InMux I__2488 (
            .O(N__18303),
            .I(N__18295));
    InMux I__2487 (
            .O(N__18302),
            .I(N__18287));
    InMux I__2486 (
            .O(N__18301),
            .I(N__18287));
    InMux I__2485 (
            .O(N__18300),
            .I(N__18287));
    LocalMux I__2484 (
            .O(N__18295),
            .I(N__18284));
    InMux I__2483 (
            .O(N__18294),
            .I(N__18281));
    LocalMux I__2482 (
            .O(N__18287),
            .I(N__18278));
    Span4Mux_h I__2481 (
            .O(N__18284),
            .I(N__18275));
    LocalMux I__2480 (
            .O(N__18281),
            .I(N__18272));
    Span12Mux_h I__2479 (
            .O(N__18278),
            .I(N__18269));
    Span4Mux_v I__2478 (
            .O(N__18275),
            .I(N__18266));
    Span4Mux_v I__2477 (
            .O(N__18272),
            .I(N__18263));
    Odrv12 I__2476 (
            .O(N__18269),
            .I(M_this_vram_read_data_1));
    Odrv4 I__2475 (
            .O(N__18266),
            .I(M_this_vram_read_data_1));
    Odrv4 I__2474 (
            .O(N__18263),
            .I(M_this_vram_read_data_1));
    CascadeMux I__2473 (
            .O(N__18256),
            .I(\this_vga_ramdac.m6_cascade_ ));
    InMux I__2472 (
            .O(N__18253),
            .I(N__18250));
    LocalMux I__2471 (
            .O(N__18250),
            .I(N__18246));
    InMux I__2470 (
            .O(N__18249),
            .I(N__18243));
    Odrv4 I__2469 (
            .O(N__18246),
            .I(\this_vga_ramdac.N_3857_reto ));
    LocalMux I__2468 (
            .O(N__18243),
            .I(\this_vga_ramdac.N_3857_reto ));
    InMux I__2467 (
            .O(N__18238),
            .I(N__18235));
    LocalMux I__2466 (
            .O(N__18235),
            .I(N__18232));
    Odrv12 I__2465 (
            .O(N__18232),
            .I(\this_ppu.oam_cache.mem_9 ));
    CascadeMux I__2464 (
            .O(N__18229),
            .I(\this_vga_signals.M_pcounter_q_ret_RNIB85CZ0Z3_cascade_ ));
    CascadeMux I__2463 (
            .O(N__18226),
            .I(\this_vga_signals.N_3_0_cascade_ ));
    InMux I__2462 (
            .O(N__18223),
            .I(N__18220));
    LocalMux I__2461 (
            .O(N__18220),
            .I(N__18217));
    Odrv4 I__2460 (
            .O(N__18217),
            .I(\this_vga_ramdac.m16 ));
    CascadeMux I__2459 (
            .O(N__18214),
            .I(M_pcounter_q_ret_1_RNIOILK7_cascade_));
    InMux I__2458 (
            .O(N__18211),
            .I(N__18208));
    LocalMux I__2457 (
            .O(N__18208),
            .I(N__18204));
    InMux I__2456 (
            .O(N__18207),
            .I(N__18201));
    Odrv4 I__2455 (
            .O(N__18204),
            .I(\this_vga_ramdac.N_3859_reto ));
    LocalMux I__2454 (
            .O(N__18201),
            .I(\this_vga_ramdac.N_3859_reto ));
    InMux I__2453 (
            .O(N__18196),
            .I(N__18193));
    LocalMux I__2452 (
            .O(N__18193),
            .I(\this_vga_signals.N_2_0 ));
    InMux I__2451 (
            .O(N__18190),
            .I(N__18187));
    LocalMux I__2450 (
            .O(N__18187),
            .I(N__18184));
    Span4Mux_h I__2449 (
            .O(N__18184),
            .I(N__18181));
    Odrv4 I__2448 (
            .O(N__18181),
            .I(M_this_oam_ram_write_data_1));
    InMux I__2447 (
            .O(N__18178),
            .I(N__18175));
    LocalMux I__2446 (
            .O(N__18175),
            .I(N__18172));
    Odrv12 I__2445 (
            .O(N__18172),
            .I(M_this_oam_ram_write_data_25));
    InMux I__2444 (
            .O(N__18169),
            .I(N__18166));
    LocalMux I__2443 (
            .O(N__18166),
            .I(M_this_data_tmp_qZ0Z_21));
    InMux I__2442 (
            .O(N__18163),
            .I(N__18160));
    LocalMux I__2441 (
            .O(N__18160),
            .I(N__18157));
    Odrv4 I__2440 (
            .O(N__18157),
            .I(M_this_data_tmp_qZ0Z_23));
    InMux I__2439 (
            .O(N__18154),
            .I(N__18151));
    LocalMux I__2438 (
            .O(N__18151),
            .I(M_this_data_tmp_qZ0Z_0));
    InMux I__2437 (
            .O(N__18148),
            .I(N__18144));
    CascadeMux I__2436 (
            .O(N__18147),
            .I(N__18141));
    LocalMux I__2435 (
            .O(N__18144),
            .I(N__18138));
    InMux I__2434 (
            .O(N__18141),
            .I(N__18135));
    Odrv12 I__2433 (
            .O(N__18138),
            .I(\this_vga_ramdac.N_3856_reto ));
    LocalMux I__2432 (
            .O(N__18135),
            .I(\this_vga_ramdac.N_3856_reto ));
    CascadeMux I__2431 (
            .O(N__18130),
            .I(\this_vga_ramdac.i2_mux_cascade_ ));
    InMux I__2430 (
            .O(N__18127),
            .I(N__18124));
    LocalMux I__2429 (
            .O(N__18124),
            .I(N__18121));
    Span4Mux_h I__2428 (
            .O(N__18121),
            .I(N__18117));
    InMux I__2427 (
            .O(N__18120),
            .I(N__18114));
    Odrv4 I__2426 (
            .O(N__18117),
            .I(\this_vga_ramdac.N_3858_reto ));
    LocalMux I__2425 (
            .O(N__18114),
            .I(\this_vga_ramdac.N_3858_reto ));
    InMux I__2424 (
            .O(N__18109),
            .I(N__18106));
    LocalMux I__2423 (
            .O(N__18106),
            .I(N__18101));
    InMux I__2422 (
            .O(N__18105),
            .I(N__18098));
    CascadeMux I__2421 (
            .O(N__18104),
            .I(N__18093));
    Span4Mux_v I__2420 (
            .O(N__18101),
            .I(N__18088));
    LocalMux I__2419 (
            .O(N__18098),
            .I(N__18085));
    InMux I__2418 (
            .O(N__18097),
            .I(N__18080));
    InMux I__2417 (
            .O(N__18096),
            .I(N__18080));
    InMux I__2416 (
            .O(N__18093),
            .I(N__18075));
    InMux I__2415 (
            .O(N__18092),
            .I(N__18075));
    InMux I__2414 (
            .O(N__18091),
            .I(N__18072));
    Odrv4 I__2413 (
            .O(N__18088),
            .I(N_852_0));
    Odrv4 I__2412 (
            .O(N__18085),
            .I(N_852_0));
    LocalMux I__2411 (
            .O(N__18080),
            .I(N_852_0));
    LocalMux I__2410 (
            .O(N__18075),
            .I(N_852_0));
    LocalMux I__2409 (
            .O(N__18072),
            .I(N_852_0));
    CascadeMux I__2408 (
            .O(N__18061),
            .I(N__18058));
    InMux I__2407 (
            .O(N__18058),
            .I(N__18054));
    InMux I__2406 (
            .O(N__18057),
            .I(N__18051));
    LocalMux I__2405 (
            .O(N__18054),
            .I(N__18048));
    LocalMux I__2404 (
            .O(N__18051),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    Odrv4 I__2403 (
            .O(N__18048),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    CascadeMux I__2402 (
            .O(N__18043),
            .I(N__18040));
    InMux I__2401 (
            .O(N__18040),
            .I(N__18037));
    LocalMux I__2400 (
            .O(N__18037),
            .I(N__18034));
    Span4Mux_h I__2399 (
            .O(N__18034),
            .I(N__18031));
    Odrv4 I__2398 (
            .O(N__18031),
            .I(M_this_vga_signals_address_5));
    InMux I__2397 (
            .O(N__18028),
            .I(N__18025));
    LocalMux I__2396 (
            .O(N__18025),
            .I(N__18022));
    Span4Mux_h I__2395 (
            .O(N__18022),
            .I(N__18019));
    Odrv4 I__2394 (
            .O(N__18019),
            .I(M_this_oam_ram_write_data_3));
    InMux I__2393 (
            .O(N__18016),
            .I(N__18013));
    LocalMux I__2392 (
            .O(N__18013),
            .I(M_this_data_tmp_qZ0Z_3));
    InMux I__2391 (
            .O(N__18010),
            .I(N__18007));
    LocalMux I__2390 (
            .O(N__18007),
            .I(N__18004));
    Span4Mux_v I__2389 (
            .O(N__18004),
            .I(N__18001));
    Odrv4 I__2388 (
            .O(N__18001),
            .I(M_this_oam_ram_write_data_4));
    InMux I__2387 (
            .O(N__17998),
            .I(N__17995));
    LocalMux I__2386 (
            .O(N__17995),
            .I(M_this_data_tmp_qZ0Z_4));
    InMux I__2385 (
            .O(N__17992),
            .I(N__17989));
    LocalMux I__2384 (
            .O(N__17989),
            .I(N__17986));
    Span4Mux_h I__2383 (
            .O(N__17986),
            .I(N__17983));
    Odrv4 I__2382 (
            .O(N__17983),
            .I(M_this_data_tmp_qZ0Z_5));
    InMux I__2381 (
            .O(N__17980),
            .I(N__17977));
    LocalMux I__2380 (
            .O(N__17977),
            .I(N__17974));
    Odrv12 I__2379 (
            .O(N__17974),
            .I(M_this_oam_ram_write_data_29));
    InMux I__2378 (
            .O(N__17971),
            .I(N__17968));
    LocalMux I__2377 (
            .O(N__17968),
            .I(N__17965));
    Span4Mux_h I__2376 (
            .O(N__17965),
            .I(N__17962));
    Odrv4 I__2375 (
            .O(N__17962),
            .I(M_this_oam_ram_write_data_21));
    CascadeMux I__2374 (
            .O(N__17959),
            .I(\this_vga_signals.mult1_un54_sum_c3_cascade_ ));
    CascadeMux I__2373 (
            .O(N__17956),
            .I(N__17953));
    InMux I__2372 (
            .O(N__17953),
            .I(N__17949));
    InMux I__2371 (
            .O(N__17952),
            .I(N__17946));
    LocalMux I__2370 (
            .O(N__17949),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_0 ));
    LocalMux I__2369 (
            .O(N__17946),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_0 ));
    InMux I__2368 (
            .O(N__17941),
            .I(N__17938));
    LocalMux I__2367 (
            .O(N__17938),
            .I(N__17934));
    InMux I__2366 (
            .O(N__17937),
            .I(N__17931));
    Span4Mux_v I__2365 (
            .O(N__17934),
            .I(N__17924));
    LocalMux I__2364 (
            .O(N__17931),
            .I(N__17924));
    InMux I__2363 (
            .O(N__17930),
            .I(N__17921));
    InMux I__2362 (
            .O(N__17929),
            .I(N__17917));
    Span4Mux_h I__2361 (
            .O(N__17924),
            .I(N__17909));
    LocalMux I__2360 (
            .O(N__17921),
            .I(N__17909));
    InMux I__2359 (
            .O(N__17920),
            .I(N__17906));
    LocalMux I__2358 (
            .O(N__17917),
            .I(N__17902));
    InMux I__2357 (
            .O(N__17916),
            .I(N__17899));
    InMux I__2356 (
            .O(N__17915),
            .I(N__17894));
    InMux I__2355 (
            .O(N__17914),
            .I(N__17894));
    Span4Mux_v I__2354 (
            .O(N__17909),
            .I(N__17889));
    LocalMux I__2353 (
            .O(N__17906),
            .I(N__17889));
    InMux I__2352 (
            .O(N__17905),
            .I(N__17886));
    Odrv4 I__2351 (
            .O(N__17902),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2350 (
            .O(N__17899),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2349 (
            .O(N__17894),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__2348 (
            .O(N__17889),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2347 (
            .O(N__17886),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__2346 (
            .O(N__17875),
            .I(N__17871));
    InMux I__2345 (
            .O(N__17874),
            .I(N__17867));
    LocalMux I__2344 (
            .O(N__17871),
            .I(N__17864));
    InMux I__2343 (
            .O(N__17870),
            .I(N__17861));
    LocalMux I__2342 (
            .O(N__17867),
            .I(N__17857));
    Span4Mux_h I__2341 (
            .O(N__17864),
            .I(N__17848));
    LocalMux I__2340 (
            .O(N__17861),
            .I(N__17848));
    InMux I__2339 (
            .O(N__17860),
            .I(N__17845));
    Span12Mux_s11_h I__2338 (
            .O(N__17857),
            .I(N__17841));
    InMux I__2337 (
            .O(N__17856),
            .I(N__17838));
    InMux I__2336 (
            .O(N__17855),
            .I(N__17835));
    InMux I__2335 (
            .O(N__17854),
            .I(N__17832));
    InMux I__2334 (
            .O(N__17853),
            .I(N__17829));
    Span4Mux_v I__2333 (
            .O(N__17848),
            .I(N__17824));
    LocalMux I__2332 (
            .O(N__17845),
            .I(N__17824));
    InMux I__2331 (
            .O(N__17844),
            .I(N__17821));
    Odrv12 I__2330 (
            .O(N__17841),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2329 (
            .O(N__17838),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2328 (
            .O(N__17835),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2327 (
            .O(N__17832),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2326 (
            .O(N__17829),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__2325 (
            .O(N__17824),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2324 (
            .O(N__17821),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    InMux I__2323 (
            .O(N__17806),
            .I(N__17802));
    CascadeMux I__2322 (
            .O(N__17805),
            .I(N__17799));
    LocalMux I__2321 (
            .O(N__17802),
            .I(N__17796));
    InMux I__2320 (
            .O(N__17799),
            .I(N__17793));
    Span4Mux_h I__2319 (
            .O(N__17796),
            .I(N__17788));
    LocalMux I__2318 (
            .O(N__17793),
            .I(N__17788));
    Span4Mux_h I__2317 (
            .O(N__17788),
            .I(N__17781));
    InMux I__2316 (
            .O(N__17787),
            .I(N__17778));
    CascadeMux I__2315 (
            .O(N__17786),
            .I(N__17775));
    InMux I__2314 (
            .O(N__17785),
            .I(N__17770));
    CascadeMux I__2313 (
            .O(N__17784),
            .I(N__17766));
    Span4Mux_v I__2312 (
            .O(N__17781),
            .I(N__17761));
    LocalMux I__2311 (
            .O(N__17778),
            .I(N__17761));
    InMux I__2310 (
            .O(N__17775),
            .I(N__17758));
    InMux I__2309 (
            .O(N__17774),
            .I(N__17755));
    InMux I__2308 (
            .O(N__17773),
            .I(N__17752));
    LocalMux I__2307 (
            .O(N__17770),
            .I(N__17749));
    InMux I__2306 (
            .O(N__17769),
            .I(N__17744));
    InMux I__2305 (
            .O(N__17766),
            .I(N__17744));
    Span4Mux_v I__2304 (
            .O(N__17761),
            .I(N__17739));
    LocalMux I__2303 (
            .O(N__17758),
            .I(N__17739));
    LocalMux I__2302 (
            .O(N__17755),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2301 (
            .O(N__17752),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__2300 (
            .O(N__17749),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2299 (
            .O(N__17744),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__2298 (
            .O(N__17739),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    InMux I__2297 (
            .O(N__17728),
            .I(N__17724));
    InMux I__2296 (
            .O(N__17727),
            .I(N__17721));
    LocalMux I__2295 (
            .O(N__17724),
            .I(\this_vga_signals.N_968 ));
    LocalMux I__2294 (
            .O(N__17721),
            .I(\this_vga_signals.N_968 ));
    CascadeMux I__2293 (
            .O(N__17716),
            .I(N__17713));
    InMux I__2292 (
            .O(N__17713),
            .I(N__17703));
    InMux I__2291 (
            .O(N__17712),
            .I(N__17694));
    InMux I__2290 (
            .O(N__17711),
            .I(N__17694));
    InMux I__2289 (
            .O(N__17710),
            .I(N__17694));
    InMux I__2288 (
            .O(N__17709),
            .I(N__17689));
    InMux I__2287 (
            .O(N__17708),
            .I(N__17689));
    InMux I__2286 (
            .O(N__17707),
            .I(N__17686));
    InMux I__2285 (
            .O(N__17706),
            .I(N__17683));
    LocalMux I__2284 (
            .O(N__17703),
            .I(N__17680));
    InMux I__2283 (
            .O(N__17702),
            .I(N__17675));
    InMux I__2282 (
            .O(N__17701),
            .I(N__17675));
    LocalMux I__2281 (
            .O(N__17694),
            .I(N__17670));
    LocalMux I__2280 (
            .O(N__17689),
            .I(N__17670));
    LocalMux I__2279 (
            .O(N__17686),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2278 (
            .O(N__17683),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__2277 (
            .O(N__17680),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2276 (
            .O(N__17675),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__2275 (
            .O(N__17670),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    CascadeMux I__2274 (
            .O(N__17659),
            .I(\this_vga_signals.N_968_cascade_ ));
    InMux I__2273 (
            .O(N__17656),
            .I(N__17650));
    InMux I__2272 (
            .O(N__17655),
            .I(N__17650));
    LocalMux I__2271 (
            .O(N__17650),
            .I(N__17646));
    InMux I__2270 (
            .O(N__17649),
            .I(N__17643));
    Odrv4 I__2269 (
            .O(N__17646),
            .I(\this_vga_signals.N_291_0 ));
    LocalMux I__2268 (
            .O(N__17643),
            .I(\this_vga_signals.N_291_0 ));
    CascadeMux I__2267 (
            .O(N__17638),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_ ));
    InMux I__2266 (
            .O(N__17635),
            .I(N__17629));
    InMux I__2265 (
            .O(N__17634),
            .I(N__17629));
    LocalMux I__2264 (
            .O(N__17629),
            .I(\this_vga_signals.mult1_un68_sum_axb1 ));
    InMux I__2263 (
            .O(N__17626),
            .I(N__17623));
    LocalMux I__2262 (
            .O(N__17623),
            .I(\this_vga_signals.mult1_un68_sum_ac0_2 ));
    CascadeMux I__2261 (
            .O(N__17620),
            .I(\this_vga_signals.mult1_un68_sum_axb1_cascade_ ));
    InMux I__2260 (
            .O(N__17617),
            .I(N__17613));
    InMux I__2259 (
            .O(N__17616),
            .I(N__17610));
    LocalMux I__2258 (
            .O(N__17613),
            .I(\this_vga_signals.mult1_un68_sum_axb2 ));
    LocalMux I__2257 (
            .O(N__17610),
            .I(\this_vga_signals.mult1_un68_sum_axb2 ));
    InMux I__2256 (
            .O(N__17605),
            .I(N__17601));
    InMux I__2255 (
            .O(N__17604),
            .I(N__17598));
    LocalMux I__2254 (
            .O(N__17601),
            .I(N__17595));
    LocalMux I__2253 (
            .O(N__17598),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    Odrv4 I__2252 (
            .O(N__17595),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    InMux I__2251 (
            .O(N__17590),
            .I(N__17587));
    LocalMux I__2250 (
            .O(N__17587),
            .I(N__17584));
    Span4Mux_h I__2249 (
            .O(N__17584),
            .I(N__17580));
    InMux I__2248 (
            .O(N__17583),
            .I(N__17577));
    Span4Mux_v I__2247 (
            .O(N__17580),
            .I(N__17572));
    LocalMux I__2246 (
            .O(N__17577),
            .I(N__17572));
    Span4Mux_h I__2245 (
            .O(N__17572),
            .I(N__17569));
    Odrv4 I__2244 (
            .O(N__17569),
            .I(M_this_oam_ram_read_data_20));
    InMux I__2243 (
            .O(N__17566),
            .I(N__17563));
    LocalMux I__2242 (
            .O(N__17563),
            .I(N__17560));
    Span4Mux_v I__2241 (
            .O(N__17560),
            .I(N__17557));
    Span4Mux_h I__2240 (
            .O(N__17557),
            .I(N__17554));
    Odrv4 I__2239 (
            .O(N__17554),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_20 ));
    InMux I__2238 (
            .O(N__17551),
            .I(N__17548));
    LocalMux I__2237 (
            .O(N__17548),
            .I(N__17545));
    Span4Mux_v I__2236 (
            .O(N__17545),
            .I(N__17542));
    Odrv4 I__2235 (
            .O(N__17542),
            .I(\this_ppu.oam_cache.mem_13 ));
    CascadeMux I__2234 (
            .O(N__17539),
            .I(N__17536));
    InMux I__2233 (
            .O(N__17536),
            .I(N__17533));
    LocalMux I__2232 (
            .O(N__17533),
            .I(N__17530));
    Odrv12 I__2231 (
            .O(N__17530),
            .I(M_this_vga_signals_address_4));
    InMux I__2230 (
            .O(N__17527),
            .I(bfn_12_18_0_));
    CascadeMux I__2229 (
            .O(N__17524),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_ ));
    InMux I__2228 (
            .O(N__17521),
            .I(N__17518));
    LocalMux I__2227 (
            .O(N__17518),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz ));
    InMux I__2226 (
            .O(N__17515),
            .I(N__17512));
    LocalMux I__2225 (
            .O(N__17512),
            .I(N__17509));
    Span4Mux_h I__2224 (
            .O(N__17509),
            .I(N__17505));
    InMux I__2223 (
            .O(N__17508),
            .I(N__17502));
    Odrv4 I__2222 (
            .O(N__17505),
            .I(\this_ppu.N_1184_7 ));
    LocalMux I__2221 (
            .O(N__17502),
            .I(\this_ppu.N_1184_7 ));
    InMux I__2220 (
            .O(N__17497),
            .I(N__17494));
    LocalMux I__2219 (
            .O(N__17494),
            .I(N__17491));
    Odrv4 I__2218 (
            .O(N__17491),
            .I(\this_ppu.un1_M_state_q_7_i_0 ));
    InMux I__2217 (
            .O(N__17488),
            .I(N__17485));
    LocalMux I__2216 (
            .O(N__17485),
            .I(N__17482));
    Span12Mux_v I__2215 (
            .O(N__17482),
            .I(N__17479));
    Odrv12 I__2214 (
            .O(N__17479),
            .I(M_this_oam_ram_read_data_11));
    InMux I__2213 (
            .O(N__17476),
            .I(N__17473));
    LocalMux I__2212 (
            .O(N__17473),
            .I(N__17470));
    Span4Mux_h I__2211 (
            .O(N__17470),
            .I(N__17467));
    Odrv4 I__2210 (
            .O(N__17467),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_11 ));
    InMux I__2209 (
            .O(N__17464),
            .I(N__17461));
    LocalMux I__2208 (
            .O(N__17461),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_12 ));
    InMux I__2207 (
            .O(N__17458),
            .I(N__17455));
    LocalMux I__2206 (
            .O(N__17455),
            .I(N__17452));
    Span4Mux_h I__2205 (
            .O(N__17452),
            .I(N__17449));
    Span4Mux_h I__2204 (
            .O(N__17449),
            .I(N__17446));
    Odrv4 I__2203 (
            .O(N__17446),
            .I(\this_ppu.oam_cache.mem_15 ));
    InMux I__2202 (
            .O(N__17443),
            .I(N__17439));
    InMux I__2201 (
            .O(N__17442),
            .I(N__17436));
    LocalMux I__2200 (
            .O(N__17439),
            .I(\this_vga_signals.N_298_0 ));
    LocalMux I__2199 (
            .O(N__17436),
            .I(\this_vga_signals.N_298_0 ));
    InMux I__2198 (
            .O(N__17431),
            .I(N__17428));
    LocalMux I__2197 (
            .O(N__17428),
            .I(\this_vga_signals.hsync_1_i_0_0_a3_0 ));
    InMux I__2196 (
            .O(N__17425),
            .I(N__17422));
    LocalMux I__2195 (
            .O(N__17422),
            .I(N__17419));
    Span4Mux_h I__2194 (
            .O(N__17419),
            .I(N__17413));
    CascadeMux I__2193 (
            .O(N__17418),
            .I(N__17410));
    InMux I__2192 (
            .O(N__17417),
            .I(N__17405));
    InMux I__2191 (
            .O(N__17416),
            .I(N__17402));
    Span4Mux_v I__2190 (
            .O(N__17413),
            .I(N__17399));
    InMux I__2189 (
            .O(N__17410),
            .I(N__17392));
    InMux I__2188 (
            .O(N__17409),
            .I(N__17392));
    InMux I__2187 (
            .O(N__17408),
            .I(N__17392));
    LocalMux I__2186 (
            .O(N__17405),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__2185 (
            .O(N__17402),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    Odrv4 I__2184 (
            .O(N__17399),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__2183 (
            .O(N__17392),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    InMux I__2182 (
            .O(N__17383),
            .I(N__17380));
    LocalMux I__2181 (
            .O(N__17380),
            .I(N__17375));
    InMux I__2180 (
            .O(N__17379),
            .I(N__17372));
    CascadeMux I__2179 (
            .O(N__17378),
            .I(N__17369));
    Span4Mux_h I__2178 (
            .O(N__17375),
            .I(N__17365));
    LocalMux I__2177 (
            .O(N__17372),
            .I(N__17362));
    InMux I__2176 (
            .O(N__17369),
            .I(N__17359));
    CascadeMux I__2175 (
            .O(N__17368),
            .I(N__17355));
    Span4Mux_h I__2174 (
            .O(N__17365),
            .I(N__17348));
    Span4Mux_h I__2173 (
            .O(N__17362),
            .I(N__17348));
    LocalMux I__2172 (
            .O(N__17359),
            .I(N__17348));
    InMux I__2171 (
            .O(N__17358),
            .I(N__17342));
    InMux I__2170 (
            .O(N__17355),
            .I(N__17339));
    Span4Mux_v I__2169 (
            .O(N__17348),
            .I(N__17336));
    InMux I__2168 (
            .O(N__17347),
            .I(N__17329));
    InMux I__2167 (
            .O(N__17346),
            .I(N__17329));
    InMux I__2166 (
            .O(N__17345),
            .I(N__17329));
    LocalMux I__2165 (
            .O(N__17342),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2164 (
            .O(N__17339),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__2163 (
            .O(N__17336),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2162 (
            .O(N__17329),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    InMux I__2161 (
            .O(N__17320),
            .I(N__17314));
    InMux I__2160 (
            .O(N__17319),
            .I(N__17307));
    InMux I__2159 (
            .O(N__17318),
            .I(N__17307));
    InMux I__2158 (
            .O(N__17317),
            .I(N__17307));
    LocalMux I__2157 (
            .O(N__17314),
            .I(N__17299));
    LocalMux I__2156 (
            .O(N__17307),
            .I(N__17299));
    InMux I__2155 (
            .O(N__17306),
            .I(N__17294));
    InMux I__2154 (
            .O(N__17305),
            .I(N__17294));
    InMux I__2153 (
            .O(N__17304),
            .I(N__17291));
    Span4Mux_v I__2152 (
            .O(N__17299),
            .I(N__17288));
    LocalMux I__2151 (
            .O(N__17294),
            .I(N__17285));
    LocalMux I__2150 (
            .O(N__17291),
            .I(N__17277));
    Span4Mux_h I__2149 (
            .O(N__17288),
            .I(N__17277));
    Span4Mux_v I__2148 (
            .O(N__17285),
            .I(N__17277));
    InMux I__2147 (
            .O(N__17284),
            .I(N__17274));
    Odrv4 I__2146 (
            .O(N__17277),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2145 (
            .O(N__17274),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__2144 (
            .O(N__17269),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__2143 (
            .O(N__17266),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__2142 (
            .O(N__17263),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__2141 (
            .O(N__17260),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__2140 (
            .O(N__17257),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__2139 (
            .O(N__17254),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__2138 (
            .O(N__17251),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__2137 (
            .O(N__17248),
            .I(N__17245));
    LocalMux I__2136 (
            .O(N__17245),
            .I(N__17242));
    Odrv4 I__2135 (
            .O(N__17242),
            .I(M_this_data_tmp_qZ0Z_20));
    InMux I__2134 (
            .O(N__17239),
            .I(N__17236));
    LocalMux I__2133 (
            .O(N__17236),
            .I(N__17233));
    Odrv4 I__2132 (
            .O(N__17233),
            .I(M_this_data_tmp_qZ0Z_18));
    InMux I__2131 (
            .O(N__17230),
            .I(N__17227));
    LocalMux I__2130 (
            .O(N__17227),
            .I(N__17224));
    Span4Mux_h I__2129 (
            .O(N__17224),
            .I(N__17221));
    Odrv4 I__2128 (
            .O(N__17221),
            .I(M_this_oam_ram_write_data_0));
    InMux I__2127 (
            .O(N__17218),
            .I(N__17213));
    InMux I__2126 (
            .O(N__17217),
            .I(N__17208));
    InMux I__2125 (
            .O(N__17216),
            .I(N__17208));
    LocalMux I__2124 (
            .O(N__17213),
            .I(N__17201));
    LocalMux I__2123 (
            .O(N__17208),
            .I(N__17201));
    InMux I__2122 (
            .O(N__17207),
            .I(N__17198));
    InMux I__2121 (
            .O(N__17206),
            .I(N__17195));
    Span4Mux_v I__2120 (
            .O(N__17201),
            .I(N__17190));
    LocalMux I__2119 (
            .O(N__17198),
            .I(N__17187));
    LocalMux I__2118 (
            .O(N__17195),
            .I(N__17184));
    InMux I__2117 (
            .O(N__17194),
            .I(N__17181));
    CascadeMux I__2116 (
            .O(N__17193),
            .I(N__17178));
    Span4Mux_h I__2115 (
            .O(N__17190),
            .I(N__17171));
    Span4Mux_v I__2114 (
            .O(N__17187),
            .I(N__17171));
    Span4Mux_v I__2113 (
            .O(N__17184),
            .I(N__17171));
    LocalMux I__2112 (
            .O(N__17181),
            .I(N__17168));
    InMux I__2111 (
            .O(N__17178),
            .I(N__17165));
    Odrv4 I__2110 (
            .O(N__17171),
            .I(\this_vga_ramdac.N_852_i_reto ));
    Odrv4 I__2109 (
            .O(N__17168),
            .I(\this_vga_ramdac.N_852_i_reto ));
    LocalMux I__2108 (
            .O(N__17165),
            .I(\this_vga_ramdac.N_852_i_reto ));
    CascadeMux I__2107 (
            .O(N__17158),
            .I(\this_vga_signals.N_298_0_cascade_ ));
    InMux I__2106 (
            .O(N__17155),
            .I(N__17152));
    LocalMux I__2105 (
            .O(N__17152),
            .I(N__17149));
    Odrv4 I__2104 (
            .O(N__17149),
            .I(\this_vga_signals.M_hcounter_d7_0_i_0_o3_0_o3_4_a2_0 ));
    CascadeMux I__2103 (
            .O(N__17146),
            .I(\this_vga_signals.N_1044_0_cascade_ ));
    InMux I__2102 (
            .O(N__17143),
            .I(N__17140));
    LocalMux I__2101 (
            .O(N__17140),
            .I(M_this_data_tmp_qZ0Z_8));
    InMux I__2100 (
            .O(N__17137),
            .I(N__17134));
    LocalMux I__2099 (
            .O(N__17134),
            .I(M_this_data_tmp_qZ0Z_9));
    InMux I__2098 (
            .O(N__17131),
            .I(N__17128));
    LocalMux I__2097 (
            .O(N__17128),
            .I(N__17125));
    Odrv12 I__2096 (
            .O(N__17125),
            .I(M_this_oam_ram_write_data_26));
    InMux I__2095 (
            .O(N__17122),
            .I(N__17119));
    LocalMux I__2094 (
            .O(N__17119),
            .I(N__17116));
    Odrv4 I__2093 (
            .O(N__17116),
            .I(M_this_oam_ram_write_data_27));
    InMux I__2092 (
            .O(N__17113),
            .I(N__17110));
    LocalMux I__2091 (
            .O(N__17110),
            .I(N__17107));
    Odrv4 I__2090 (
            .O(N__17107),
            .I(M_this_oam_ram_write_data_30));
    InMux I__2089 (
            .O(N__17104),
            .I(N__17101));
    LocalMux I__2088 (
            .O(N__17101),
            .I(M_this_data_tmp_qZ0Z_15));
    InMux I__2087 (
            .O(N__17098),
            .I(N__17095));
    LocalMux I__2086 (
            .O(N__17095),
            .I(N__17092));
    Span4Mux_h I__2085 (
            .O(N__17092),
            .I(N__17089));
    Odrv4 I__2084 (
            .O(N__17089),
            .I(M_this_oam_ram_write_data_15));
    InMux I__2083 (
            .O(N__17086),
            .I(N__17083));
    LocalMux I__2082 (
            .O(N__17083),
            .I(M_this_data_tmp_qZ0Z_16));
    InMux I__2081 (
            .O(N__17080),
            .I(N__17077));
    LocalMux I__2080 (
            .O(N__17077),
            .I(N__17074));
    Span4Mux_h I__2079 (
            .O(N__17074),
            .I(N__17071));
    Odrv4 I__2078 (
            .O(N__17071),
            .I(M_this_data_tmp_qZ0Z_17));
    InMux I__2077 (
            .O(N__17068),
            .I(N__17065));
    LocalMux I__2076 (
            .O(N__17065),
            .I(N__17062));
    Odrv4 I__2075 (
            .O(N__17062),
            .I(M_this_data_tmp_qZ0Z_19));
    InMux I__2074 (
            .O(N__17059),
            .I(N__17056));
    LocalMux I__2073 (
            .O(N__17056),
            .I(N__17053));
    Odrv4 I__2072 (
            .O(N__17053),
            .I(\this_ppu.un1_oam_data_1_axb_7 ));
    InMux I__2071 (
            .O(N__17050),
            .I(N__17047));
    LocalMux I__2070 (
            .O(N__17047),
            .I(N__17044));
    Span4Mux_v I__2069 (
            .O(N__17044),
            .I(N__17041));
    Span4Mux_h I__2068 (
            .O(N__17041),
            .I(N__17038));
    Odrv4 I__2067 (
            .O(N__17038),
            .I(M_this_oam_ram_write_data_6));
    InMux I__2066 (
            .O(N__17035),
            .I(N__17032));
    LocalMux I__2065 (
            .O(N__17032),
            .I(M_this_data_tmp_qZ0Z_6));
    InMux I__2064 (
            .O(N__17029),
            .I(N__17026));
    LocalMux I__2063 (
            .O(N__17026),
            .I(N__17023));
    Span4Mux_h I__2062 (
            .O(N__17023),
            .I(N__17020));
    Odrv4 I__2061 (
            .O(N__17020),
            .I(M_this_oam_ram_write_data_7));
    InMux I__2060 (
            .O(N__17017),
            .I(N__17014));
    LocalMux I__2059 (
            .O(N__17014),
            .I(M_this_data_tmp_qZ0Z_7));
    InMux I__2058 (
            .O(N__17011),
            .I(N__17007));
    InMux I__2057 (
            .O(N__17010),
            .I(N__17004));
    LocalMux I__2056 (
            .O(N__17007),
            .I(N__17001));
    LocalMux I__2055 (
            .O(N__17004),
            .I(N__16998));
    Span4Mux_h I__2054 (
            .O(N__17001),
            .I(N__16995));
    Span12Mux_v I__2053 (
            .O(N__16998),
            .I(N__16992));
    Odrv4 I__2052 (
            .O(N__16995),
            .I(M_this_oam_ram_read_data_17));
    Odrv12 I__2051 (
            .O(N__16992),
            .I(M_this_oam_ram_read_data_17));
    InMux I__2050 (
            .O(N__16987),
            .I(N__16984));
    LocalMux I__2049 (
            .O(N__16984),
            .I(N__16981));
    Span12Mux_v I__2048 (
            .O(N__16981),
            .I(N__16978));
    Odrv12 I__2047 (
            .O(N__16978),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_17 ));
    InMux I__2046 (
            .O(N__16975),
            .I(N__16972));
    LocalMux I__2045 (
            .O(N__16972),
            .I(M_this_data_tmp_qZ0Z_10));
    CascadeMux I__2044 (
            .O(N__16969),
            .I(\this_vga_signals.mult1_un68_sum_ac0_2_cascade_ ));
    InMux I__2043 (
            .O(N__16966),
            .I(N__16963));
    LocalMux I__2042 (
            .O(N__16963),
            .I(\this_vga_signals.mult1_un68_sum_c3_1 ));
    InMux I__2041 (
            .O(N__16960),
            .I(N__16952));
    InMux I__2040 (
            .O(N__16959),
            .I(N__16947));
    InMux I__2039 (
            .O(N__16958),
            .I(N__16947));
    InMux I__2038 (
            .O(N__16957),
            .I(N__16942));
    InMux I__2037 (
            .O(N__16956),
            .I(N__16942));
    InMux I__2036 (
            .O(N__16955),
            .I(N__16939));
    LocalMux I__2035 (
            .O(N__16952),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    LocalMux I__2034 (
            .O(N__16947),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    LocalMux I__2033 (
            .O(N__16942),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    LocalMux I__2032 (
            .O(N__16939),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    InMux I__2031 (
            .O(N__16930),
            .I(N__16927));
    LocalMux I__2030 (
            .O(N__16927),
            .I(\this_vga_signals.mult1_un75_sum_c2_0 ));
    CascadeMux I__2029 (
            .O(N__16924),
            .I(\this_vga_signals.mult1_un75_sum_c2_0_cascade_ ));
    InMux I__2028 (
            .O(N__16921),
            .I(N__16918));
    LocalMux I__2027 (
            .O(N__16918),
            .I(\this_vga_signals.if_N_8_i ));
    InMux I__2026 (
            .O(N__16915),
            .I(N__16912));
    LocalMux I__2025 (
            .O(N__16912),
            .I(N__16909));
    Span4Mux_v I__2024 (
            .O(N__16909),
            .I(N__16906));
    Odrv4 I__2023 (
            .O(N__16906),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    InMux I__2022 (
            .O(N__16903),
            .I(N__16900));
    LocalMux I__2021 (
            .O(N__16900),
            .I(N__16897));
    Span4Mux_v I__2020 (
            .O(N__16897),
            .I(N__16894));
    Span4Mux_h I__2019 (
            .O(N__16894),
            .I(N__16891));
    Odrv4 I__2018 (
            .O(N__16891),
            .I(M_this_oam_ram_read_data_27));
    InMux I__2017 (
            .O(N__16888),
            .I(N__16885));
    LocalMux I__2016 (
            .O(N__16885),
            .I(N__16882));
    Span4Mux_h I__2015 (
            .O(N__16882),
            .I(N__16879));
    Odrv4 I__2014 (
            .O(N__16879),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_27 ));
    InMux I__2013 (
            .O(N__16876),
            .I(N__16873));
    LocalMux I__2012 (
            .O(N__16873),
            .I(N__16870));
    Span4Mux_v I__2011 (
            .O(N__16870),
            .I(N__16867));
    Odrv4 I__2010 (
            .O(N__16867),
            .I(\this_ppu.oam_cache.mem_0 ));
    InMux I__2009 (
            .O(N__16864),
            .I(N__16861));
    LocalMux I__2008 (
            .O(N__16861),
            .I(N__16857));
    InMux I__2007 (
            .O(N__16860),
            .I(N__16854));
    Span4Mux_h I__2006 (
            .O(N__16857),
            .I(N__16851));
    LocalMux I__2005 (
            .O(N__16854),
            .I(N__16848));
    Span4Mux_v I__2004 (
            .O(N__16851),
            .I(N__16845));
    Odrv4 I__2003 (
            .O(N__16848),
            .I(M_this_oam_ram_read_data_2));
    Odrv4 I__2002 (
            .O(N__16845),
            .I(M_this_oam_ram_read_data_2));
    InMux I__2001 (
            .O(N__16840),
            .I(N__16837));
    LocalMux I__2000 (
            .O(N__16837),
            .I(N__16834));
    Span4Mux_h I__1999 (
            .O(N__16834),
            .I(N__16831));
    Odrv4 I__1998 (
            .O(N__16831),
            .I(\this_ppu.m28_e_i_a3_4 ));
    InMux I__1997 (
            .O(N__16828),
            .I(N__16825));
    LocalMux I__1996 (
            .O(N__16825),
            .I(\this_ppu.m28_e_i_a3_3 ));
    CascadeMux I__1995 (
            .O(N__16822),
            .I(\this_ppu.N_1184_7_cascade_ ));
    InMux I__1994 (
            .O(N__16819),
            .I(N__16816));
    LocalMux I__1993 (
            .O(N__16816),
            .I(\this_ppu.m18_i_1 ));
    InMux I__1992 (
            .O(N__16813),
            .I(N__16810));
    LocalMux I__1991 (
            .O(N__16810),
            .I(N__16806));
    InMux I__1990 (
            .O(N__16809),
            .I(N__16803));
    Odrv4 I__1989 (
            .O(N__16806),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_2 ));
    LocalMux I__1988 (
            .O(N__16803),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_2 ));
    InMux I__1987 (
            .O(N__16798),
            .I(N__16795));
    LocalMux I__1986 (
            .O(N__16795),
            .I(N__16792));
    Span4Mux_v I__1985 (
            .O(N__16792),
            .I(N__16789));
    Odrv4 I__1984 (
            .O(N__16789),
            .I(\this_ppu.oam_cache.mem_12 ));
    CascadeMux I__1983 (
            .O(N__16786),
            .I(N__16782));
    InMux I__1982 (
            .O(N__16785),
            .I(N__16777));
    InMux I__1981 (
            .O(N__16782),
            .I(N__16777));
    LocalMux I__1980 (
            .O(N__16777),
            .I(N__16774));
    Span4Mux_h I__1979 (
            .O(N__16774),
            .I(N__16771));
    Span4Mux_v I__1978 (
            .O(N__16771),
            .I(N__16768));
    Odrv4 I__1977 (
            .O(N__16768),
            .I(M_this_oam_ram_read_data_5));
    InMux I__1976 (
            .O(N__16765),
            .I(N__16762));
    LocalMux I__1975 (
            .O(N__16762),
            .I(N__16759));
    Span4Mux_h I__1974 (
            .O(N__16759),
            .I(N__16756));
    Odrv4 I__1973 (
            .O(N__16756),
            .I(\this_ppu.oam_cache.N_569_0 ));
    InMux I__1972 (
            .O(N__16753),
            .I(N__16749));
    InMux I__1971 (
            .O(N__16752),
            .I(N__16746));
    LocalMux I__1970 (
            .O(N__16749),
            .I(N__16741));
    LocalMux I__1969 (
            .O(N__16746),
            .I(N__16741));
    Span4Mux_h I__1968 (
            .O(N__16741),
            .I(N__16738));
    Span4Mux_v I__1967 (
            .O(N__16738),
            .I(N__16735));
    Odrv4 I__1966 (
            .O(N__16735),
            .I(M_this_oam_ram_read_data_4));
    InMux I__1965 (
            .O(N__16732),
            .I(N__16729));
    LocalMux I__1964 (
            .O(N__16729),
            .I(N__16726));
    Span4Mux_h I__1963 (
            .O(N__16726),
            .I(N__16723));
    Odrv4 I__1962 (
            .O(N__16723),
            .I(\this_ppu.oam_cache.N_575_0 ));
    InMux I__1961 (
            .O(N__16720),
            .I(N__16717));
    LocalMux I__1960 (
            .O(N__16717),
            .I(\this_ppu.N_1182 ));
    CascadeMux I__1959 (
            .O(N__16714),
            .I(\this_vga_signals.if_N_9_0_0_cascade_ ));
    InMux I__1958 (
            .O(N__16711),
            .I(N__16708));
    LocalMux I__1957 (
            .O(N__16708),
            .I(\this_vga_signals.mult1_un82_sum_c3 ));
    InMux I__1956 (
            .O(N__16705),
            .I(N__16702));
    LocalMux I__1955 (
            .O(N__16702),
            .I(\this_vga_signals.N_811_0 ));
    IoInMux I__1954 (
            .O(N__16699),
            .I(N__16696));
    LocalMux I__1953 (
            .O(N__16696),
            .I(N__16693));
    Span4Mux_s3_h I__1952 (
            .O(N__16693),
            .I(N__16690));
    Span4Mux_v I__1951 (
            .O(N__16690),
            .I(N__16687));
    Span4Mux_v I__1950 (
            .O(N__16687),
            .I(N__16684));
    Span4Mux_h I__1949 (
            .O(N__16684),
            .I(N__16681));
    Odrv4 I__1948 (
            .O(N__16681),
            .I(rgb_c_3));
    CascadeMux I__1947 (
            .O(N__16678),
            .I(N__16675));
    CascadeBuf I__1946 (
            .O(N__16675),
            .I(N__16672));
    CascadeMux I__1945 (
            .O(N__16672),
            .I(N__16669));
    InMux I__1944 (
            .O(N__16669),
            .I(N__16666));
    LocalMux I__1943 (
            .O(N__16666),
            .I(N__16663));
    Span4Mux_h I__1942 (
            .O(N__16663),
            .I(N__16657));
    InMux I__1941 (
            .O(N__16662),
            .I(N__16652));
    InMux I__1940 (
            .O(N__16661),
            .I(N__16652));
    InMux I__1939 (
            .O(N__16660),
            .I(N__16649));
    Span4Mux_v I__1938 (
            .O(N__16657),
            .I(N__16646));
    LocalMux I__1937 (
            .O(N__16652),
            .I(M_this_ppu_oam_addr_5));
    LocalMux I__1936 (
            .O(N__16649),
            .I(M_this_ppu_oam_addr_5));
    Odrv4 I__1935 (
            .O(N__16646),
            .I(M_this_ppu_oam_addr_5));
    CascadeMux I__1934 (
            .O(N__16639),
            .I(N__16636));
    CascadeBuf I__1933 (
            .O(N__16636),
            .I(N__16633));
    CascadeMux I__1932 (
            .O(N__16633),
            .I(N__16628));
    CascadeMux I__1931 (
            .O(N__16632),
            .I(N__16625));
    InMux I__1930 (
            .O(N__16631),
            .I(N__16620));
    InMux I__1929 (
            .O(N__16628),
            .I(N__16617));
    InMux I__1928 (
            .O(N__16625),
            .I(N__16610));
    InMux I__1927 (
            .O(N__16624),
            .I(N__16610));
    InMux I__1926 (
            .O(N__16623),
            .I(N__16610));
    LocalMux I__1925 (
            .O(N__16620),
            .I(N__16604));
    LocalMux I__1924 (
            .O(N__16617),
            .I(N__16601));
    LocalMux I__1923 (
            .O(N__16610),
            .I(N__16598));
    InMux I__1922 (
            .O(N__16609),
            .I(N__16593));
    InMux I__1921 (
            .O(N__16608),
            .I(N__16593));
    InMux I__1920 (
            .O(N__16607),
            .I(N__16590));
    Span4Mux_h I__1919 (
            .O(N__16604),
            .I(N__16585));
    Span4Mux_v I__1918 (
            .O(N__16601),
            .I(N__16585));
    Odrv4 I__1917 (
            .O(N__16598),
            .I(M_this_ppu_oam_addr_0));
    LocalMux I__1916 (
            .O(N__16593),
            .I(M_this_ppu_oam_addr_0));
    LocalMux I__1915 (
            .O(N__16590),
            .I(M_this_ppu_oam_addr_0));
    Odrv4 I__1914 (
            .O(N__16585),
            .I(M_this_ppu_oam_addr_0));
    InMux I__1913 (
            .O(N__16576),
            .I(N__16573));
    LocalMux I__1912 (
            .O(N__16573),
            .I(N__16570));
    Odrv4 I__1911 (
            .O(N__16570),
            .I(\this_ppu.m35_i_0_a3_1_3 ));
    InMux I__1910 (
            .O(N__16567),
            .I(N__16563));
    InMux I__1909 (
            .O(N__16566),
            .I(N__16560));
    LocalMux I__1908 (
            .O(N__16563),
            .I(N__16557));
    LocalMux I__1907 (
            .O(N__16560),
            .I(N__16554));
    Odrv4 I__1906 (
            .O(N__16557),
            .I(\this_ppu.N_1394 ));
    Odrv4 I__1905 (
            .O(N__16554),
            .I(\this_ppu.N_1394 ));
    InMux I__1904 (
            .O(N__16549),
            .I(N__16546));
    LocalMux I__1903 (
            .O(N__16546),
            .I(N__16543));
    Span4Mux_h I__1902 (
            .O(N__16543),
            .I(N__16540));
    Odrv4 I__1901 (
            .O(N__16540),
            .I(M_this_oam_ram_write_data_9));
    InMux I__1900 (
            .O(N__16537),
            .I(N__16534));
    LocalMux I__1899 (
            .O(N__16534),
            .I(N__16531));
    Odrv4 I__1898 (
            .O(N__16531),
            .I(M_this_oam_ram_read_data_i_20));
    InMux I__1897 (
            .O(N__16528),
            .I(N__16525));
    LocalMux I__1896 (
            .O(N__16525),
            .I(N__16522));
    Odrv4 I__1895 (
            .O(N__16522),
            .I(M_this_oam_ram_write_data_28));
    InMux I__1894 (
            .O(N__16519),
            .I(N__16516));
    LocalMux I__1893 (
            .O(N__16516),
            .I(N__16513));
    Span4Mux_h I__1892 (
            .O(N__16513),
            .I(N__16510));
    Odrv4 I__1891 (
            .O(N__16510),
            .I(M_this_oam_ram_write_data_8));
    InMux I__1890 (
            .O(N__16507),
            .I(N__16504));
    LocalMux I__1889 (
            .O(N__16504),
            .I(N__16501));
    Odrv4 I__1888 (
            .O(N__16501),
            .I(M_this_oam_ram_write_data_31));
    InMux I__1887 (
            .O(N__16498),
            .I(N__16495));
    LocalMux I__1886 (
            .O(N__16495),
            .I(N__16492));
    Odrv4 I__1885 (
            .O(N__16492),
            .I(M_this_oam_ram_write_data_16));
    InMux I__1884 (
            .O(N__16489),
            .I(N__16486));
    LocalMux I__1883 (
            .O(N__16486),
            .I(N__16483));
    Span4Mux_h I__1882 (
            .O(N__16483),
            .I(N__16480));
    Odrv4 I__1881 (
            .O(N__16480),
            .I(M_this_oam_ram_write_data_24));
    InMux I__1880 (
            .O(N__16477),
            .I(N__16474));
    LocalMux I__1879 (
            .O(N__16474),
            .I(N__16471));
    Sp12to4 I__1878 (
            .O(N__16471),
            .I(N__16468));
    Odrv12 I__1877 (
            .O(N__16468),
            .I(\this_vga_signals.hsync_1_i_0_0_1 ));
    InMux I__1876 (
            .O(N__16465),
            .I(N__16462));
    LocalMux I__1875 (
            .O(N__16462),
            .I(N__16459));
    Span4Mux_h I__1874 (
            .O(N__16459),
            .I(N__16456));
    Span4Mux_v I__1873 (
            .O(N__16456),
            .I(N__16453));
    Odrv4 I__1872 (
            .O(N__16453),
            .I(M_this_oam_ram_read_data_14));
    InMux I__1871 (
            .O(N__16450),
            .I(N__16447));
    LocalMux I__1870 (
            .O(N__16447),
            .I(N__16444));
    Span4Mux_h I__1869 (
            .O(N__16444),
            .I(N__16441));
    Odrv4 I__1868 (
            .O(N__16441),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_14 ));
    InMux I__1867 (
            .O(N__16438),
            .I(N__16435));
    LocalMux I__1866 (
            .O(N__16435),
            .I(\this_vga_signals.hsync_1_i_0_0_a3_0_0 ));
    InMux I__1865 (
            .O(N__16432),
            .I(N__16429));
    LocalMux I__1864 (
            .O(N__16429),
            .I(N__16426));
    Span12Mux_h I__1863 (
            .O(N__16426),
            .I(N__16423));
    Odrv12 I__1862 (
            .O(N__16423),
            .I(M_this_oam_ram_read_data_29));
    InMux I__1861 (
            .O(N__16420),
            .I(N__16417));
    LocalMux I__1860 (
            .O(N__16417),
            .I(N__16414));
    Span4Mux_h I__1859 (
            .O(N__16414),
            .I(N__16411));
    Odrv4 I__1858 (
            .O(N__16411),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_29 ));
    InMux I__1857 (
            .O(N__16408),
            .I(N__16404));
    InMux I__1856 (
            .O(N__16407),
            .I(N__16401));
    LocalMux I__1855 (
            .O(N__16404),
            .I(N__16398));
    LocalMux I__1854 (
            .O(N__16401),
            .I(N__16395));
    Span4Mux_v I__1853 (
            .O(N__16398),
            .I(N__16392));
    Span4Mux_h I__1852 (
            .O(N__16395),
            .I(N__16389));
    Odrv4 I__1851 (
            .O(N__16392),
            .I(M_this_oam_ram_read_data_21));
    Odrv4 I__1850 (
            .O(N__16389),
            .I(M_this_oam_ram_read_data_21));
    CascadeMux I__1849 (
            .O(N__16384),
            .I(N__16381));
    InMux I__1848 (
            .O(N__16381),
            .I(N__16378));
    LocalMux I__1847 (
            .O(N__16378),
            .I(M_this_oam_ram_read_data_i_21));
    InMux I__1846 (
            .O(N__16375),
            .I(N__16372));
    LocalMux I__1845 (
            .O(N__16372),
            .I(N__16369));
    Span4Mux_h I__1844 (
            .O(N__16369),
            .I(N__16366));
    Odrv4 I__1843 (
            .O(N__16366),
            .I(M_this_oam_ram_read_data_31));
    InMux I__1842 (
            .O(N__16363),
            .I(N__16360));
    LocalMux I__1841 (
            .O(N__16360),
            .I(N__16357));
    Span4Mux_h I__1840 (
            .O(N__16357),
            .I(N__16354));
    Odrv4 I__1839 (
            .O(N__16354),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_31 ));
    InMux I__1838 (
            .O(N__16351),
            .I(N__16348));
    LocalMux I__1837 (
            .O(N__16348),
            .I(N__16345));
    Span4Mux_h I__1836 (
            .O(N__16345),
            .I(N__16342));
    Odrv4 I__1835 (
            .O(N__16342),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_19 ));
    InMux I__1834 (
            .O(N__16339),
            .I(N__16333));
    InMux I__1833 (
            .O(N__16338),
            .I(N__16333));
    LocalMux I__1832 (
            .O(N__16333),
            .I(N__16330));
    Span4Mux_v I__1831 (
            .O(N__16330),
            .I(N__16327));
    Odrv4 I__1830 (
            .O(N__16327),
            .I(M_this_oam_ram_read_data_19));
    InMux I__1829 (
            .O(N__16324),
            .I(N__16321));
    LocalMux I__1828 (
            .O(N__16321),
            .I(M_this_oam_ram_read_data_i_19));
    InMux I__1827 (
            .O(N__16318),
            .I(N__16315));
    LocalMux I__1826 (
            .O(N__16315),
            .I(N__16312));
    Span4Mux_h I__1825 (
            .O(N__16312),
            .I(N__16309));
    Odrv4 I__1824 (
            .O(N__16309),
            .I(M_this_oam_ram_write_data_10));
    IoInMux I__1823 (
            .O(N__16306),
            .I(N__16303));
    LocalMux I__1822 (
            .O(N__16303),
            .I(N__16300));
    Span12Mux_s8_v I__1821 (
            .O(N__16300),
            .I(N__16297));
    Odrv12 I__1820 (
            .O(N__16297),
            .I(N_260));
    InMux I__1819 (
            .O(N__16294),
            .I(N__16291));
    LocalMux I__1818 (
            .O(N__16291),
            .I(N__16288));
    Span4Mux_h I__1817 (
            .O(N__16288),
            .I(N__16285));
    Odrv4 I__1816 (
            .O(N__16285),
            .I(M_this_oam_ram_read_data_28));
    InMux I__1815 (
            .O(N__16282),
            .I(N__16279));
    LocalMux I__1814 (
            .O(N__16279),
            .I(N__16276));
    Span12Mux_v I__1813 (
            .O(N__16276),
            .I(N__16273));
    Odrv12 I__1812 (
            .O(N__16273),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_28 ));
    InMux I__1811 (
            .O(N__16270),
            .I(N__16267));
    LocalMux I__1810 (
            .O(N__16267),
            .I(\this_ppu.M_this_oam_ram_read_data_i_18 ));
    InMux I__1809 (
            .O(N__16264),
            .I(\this_ppu.un1_oam_data_1_cry_2 ));
    InMux I__1808 (
            .O(N__16261),
            .I(\this_ppu.un1_oam_data_1_cry_3 ));
    InMux I__1807 (
            .O(N__16258),
            .I(N__16255));
    LocalMux I__1806 (
            .O(N__16255),
            .I(N__16251));
    InMux I__1805 (
            .O(N__16254),
            .I(N__16248));
    Odrv12 I__1804 (
            .O(N__16251),
            .I(\this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0 ));
    LocalMux I__1803 (
            .O(N__16248),
            .I(\this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0 ));
    InMux I__1802 (
            .O(N__16243),
            .I(\this_ppu.un1_oam_data_1_cry_4 ));
    InMux I__1801 (
            .O(N__16240),
            .I(N__16237));
    LocalMux I__1800 (
            .O(N__16237),
            .I(N__16234));
    Span4Mux_v I__1799 (
            .O(N__16234),
            .I(N__16230));
    InMux I__1798 (
            .O(N__16233),
            .I(N__16227));
    Odrv4 I__1797 (
            .O(N__16230),
            .I(\this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0 ));
    LocalMux I__1796 (
            .O(N__16227),
            .I(\this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0 ));
    InMux I__1795 (
            .O(N__16222),
            .I(\this_ppu.un1_oam_data_1_cry_5 ));
    InMux I__1794 (
            .O(N__16219),
            .I(N__16216));
    LocalMux I__1793 (
            .O(N__16216),
            .I(\this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0 ));
    CascadeMux I__1792 (
            .O(N__16213),
            .I(N__16210));
    InMux I__1791 (
            .O(N__16210),
            .I(N__16207));
    LocalMux I__1790 (
            .O(N__16207),
            .I(\this_ppu.un1_oam_data_1_cry_2_c_RNIR4HDZ0 ));
    InMux I__1789 (
            .O(N__16204),
            .I(\this_ppu.un1_oam_data_1_cry_6 ));
    InMux I__1788 (
            .O(N__16201),
            .I(N__16198));
    LocalMux I__1787 (
            .O(N__16198),
            .I(N__16195));
    Span4Mux_v I__1786 (
            .O(N__16195),
            .I(N__16191));
    InMux I__1785 (
            .O(N__16194),
            .I(N__16188));
    Odrv4 I__1784 (
            .O(N__16191),
            .I(\this_ppu.m28_e_i_o3_2 ));
    LocalMux I__1783 (
            .O(N__16188),
            .I(\this_ppu.m28_e_i_o3_2 ));
    InMux I__1782 (
            .O(N__16183),
            .I(N__16179));
    InMux I__1781 (
            .O(N__16182),
            .I(N__16176));
    LocalMux I__1780 (
            .O(N__16179),
            .I(N__16173));
    LocalMux I__1779 (
            .O(N__16176),
            .I(N__16170));
    Span4Mux_v I__1778 (
            .O(N__16173),
            .I(N__16167));
    Span4Mux_h I__1777 (
            .O(N__16170),
            .I(N__16164));
    Odrv4 I__1776 (
            .O(N__16167),
            .I(M_this_oam_ram_read_data_18));
    Odrv4 I__1775 (
            .O(N__16164),
            .I(M_this_oam_ram_read_data_18));
    InMux I__1774 (
            .O(N__16159),
            .I(N__16156));
    LocalMux I__1773 (
            .O(N__16156),
            .I(N__16153));
    Span4Mux_h I__1772 (
            .O(N__16153),
            .I(N__16150));
    Odrv4 I__1771 (
            .O(N__16150),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_18 ));
    InMux I__1770 (
            .O(N__16147),
            .I(N__16144));
    LocalMux I__1769 (
            .O(N__16144),
            .I(N__16141));
    Span4Mux_h I__1768 (
            .O(N__16141),
            .I(N__16138));
    Odrv4 I__1767 (
            .O(N__16138),
            .I(M_this_oam_ram_write_data_5));
    InMux I__1766 (
            .O(N__16135),
            .I(N__16131));
    InMux I__1765 (
            .O(N__16134),
            .I(N__16128));
    LocalMux I__1764 (
            .O(N__16131),
            .I(N__16125));
    LocalMux I__1763 (
            .O(N__16128),
            .I(N__16122));
    Span4Mux_v I__1762 (
            .O(N__16125),
            .I(N__16119));
    Span4Mux_h I__1761 (
            .O(N__16122),
            .I(N__16116));
    Odrv4 I__1760 (
            .O(N__16119),
            .I(M_this_oam_ram_read_data_22));
    Odrv4 I__1759 (
            .O(N__16116),
            .I(M_this_oam_ram_read_data_22));
    CascadeMux I__1758 (
            .O(N__16111),
            .I(N__16108));
    InMux I__1757 (
            .O(N__16108),
            .I(N__16105));
    LocalMux I__1756 (
            .O(N__16105),
            .I(M_this_oam_ram_read_data_i_22));
    CascadeMux I__1755 (
            .O(N__16102),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_cascade_ ));
    InMux I__1754 (
            .O(N__16099),
            .I(N__16093));
    InMux I__1753 (
            .O(N__16098),
            .I(N__16093));
    LocalMux I__1752 (
            .O(N__16093),
            .I(\this_vga_signals.if_m2 ));
    InMux I__1751 (
            .O(N__16090),
            .I(N__16086));
    InMux I__1750 (
            .O(N__16089),
            .I(N__16083));
    LocalMux I__1749 (
            .O(N__16086),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__1748 (
            .O(N__16083),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    CascadeMux I__1747 (
            .O(N__16078),
            .I(N__16075));
    InMux I__1746 (
            .O(N__16075),
            .I(N__16072));
    LocalMux I__1745 (
            .O(N__16072),
            .I(N__16069));
    Odrv12 I__1744 (
            .O(N__16069),
            .I(M_this_vga_signals_address_1));
    InMux I__1743 (
            .O(N__16066),
            .I(N__16063));
    LocalMux I__1742 (
            .O(N__16063),
            .I(\this_vga_signals.mult1_un75_sum_axb1 ));
    CascadeMux I__1741 (
            .O(N__16060),
            .I(N__16057));
    CascadeBuf I__1740 (
            .O(N__16057),
            .I(N__16054));
    CascadeMux I__1739 (
            .O(N__16054),
            .I(N__16050));
    CascadeMux I__1738 (
            .O(N__16053),
            .I(N__16045));
    InMux I__1737 (
            .O(N__16050),
            .I(N__16042));
    CascadeMux I__1736 (
            .O(N__16049),
            .I(N__16039));
    InMux I__1735 (
            .O(N__16048),
            .I(N__16036));
    InMux I__1734 (
            .O(N__16045),
            .I(N__16033));
    LocalMux I__1733 (
            .O(N__16042),
            .I(N__16030));
    InMux I__1732 (
            .O(N__16039),
            .I(N__16027));
    LocalMux I__1731 (
            .O(N__16036),
            .I(N__16022));
    LocalMux I__1730 (
            .O(N__16033),
            .I(N__16022));
    Span4Mux_h I__1729 (
            .O(N__16030),
            .I(N__16019));
    LocalMux I__1728 (
            .O(N__16027),
            .I(\this_ppu.M_oam_cache_cnt_qZ1Z_0 ));
    Odrv12 I__1727 (
            .O(N__16022),
            .I(\this_ppu.M_oam_cache_cnt_qZ1Z_0 ));
    Odrv4 I__1726 (
            .O(N__16019),
            .I(\this_ppu.M_oam_cache_cnt_qZ1Z_0 ));
    CascadeMux I__1725 (
            .O(N__16012),
            .I(N__16009));
    InMux I__1724 (
            .O(N__16009),
            .I(N__16006));
    LocalMux I__1723 (
            .O(N__16006),
            .I(N__16003));
    Odrv4 I__1722 (
            .O(N__16003),
            .I(M_this_vga_signals_address_3));
    InMux I__1721 (
            .O(N__16000),
            .I(N__15996));
    InMux I__1720 (
            .O(N__15999),
            .I(N__15993));
    LocalMux I__1719 (
            .O(N__15996),
            .I(N__15990));
    LocalMux I__1718 (
            .O(N__15993),
            .I(N__15987));
    Span4Mux_h I__1717 (
            .O(N__15990),
            .I(N__15984));
    Span12Mux_v I__1716 (
            .O(N__15987),
            .I(N__15981));
    Span4Mux_v I__1715 (
            .O(N__15984),
            .I(N__15978));
    Odrv12 I__1714 (
            .O(N__15981),
            .I(M_this_oam_ram_read_data_16));
    Odrv4 I__1713 (
            .O(N__15978),
            .I(M_this_oam_ram_read_data_16));
    InMux I__1712 (
            .O(N__15973),
            .I(N__15970));
    LocalMux I__1711 (
            .O(N__15970),
            .I(\this_ppu.M_this_oam_ram_read_data_i_16 ));
    InMux I__1710 (
            .O(N__15967),
            .I(N__15964));
    LocalMux I__1709 (
            .O(N__15964),
            .I(\this_ppu.M_this_oam_ram_read_data_i_17 ));
    InMux I__1708 (
            .O(N__15961),
            .I(N__15958));
    LocalMux I__1707 (
            .O(N__15958),
            .I(N__15955));
    Span4Mux_v I__1706 (
            .O(N__15955),
            .I(N__15952));
    Span4Mux_v I__1705 (
            .O(N__15952),
            .I(N__15949));
    Odrv4 I__1704 (
            .O(N__15949),
            .I(M_this_oam_ram_read_data_24));
    InMux I__1703 (
            .O(N__15946),
            .I(N__15943));
    LocalMux I__1702 (
            .O(N__15943),
            .I(N__15940));
    Odrv4 I__1701 (
            .O(N__15940),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_24 ));
    InMux I__1700 (
            .O(N__15937),
            .I(N__15934));
    LocalMux I__1699 (
            .O(N__15934),
            .I(N__15931));
    Span4Mux_h I__1698 (
            .O(N__15931),
            .I(N__15928));
    Odrv4 I__1697 (
            .O(N__15928),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    InMux I__1696 (
            .O(N__15925),
            .I(N__15921));
    InMux I__1695 (
            .O(N__15924),
            .I(N__15918));
    LocalMux I__1694 (
            .O(N__15921),
            .I(N__15915));
    LocalMux I__1693 (
            .O(N__15918),
            .I(N__15912));
    Span4Mux_v I__1692 (
            .O(N__15915),
            .I(N__15909));
    Span4Mux_v I__1691 (
            .O(N__15912),
            .I(N__15906));
    Span4Mux_v I__1690 (
            .O(N__15909),
            .I(N__15903));
    Odrv4 I__1689 (
            .O(N__15906),
            .I(M_this_oam_ram_read_data_7));
    Odrv4 I__1688 (
            .O(N__15903),
            .I(M_this_oam_ram_read_data_7));
    CascadeMux I__1687 (
            .O(N__15898),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ));
    CascadeMux I__1686 (
            .O(N__15895),
            .I(\this_vga_signals.mult1_un82_sum_axb1_cascade_ ));
    CascadeMux I__1685 (
            .O(N__15892),
            .I(\this_vga_signals.mult1_un89_sum_c3_cascade_ ));
    InMux I__1684 (
            .O(N__15889),
            .I(N__15886));
    LocalMux I__1683 (
            .O(N__15886),
            .I(\this_vga_signals.haddress_1_0 ));
    CascadeMux I__1682 (
            .O(N__15883),
            .I(N__15880));
    InMux I__1681 (
            .O(N__15880),
            .I(N__15877));
    LocalMux I__1680 (
            .O(N__15877),
            .I(N__15874));
    Span4Mux_v I__1679 (
            .O(N__15874),
            .I(N__15871));
    Odrv4 I__1678 (
            .O(N__15871),
            .I(M_this_vga_signals_address_0));
    InMux I__1677 (
            .O(N__15868),
            .I(N__15862));
    InMux I__1676 (
            .O(N__15867),
            .I(N__15862));
    LocalMux I__1675 (
            .O(N__15862),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0_0 ));
    InMux I__1674 (
            .O(N__15859),
            .I(N__15856));
    LocalMux I__1673 (
            .O(N__15856),
            .I(\this_ppu.un1_M_oam_curr_q_1_c4 ));
    CascadeMux I__1672 (
            .O(N__15853),
            .I(N__15848));
    InMux I__1671 (
            .O(N__15852),
            .I(N__15836));
    InMux I__1670 (
            .O(N__15851),
            .I(N__15836));
    InMux I__1669 (
            .O(N__15848),
            .I(N__15836));
    InMux I__1668 (
            .O(N__15847),
            .I(N__15836));
    InMux I__1667 (
            .O(N__15846),
            .I(N__15830));
    InMux I__1666 (
            .O(N__15845),
            .I(N__15830));
    LocalMux I__1665 (
            .O(N__15836),
            .I(N__15827));
    InMux I__1664 (
            .O(N__15835),
            .I(N__15824));
    LocalMux I__1663 (
            .O(N__15830),
            .I(\this_ppu.M_oam_curr_qc_0_1 ));
    Odrv4 I__1662 (
            .O(N__15827),
            .I(\this_ppu.M_oam_curr_qc_0_1 ));
    LocalMux I__1661 (
            .O(N__15824),
            .I(\this_ppu.M_oam_curr_qc_0_1 ));
    CascadeMux I__1660 (
            .O(N__15817),
            .I(N__15814));
    InMux I__1659 (
            .O(N__15814),
            .I(N__15811));
    LocalMux I__1658 (
            .O(N__15811),
            .I(N__15808));
    Odrv4 I__1657 (
            .O(N__15808),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO ));
    CascadeMux I__1656 (
            .O(N__15805),
            .I(N__15802));
    CascadeBuf I__1655 (
            .O(N__15802),
            .I(N__15799));
    CascadeMux I__1654 (
            .O(N__15799),
            .I(N__15796));
    InMux I__1653 (
            .O(N__15796),
            .I(N__15791));
    InMux I__1652 (
            .O(N__15795),
            .I(N__15787));
    InMux I__1651 (
            .O(N__15794),
            .I(N__15784));
    LocalMux I__1650 (
            .O(N__15791),
            .I(N__15781));
    InMux I__1649 (
            .O(N__15790),
            .I(N__15778));
    LocalMux I__1648 (
            .O(N__15787),
            .I(N__15775));
    LocalMux I__1647 (
            .O(N__15784),
            .I(N__15770));
    Span4Mux_h I__1646 (
            .O(N__15781),
            .I(N__15770));
    LocalMux I__1645 (
            .O(N__15778),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_1 ));
    Odrv4 I__1644 (
            .O(N__15775),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_1 ));
    Odrv4 I__1643 (
            .O(N__15770),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_1 ));
    InMux I__1642 (
            .O(N__15763),
            .I(N__15760));
    LocalMux I__1641 (
            .O(N__15760),
            .I(\this_ppu.m62_0_a2_0_o2_1 ));
    CascadeMux I__1640 (
            .O(N__15757),
            .I(N__15754));
    CascadeBuf I__1639 (
            .O(N__15754),
            .I(N__15751));
    CascadeMux I__1638 (
            .O(N__15751),
            .I(N__15748));
    InMux I__1637 (
            .O(N__15748),
            .I(N__15743));
    InMux I__1636 (
            .O(N__15747),
            .I(N__15738));
    InMux I__1635 (
            .O(N__15746),
            .I(N__15738));
    LocalMux I__1634 (
            .O(N__15743),
            .I(N__15734));
    LocalMux I__1633 (
            .O(N__15738),
            .I(N__15729));
    InMux I__1632 (
            .O(N__15737),
            .I(N__15725));
    Span4Mux_h I__1631 (
            .O(N__15734),
            .I(N__15722));
    InMux I__1630 (
            .O(N__15733),
            .I(N__15719));
    InMux I__1629 (
            .O(N__15732),
            .I(N__15716));
    Span4Mux_h I__1628 (
            .O(N__15729),
            .I(N__15713));
    InMux I__1627 (
            .O(N__15728),
            .I(N__15710));
    LocalMux I__1626 (
            .O(N__15725),
            .I(N__15705));
    Span4Mux_v I__1625 (
            .O(N__15722),
            .I(N__15705));
    LocalMux I__1624 (
            .O(N__15719),
            .I(M_this_ppu_oam_addr_3));
    LocalMux I__1623 (
            .O(N__15716),
            .I(M_this_ppu_oam_addr_3));
    Odrv4 I__1622 (
            .O(N__15713),
            .I(M_this_ppu_oam_addr_3));
    LocalMux I__1621 (
            .O(N__15710),
            .I(M_this_ppu_oam_addr_3));
    Odrv4 I__1620 (
            .O(N__15705),
            .I(M_this_ppu_oam_addr_3));
    CascadeMux I__1619 (
            .O(N__15694),
            .I(N__15691));
    CascadeBuf I__1618 (
            .O(N__15691),
            .I(N__15688));
    CascadeMux I__1617 (
            .O(N__15688),
            .I(N__15685));
    InMux I__1616 (
            .O(N__15685),
            .I(N__15682));
    LocalMux I__1615 (
            .O(N__15682),
            .I(N__15679));
    Span4Mux_h I__1614 (
            .O(N__15679),
            .I(N__15668));
    InMux I__1613 (
            .O(N__15678),
            .I(N__15665));
    InMux I__1612 (
            .O(N__15677),
            .I(N__15662));
    InMux I__1611 (
            .O(N__15676),
            .I(N__15657));
    InMux I__1610 (
            .O(N__15675),
            .I(N__15657));
    InMux I__1609 (
            .O(N__15674),
            .I(N__15650));
    InMux I__1608 (
            .O(N__15673),
            .I(N__15650));
    InMux I__1607 (
            .O(N__15672),
            .I(N__15650));
    InMux I__1606 (
            .O(N__15671),
            .I(N__15647));
    Span4Mux_v I__1605 (
            .O(N__15668),
            .I(N__15644));
    LocalMux I__1604 (
            .O(N__15665),
            .I(M_this_ppu_oam_addr_2));
    LocalMux I__1603 (
            .O(N__15662),
            .I(M_this_ppu_oam_addr_2));
    LocalMux I__1602 (
            .O(N__15657),
            .I(M_this_ppu_oam_addr_2));
    LocalMux I__1601 (
            .O(N__15650),
            .I(M_this_ppu_oam_addr_2));
    LocalMux I__1600 (
            .O(N__15647),
            .I(M_this_ppu_oam_addr_2));
    Odrv4 I__1599 (
            .O(N__15644),
            .I(M_this_ppu_oam_addr_2));
    CascadeMux I__1598 (
            .O(N__15631),
            .I(N__15628));
    CascadeBuf I__1597 (
            .O(N__15628),
            .I(N__15625));
    CascadeMux I__1596 (
            .O(N__15625),
            .I(N__15622));
    InMux I__1595 (
            .O(N__15622),
            .I(N__15616));
    CascadeMux I__1594 (
            .O(N__15621),
            .I(N__15612));
    CascadeMux I__1593 (
            .O(N__15620),
            .I(N__15609));
    CascadeMux I__1592 (
            .O(N__15619),
            .I(N__15605));
    LocalMux I__1591 (
            .O(N__15616),
            .I(N__15602));
    InMux I__1590 (
            .O(N__15615),
            .I(N__15599));
    InMux I__1589 (
            .O(N__15612),
            .I(N__15596));
    InMux I__1588 (
            .O(N__15609),
            .I(N__15591));
    InMux I__1587 (
            .O(N__15608),
            .I(N__15591));
    InMux I__1586 (
            .O(N__15605),
            .I(N__15588));
    Span4Mux_v I__1585 (
            .O(N__15602),
            .I(N__15585));
    LocalMux I__1584 (
            .O(N__15599),
            .I(M_this_ppu_oam_addr_4));
    LocalMux I__1583 (
            .O(N__15596),
            .I(M_this_ppu_oam_addr_4));
    LocalMux I__1582 (
            .O(N__15591),
            .I(M_this_ppu_oam_addr_4));
    LocalMux I__1581 (
            .O(N__15588),
            .I(M_this_ppu_oam_addr_4));
    Odrv4 I__1580 (
            .O(N__15585),
            .I(M_this_ppu_oam_addr_4));
    InMux I__1579 (
            .O(N__15574),
            .I(N__15565));
    InMux I__1578 (
            .O(N__15573),
            .I(N__15565));
    InMux I__1577 (
            .O(N__15572),
            .I(N__15562));
    InMux I__1576 (
            .O(N__15571),
            .I(N__15557));
    InMux I__1575 (
            .O(N__15570),
            .I(N__15557));
    LocalMux I__1574 (
            .O(N__15565),
            .I(\this_ppu.un1_M_oam_curr_q_1_c2 ));
    LocalMux I__1573 (
            .O(N__15562),
            .I(\this_ppu.un1_M_oam_curr_q_1_c2 ));
    LocalMux I__1572 (
            .O(N__15557),
            .I(\this_ppu.un1_M_oam_curr_q_1_c2 ));
    InMux I__1571 (
            .O(N__15550),
            .I(N__15547));
    LocalMux I__1570 (
            .O(N__15547),
            .I(\this_ppu.un1_M_oam_curr_q_1_c5 ));
    InMux I__1569 (
            .O(N__15544),
            .I(N__15541));
    LocalMux I__1568 (
            .O(N__15541),
            .I(N__15538));
    Odrv12 I__1567 (
            .O(N__15538),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO ));
    CascadeMux I__1566 (
            .O(N__15535),
            .I(N__15532));
    CascadeBuf I__1565 (
            .O(N__15532),
            .I(N__15529));
    CascadeMux I__1564 (
            .O(N__15529),
            .I(N__15524));
    CascadeMux I__1563 (
            .O(N__15528),
            .I(N__15520));
    CascadeMux I__1562 (
            .O(N__15527),
            .I(N__15517));
    InMux I__1561 (
            .O(N__15524),
            .I(N__15514));
    InMux I__1560 (
            .O(N__15523),
            .I(N__15511));
    InMux I__1559 (
            .O(N__15520),
            .I(N__15506));
    InMux I__1558 (
            .O(N__15517),
            .I(N__15506));
    LocalMux I__1557 (
            .O(N__15514),
            .I(N__15503));
    LocalMux I__1556 (
            .O(N__15511),
            .I(N__15500));
    LocalMux I__1555 (
            .O(N__15506),
            .I(N__15495));
    Span4Mux_v I__1554 (
            .O(N__15503),
            .I(N__15495));
    Odrv12 I__1553 (
            .O(N__15500),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_3 ));
    Odrv4 I__1552 (
            .O(N__15495),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_3 ));
    InMux I__1551 (
            .O(N__15490),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_0 ));
    InMux I__1550 (
            .O(N__15487),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_1 ));
    InMux I__1549 (
            .O(N__15484),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_2 ));
    InMux I__1548 (
            .O(N__15481),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_3 ));
    InMux I__1547 (
            .O(N__15478),
            .I(N__15475));
    LocalMux I__1546 (
            .O(N__15475),
            .I(N__15472));
    Span4Mux_v I__1545 (
            .O(N__15472),
            .I(N__15469));
    Odrv4 I__1544 (
            .O(N__15469),
            .I(\this_ppu.oam_cache.mem_7 ));
    CascadeMux I__1543 (
            .O(N__15466),
            .I(N__15463));
    InMux I__1542 (
            .O(N__15463),
            .I(N__15460));
    LocalMux I__1541 (
            .O(N__15460),
            .I(N__15457));
    Span4Mux_v I__1540 (
            .O(N__15457),
            .I(N__15454));
    Odrv4 I__1539 (
            .O(N__15454),
            .I(N_41_0));
    CascadeMux I__1538 (
            .O(N__15451),
            .I(N__15448));
    CascadeBuf I__1537 (
            .O(N__15448),
            .I(N__15445));
    CascadeMux I__1536 (
            .O(N__15445),
            .I(N__15442));
    InMux I__1535 (
            .O(N__15442),
            .I(N__15436));
    CascadeMux I__1534 (
            .O(N__15441),
            .I(N__15432));
    InMux I__1533 (
            .O(N__15440),
            .I(N__15428));
    InMux I__1532 (
            .O(N__15439),
            .I(N__15425));
    LocalMux I__1531 (
            .O(N__15436),
            .I(N__15422));
    InMux I__1530 (
            .O(N__15435),
            .I(N__15419));
    InMux I__1529 (
            .O(N__15432),
            .I(N__15414));
    InMux I__1528 (
            .O(N__15431),
            .I(N__15414));
    LocalMux I__1527 (
            .O(N__15428),
            .I(N__15411));
    LocalMux I__1526 (
            .O(N__15425),
            .I(N__15408));
    Span4Mux_v I__1525 (
            .O(N__15422),
            .I(N__15405));
    LocalMux I__1524 (
            .O(N__15419),
            .I(M_this_ppu_oam_addr_1));
    LocalMux I__1523 (
            .O(N__15414),
            .I(M_this_ppu_oam_addr_1));
    Odrv4 I__1522 (
            .O(N__15411),
            .I(M_this_ppu_oam_addr_1));
    Odrv4 I__1521 (
            .O(N__15408),
            .I(M_this_ppu_oam_addr_1));
    Odrv4 I__1520 (
            .O(N__15405),
            .I(M_this_ppu_oam_addr_1));
    InMux I__1519 (
            .O(N__15394),
            .I(N__15390));
    InMux I__1518 (
            .O(N__15393),
            .I(N__15387));
    LocalMux I__1517 (
            .O(N__15390),
            .I(N__15384));
    LocalMux I__1516 (
            .O(N__15387),
            .I(N__15381));
    Odrv4 I__1515 (
            .O(N__15384),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_4 ));
    Odrv4 I__1514 (
            .O(N__15381),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_4 ));
    CascadeMux I__1513 (
            .O(N__15376),
            .I(\this_ppu.m62_0_a2_0_o2_0_cascade_ ));
    InMux I__1512 (
            .O(N__15373),
            .I(N__15370));
    LocalMux I__1511 (
            .O(N__15370),
            .I(M_this_oam_ram_write_data_23));
    InMux I__1510 (
            .O(N__15367),
            .I(N__15364));
    LocalMux I__1509 (
            .O(N__15364),
            .I(M_this_oam_ram_write_data_20));
    InMux I__1508 (
            .O(N__15361),
            .I(N__15358));
    LocalMux I__1507 (
            .O(N__15358),
            .I(M_this_oam_ram_write_data_19));
    InMux I__1506 (
            .O(N__15355),
            .I(N__15352));
    LocalMux I__1505 (
            .O(N__15352),
            .I(M_this_oam_ram_write_data_17));
    IoInMux I__1504 (
            .O(N__15349),
            .I(N__15346));
    LocalMux I__1503 (
            .O(N__15346),
            .I(N__15343));
    IoSpan4Mux I__1502 (
            .O(N__15343),
            .I(N__15340));
    Span4Mux_s3_h I__1501 (
            .O(N__15340),
            .I(N__15337));
    Span4Mux_h I__1500 (
            .O(N__15337),
            .I(N__15334));
    Odrv4 I__1499 (
            .O(N__15334),
            .I(rgb_c_1));
    InMux I__1498 (
            .O(N__15331),
            .I(N__15328));
    LocalMux I__1497 (
            .O(N__15328),
            .I(N__15325));
    Span4Mux_h I__1496 (
            .O(N__15325),
            .I(N__15321));
    InMux I__1495 (
            .O(N__15324),
            .I(N__15318));
    Span4Mux_v I__1494 (
            .O(N__15321),
            .I(N__15315));
    LocalMux I__1493 (
            .O(N__15318),
            .I(N__15312));
    Span4Mux_v I__1492 (
            .O(N__15315),
            .I(N__15309));
    Span4Mux_h I__1491 (
            .O(N__15312),
            .I(N__15306));
    Odrv4 I__1490 (
            .O(N__15309),
            .I(M_this_oam_ram_read_data_0));
    Odrv4 I__1489 (
            .O(N__15306),
            .I(M_this_oam_ram_read_data_0));
    InMux I__1488 (
            .O(N__15301),
            .I(N__15298));
    LocalMux I__1487 (
            .O(N__15298),
            .I(N__15295));
    Span4Mux_h I__1486 (
            .O(N__15295),
            .I(N__15292));
    Odrv4 I__1485 (
            .O(N__15292),
            .I(\this_ppu.oam_cache.N_586_0 ));
    InMux I__1484 (
            .O(N__15289),
            .I(N__15286));
    LocalMux I__1483 (
            .O(N__15286),
            .I(N__15283));
    Span4Mux_h I__1482 (
            .O(N__15283),
            .I(N__15280));
    Odrv4 I__1481 (
            .O(N__15280),
            .I(\this_ppu.oam_cache.mem_10 ));
    InMux I__1480 (
            .O(N__15277),
            .I(N__15274));
    LocalMux I__1479 (
            .O(N__15274),
            .I(\this_ppu.N_844_0 ));
    InMux I__1478 (
            .O(N__15271),
            .I(N__15268));
    LocalMux I__1477 (
            .O(N__15268),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_10 ));
    InMux I__1476 (
            .O(N__15265),
            .I(un1_M_this_warmup_d_cry_20));
    InMux I__1475 (
            .O(N__15262),
            .I(N__15259));
    LocalMux I__1474 (
            .O(N__15259),
            .I(M_this_warmup_qZ0Z_22));
    InMux I__1473 (
            .O(N__15256),
            .I(un1_M_this_warmup_d_cry_21));
    InMux I__1472 (
            .O(N__15253),
            .I(N__15250));
    LocalMux I__1471 (
            .O(N__15250),
            .I(M_this_warmup_qZ0Z_23));
    InMux I__1470 (
            .O(N__15247),
            .I(un1_M_this_warmup_d_cry_22));
    InMux I__1469 (
            .O(N__15244),
            .I(N__15241));
    LocalMux I__1468 (
            .O(N__15241),
            .I(M_this_warmup_qZ0Z_24));
    InMux I__1467 (
            .O(N__15238),
            .I(un1_M_this_warmup_d_cry_23));
    InMux I__1466 (
            .O(N__15235),
            .I(N__15232));
    LocalMux I__1465 (
            .O(N__15232),
            .I(M_this_warmup_qZ0Z_25));
    InMux I__1464 (
            .O(N__15229),
            .I(bfn_9_25_0_));
    InMux I__1463 (
            .O(N__15226),
            .I(N__15223));
    LocalMux I__1462 (
            .O(N__15223),
            .I(M_this_warmup_qZ0Z_26));
    InMux I__1461 (
            .O(N__15220),
            .I(un1_M_this_warmup_d_cry_25));
    InMux I__1460 (
            .O(N__15217),
            .I(un1_M_this_warmup_d_cry_26));
    InMux I__1459 (
            .O(N__15214),
            .I(N__15208));
    InMux I__1458 (
            .O(N__15213),
            .I(N__15208));
    LocalMux I__1457 (
            .O(N__15208),
            .I(M_this_warmup_qZ0Z_27));
    InMux I__1456 (
            .O(N__15205),
            .I(N__15202));
    LocalMux I__1455 (
            .O(N__15202),
            .I(M_this_oam_ram_write_data_18));
    InMux I__1454 (
            .O(N__15199),
            .I(N__15196));
    LocalMux I__1453 (
            .O(N__15196),
            .I(M_this_warmup_qZ0Z_13));
    InMux I__1452 (
            .O(N__15193),
            .I(un1_M_this_warmup_d_cry_12));
    InMux I__1451 (
            .O(N__15190),
            .I(N__15187));
    LocalMux I__1450 (
            .O(N__15187),
            .I(M_this_warmup_qZ0Z_14));
    InMux I__1449 (
            .O(N__15184),
            .I(un1_M_this_warmup_d_cry_13));
    InMux I__1448 (
            .O(N__15181),
            .I(N__15178));
    LocalMux I__1447 (
            .O(N__15178),
            .I(M_this_warmup_qZ0Z_15));
    InMux I__1446 (
            .O(N__15175),
            .I(un1_M_this_warmup_d_cry_14));
    InMux I__1445 (
            .O(N__15172),
            .I(N__15169));
    LocalMux I__1444 (
            .O(N__15169),
            .I(M_this_warmup_qZ0Z_16));
    InMux I__1443 (
            .O(N__15166),
            .I(un1_M_this_warmup_d_cry_15));
    InMux I__1442 (
            .O(N__15163),
            .I(N__15160));
    LocalMux I__1441 (
            .O(N__15160),
            .I(M_this_warmup_qZ0Z_17));
    InMux I__1440 (
            .O(N__15157),
            .I(bfn_9_24_0_));
    InMux I__1439 (
            .O(N__15154),
            .I(N__15151));
    LocalMux I__1438 (
            .O(N__15151),
            .I(M_this_warmup_qZ0Z_18));
    InMux I__1437 (
            .O(N__15148),
            .I(un1_M_this_warmup_d_cry_17));
    InMux I__1436 (
            .O(N__15145),
            .I(N__15142));
    LocalMux I__1435 (
            .O(N__15142),
            .I(M_this_warmup_qZ0Z_19));
    InMux I__1434 (
            .O(N__15139),
            .I(un1_M_this_warmup_d_cry_18));
    InMux I__1433 (
            .O(N__15136),
            .I(N__15133));
    LocalMux I__1432 (
            .O(N__15133),
            .I(M_this_warmup_qZ0Z_20));
    InMux I__1431 (
            .O(N__15130),
            .I(un1_M_this_warmup_d_cry_19));
    InMux I__1430 (
            .O(N__15127),
            .I(N__15124));
    LocalMux I__1429 (
            .O(N__15124),
            .I(M_this_warmup_qZ0Z_21));
    InMux I__1428 (
            .O(N__15121),
            .I(N__15118));
    LocalMux I__1427 (
            .O(N__15118),
            .I(M_this_warmup_qZ0Z_5));
    InMux I__1426 (
            .O(N__15115),
            .I(un1_M_this_warmup_d_cry_4));
    InMux I__1425 (
            .O(N__15112),
            .I(N__15109));
    LocalMux I__1424 (
            .O(N__15109),
            .I(M_this_warmup_qZ0Z_6));
    InMux I__1423 (
            .O(N__15106),
            .I(un1_M_this_warmup_d_cry_5));
    InMux I__1422 (
            .O(N__15103),
            .I(N__15100));
    LocalMux I__1421 (
            .O(N__15100),
            .I(M_this_warmup_qZ0Z_7));
    InMux I__1420 (
            .O(N__15097),
            .I(un1_M_this_warmup_d_cry_6));
    InMux I__1419 (
            .O(N__15094),
            .I(N__15091));
    LocalMux I__1418 (
            .O(N__15091),
            .I(M_this_warmup_qZ0Z_8));
    InMux I__1417 (
            .O(N__15088),
            .I(un1_M_this_warmup_d_cry_7));
    InMux I__1416 (
            .O(N__15085),
            .I(N__15082));
    LocalMux I__1415 (
            .O(N__15082),
            .I(M_this_warmup_qZ0Z_9));
    InMux I__1414 (
            .O(N__15079),
            .I(bfn_9_23_0_));
    InMux I__1413 (
            .O(N__15076),
            .I(N__15073));
    LocalMux I__1412 (
            .O(N__15073),
            .I(M_this_warmup_qZ0Z_10));
    InMux I__1411 (
            .O(N__15070),
            .I(un1_M_this_warmup_d_cry_9));
    InMux I__1410 (
            .O(N__15067),
            .I(N__15064));
    LocalMux I__1409 (
            .O(N__15064),
            .I(M_this_warmup_qZ0Z_11));
    InMux I__1408 (
            .O(N__15061),
            .I(un1_M_this_warmup_d_cry_10));
    InMux I__1407 (
            .O(N__15058),
            .I(N__15055));
    LocalMux I__1406 (
            .O(N__15055),
            .I(M_this_warmup_qZ0Z_12));
    InMux I__1405 (
            .O(N__15052),
            .I(un1_M_this_warmup_d_cry_11));
    InMux I__1404 (
            .O(N__15049),
            .I(N__15046));
    LocalMux I__1403 (
            .O(N__15046),
            .I(N__15043));
    Span4Mux_h I__1402 (
            .O(N__15043),
            .I(N__15040));
    Odrv4 I__1401 (
            .O(N__15040),
            .I(\this_ppu.oam_cache.mem_2 ));
    InMux I__1400 (
            .O(N__15037),
            .I(N__15034));
    LocalMux I__1399 (
            .O(N__15034),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_21 ));
    InMux I__1398 (
            .O(N__15031),
            .I(N__15028));
    LocalMux I__1397 (
            .O(N__15028),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_22 ));
    InMux I__1396 (
            .O(N__15025),
            .I(N__15022));
    LocalMux I__1395 (
            .O(N__15022),
            .I(N__15018));
    InMux I__1394 (
            .O(N__15021),
            .I(N__15015));
    Span4Mux_v I__1393 (
            .O(N__15018),
            .I(N__15010));
    LocalMux I__1392 (
            .O(N__15015),
            .I(N__15010));
    Odrv4 I__1391 (
            .O(N__15010),
            .I(M_this_oam_ram_read_data_3));
    InMux I__1390 (
            .O(N__15007),
            .I(N__15003));
    CascadeMux I__1389 (
            .O(N__15006),
            .I(N__15000));
    LocalMux I__1388 (
            .O(N__15003),
            .I(N__14997));
    InMux I__1387 (
            .O(N__15000),
            .I(N__14994));
    Span4Mux_v I__1386 (
            .O(N__14997),
            .I(N__14989));
    LocalMux I__1385 (
            .O(N__14994),
            .I(N__14989));
    Odrv4 I__1384 (
            .O(N__14989),
            .I(M_this_oam_ram_read_data_6));
    InMux I__1383 (
            .O(N__14986),
            .I(N__14983));
    LocalMux I__1382 (
            .O(N__14983),
            .I(N__14980));
    Span4Mux_v I__1381 (
            .O(N__14980),
            .I(N__14977));
    Odrv4 I__1380 (
            .O(N__14977),
            .I(M_this_oam_ram_read_data_25));
    InMux I__1379 (
            .O(N__14974),
            .I(N__14971));
    LocalMux I__1378 (
            .O(N__14971),
            .I(N__14968));
    Span4Mux_h I__1377 (
            .O(N__14968),
            .I(N__14965));
    Odrv4 I__1376 (
            .O(N__14965),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_25 ));
    InMux I__1375 (
            .O(N__14962),
            .I(N__14958));
    InMux I__1374 (
            .O(N__14961),
            .I(N__14955));
    LocalMux I__1373 (
            .O(N__14958),
            .I(N__14952));
    LocalMux I__1372 (
            .O(N__14955),
            .I(M_this_warmup_qZ0Z_1));
    Odrv4 I__1371 (
            .O(N__14952),
            .I(M_this_warmup_qZ0Z_1));
    CascadeMux I__1370 (
            .O(N__14947),
            .I(N__14942));
    InMux I__1369 (
            .O(N__14946),
            .I(N__14937));
    InMux I__1368 (
            .O(N__14945),
            .I(N__14937));
    InMux I__1367 (
            .O(N__14942),
            .I(N__14934));
    LocalMux I__1366 (
            .O(N__14937),
            .I(N__14929));
    LocalMux I__1365 (
            .O(N__14934),
            .I(N__14929));
    Odrv4 I__1364 (
            .O(N__14929),
            .I(M_this_warmup_qZ0Z_0));
    InMux I__1363 (
            .O(N__14926),
            .I(N__14923));
    LocalMux I__1362 (
            .O(N__14923),
            .I(M_this_warmup_qZ0Z_2));
    InMux I__1361 (
            .O(N__14920),
            .I(un1_M_this_warmup_d_cry_1));
    InMux I__1360 (
            .O(N__14917),
            .I(N__14914));
    LocalMux I__1359 (
            .O(N__14914),
            .I(M_this_warmup_qZ0Z_3));
    InMux I__1358 (
            .O(N__14911),
            .I(un1_M_this_warmup_d_cry_2));
    InMux I__1357 (
            .O(N__14908),
            .I(N__14905));
    LocalMux I__1356 (
            .O(N__14905),
            .I(M_this_warmup_qZ0Z_4));
    InMux I__1355 (
            .O(N__14902),
            .I(un1_M_this_warmup_d_cry_3));
    CascadeMux I__1354 (
            .O(N__14899),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_cascade_ ));
    InMux I__1353 (
            .O(N__14896),
            .I(N__14891));
    InMux I__1352 (
            .O(N__14895),
            .I(N__14886));
    InMux I__1351 (
            .O(N__14894),
            .I(N__14886));
    LocalMux I__1350 (
            .O(N__14891),
            .I(N__14883));
    LocalMux I__1349 (
            .O(N__14886),
            .I(\this_ppu.N_841_0 ));
    Odrv4 I__1348 (
            .O(N__14883),
            .I(\this_ppu.N_841_0 ));
    CascadeMux I__1347 (
            .O(N__14878),
            .I(\this_ppu.N_841_0_cascade_ ));
    CascadeMux I__1346 (
            .O(N__14875),
            .I(N__14872));
    CascadeBuf I__1345 (
            .O(N__14872),
            .I(N__14869));
    CascadeMux I__1344 (
            .O(N__14869),
            .I(N__14866));
    InMux I__1343 (
            .O(N__14866),
            .I(N__14863));
    LocalMux I__1342 (
            .O(N__14863),
            .I(\this_ppu.N_669_0 ));
    CascadeMux I__1341 (
            .O(N__14860),
            .I(\this_ppu.m18_i_o2_1_cascade_ ));
    InMux I__1340 (
            .O(N__14857),
            .I(N__14851));
    InMux I__1339 (
            .O(N__14856),
            .I(N__14844));
    InMux I__1338 (
            .O(N__14855),
            .I(N__14844));
    InMux I__1337 (
            .O(N__14854),
            .I(N__14844));
    LocalMux I__1336 (
            .O(N__14851),
            .I(\this_ppu.N_426_0 ));
    LocalMux I__1335 (
            .O(N__14844),
            .I(\this_ppu.N_426_0 ));
    CascadeMux I__1334 (
            .O(N__14839),
            .I(N__14836));
    InMux I__1333 (
            .O(N__14836),
            .I(N__14833));
    LocalMux I__1332 (
            .O(N__14833),
            .I(M_this_vga_signals_address_2));
    InMux I__1331 (
            .O(N__14830),
            .I(N__14827));
    LocalMux I__1330 (
            .O(N__14827),
            .I(\this_ppu.oam_cache.mem_4 ));
    CascadeMux I__1329 (
            .O(N__14824),
            .I(N__14821));
    CascadeBuf I__1328 (
            .O(N__14821),
            .I(N__14818));
    CascadeMux I__1327 (
            .O(N__14818),
            .I(N__14815));
    InMux I__1326 (
            .O(N__14815),
            .I(N__14812));
    LocalMux I__1325 (
            .O(N__14812),
            .I(\this_ppu.N_985_0 ));
    CascadeMux I__1324 (
            .O(N__14809),
            .I(N__14806));
    CascadeBuf I__1323 (
            .O(N__14806),
            .I(N__14803));
    CascadeMux I__1322 (
            .O(N__14803),
            .I(N__14800));
    InMux I__1321 (
            .O(N__14800),
            .I(N__14797));
    LocalMux I__1320 (
            .O(N__14797),
            .I(\this_ppu.N_671_0 ));
    CascadeMux I__1319 (
            .O(N__14794),
            .I(\this_ppu.N_426_0_cascade_ ));
    CascadeMux I__1318 (
            .O(N__14791),
            .I(\this_ppu.un1_M_oam_curr_q_1_c2_cascade_ ));
    CascadeMux I__1317 (
            .O(N__14788),
            .I(N__14785));
    CascadeBuf I__1316 (
            .O(N__14785),
            .I(N__14782));
    CascadeMux I__1315 (
            .O(N__14782),
            .I(N__14779));
    InMux I__1314 (
            .O(N__14779),
            .I(N__14776));
    LocalMux I__1313 (
            .O(N__14776),
            .I(\this_ppu.N_986_0 ));
    CascadeMux I__1312 (
            .O(N__14773),
            .I(\this_ppu.un1_M_oam_curr_q_1_c4_cascade_ ));
    IoInMux I__1311 (
            .O(N__14770),
            .I(N__14767));
    LocalMux I__1310 (
            .O(N__14767),
            .I(N__14764));
    IoSpan4Mux I__1309 (
            .O(N__14764),
            .I(N__14761));
    Span4Mux_s2_h I__1308 (
            .O(N__14761),
            .I(N__14758));
    Sp12to4 I__1307 (
            .O(N__14758),
            .I(N__14755));
    Span12Mux_s8_h I__1306 (
            .O(N__14755),
            .I(N__14752));
    Odrv12 I__1305 (
            .O(N__14752),
            .I(rgb_c_0));
    InMux I__1304 (
            .O(N__14749),
            .I(N__14746));
    LocalMux I__1303 (
            .O(N__14746),
            .I(N__14743));
    Span4Mux_v I__1302 (
            .O(N__14743),
            .I(N__14740));
    Odrv4 I__1301 (
            .O(N__14740),
            .I(M_this_oam_ram_read_data_15));
    InMux I__1300 (
            .O(N__14737),
            .I(N__14734));
    LocalMux I__1299 (
            .O(N__14734),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_15 ));
    InMux I__1298 (
            .O(N__14731),
            .I(N__14728));
    LocalMux I__1297 (
            .O(N__14728),
            .I(\this_ppu.oam_cache.N_577_0 ));
    InMux I__1296 (
            .O(N__14725),
            .I(N__14722));
    LocalMux I__1295 (
            .O(N__14722),
            .I(\this_ppu.oam_cache.N_567_0 ));
    InMux I__1294 (
            .O(N__14719),
            .I(N__14716));
    LocalMux I__1293 (
            .O(N__14716),
            .I(N__14713));
    Span4Mux_v I__1292 (
            .O(N__14713),
            .I(N__14710));
    Odrv4 I__1291 (
            .O(N__14710),
            .I(M_this_oam_ram_read_data_8));
    InMux I__1290 (
            .O(N__14707),
            .I(N__14704));
    LocalMux I__1289 (
            .O(N__14704),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_8 ));
    InMux I__1288 (
            .O(N__14701),
            .I(N__14698));
    LocalMux I__1287 (
            .O(N__14698),
            .I(N__14695));
    Span12Mux_h I__1286 (
            .O(N__14695),
            .I(N__14692));
    Odrv12 I__1285 (
            .O(N__14692),
            .I(M_this_oam_ram_read_data_9));
    InMux I__1284 (
            .O(N__14689),
            .I(N__14686));
    LocalMux I__1283 (
            .O(N__14686),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_9 ));
    InMux I__1282 (
            .O(N__14683),
            .I(N__14680));
    LocalMux I__1281 (
            .O(N__14680),
            .I(N__14677));
    Span4Mux_h I__1280 (
            .O(N__14677),
            .I(N__14674));
    Span4Mux_v I__1279 (
            .O(N__14674),
            .I(N__14671));
    Odrv4 I__1278 (
            .O(N__14671),
            .I(M_this_oam_ram_read_data_10));
    InMux I__1277 (
            .O(N__14668),
            .I(N__14665));
    LocalMux I__1276 (
            .O(N__14665),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_10 ));
    InMux I__1275 (
            .O(N__14662),
            .I(N__14659));
    LocalMux I__1274 (
            .O(N__14659),
            .I(N__14656));
    Span4Mux_h I__1273 (
            .O(N__14656),
            .I(N__14653));
    Odrv4 I__1272 (
            .O(N__14653),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_16 ));
    InMux I__1271 (
            .O(N__14650),
            .I(N__14647));
    LocalMux I__1270 (
            .O(N__14647),
            .I(\this_ppu.oam_cache.mem_18 ));
    InMux I__1269 (
            .O(N__14644),
            .I(N__14641));
    LocalMux I__1268 (
            .O(N__14641),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_18 ));
    InMux I__1267 (
            .O(N__14638),
            .I(N__14635));
    LocalMux I__1266 (
            .O(N__14635),
            .I(N__14632));
    Odrv12 I__1265 (
            .O(N__14632),
            .I(port_clk_c));
    InMux I__1264 (
            .O(N__14629),
            .I(N__14626));
    LocalMux I__1263 (
            .O(N__14626),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    InMux I__1262 (
            .O(N__14623),
            .I(N__14620));
    LocalMux I__1261 (
            .O(N__14620),
            .I(N__14617));
    Odrv4 I__1260 (
            .O(N__14617),
            .I(M_this_oam_ram_read_data_12));
    InMux I__1259 (
            .O(N__14614),
            .I(N__14611));
    LocalMux I__1258 (
            .O(N__14611),
            .I(N__14608));
    Span4Mux_h I__1257 (
            .O(N__14608),
            .I(N__14605));
    Odrv4 I__1256 (
            .O(N__14605),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_12 ));
    InMux I__1255 (
            .O(N__14602),
            .I(N__14599));
    LocalMux I__1254 (
            .O(N__14599),
            .I(N__14596));
    Span4Mux_h I__1253 (
            .O(N__14596),
            .I(N__14593));
    Odrv4 I__1252 (
            .O(N__14593),
            .I(\this_ppu.oam_cache.N_579_0 ));
    InMux I__1251 (
            .O(N__14590),
            .I(N__14587));
    LocalMux I__1250 (
            .O(N__14587),
            .I(N__14584));
    Span4Mux_h I__1249 (
            .O(N__14584),
            .I(N__14581));
    Odrv4 I__1248 (
            .O(N__14581),
            .I(M_this_oam_ram_read_data_26));
    InMux I__1247 (
            .O(N__14578),
            .I(N__14575));
    LocalMux I__1246 (
            .O(N__14575),
            .I(N__14572));
    Odrv4 I__1245 (
            .O(N__14572),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_26 ));
    IoInMux I__1244 (
            .O(N__14569),
            .I(N__14566));
    LocalMux I__1243 (
            .O(N__14566),
            .I(N__14563));
    IoSpan4Mux I__1242 (
            .O(N__14563),
            .I(N__14560));
    Span4Mux_s1_v I__1241 (
            .O(N__14560),
            .I(N__14557));
    Span4Mux_v I__1240 (
            .O(N__14557),
            .I(N__14554));
    Odrv4 I__1239 (
            .O(N__14554),
            .I(N_84));
    IoInMux I__1238 (
            .O(N__14551),
            .I(N__14548));
    LocalMux I__1237 (
            .O(N__14548),
            .I(N__14545));
    Span4Mux_s2_h I__1236 (
            .O(N__14545),
            .I(N__14542));
    Span4Mux_h I__1235 (
            .O(N__14542),
            .I(N__14539));
    Span4Mux_v I__1234 (
            .O(N__14539),
            .I(N__14536));
    Span4Mux_v I__1233 (
            .O(N__14536),
            .I(N__14533));
    Odrv4 I__1232 (
            .O(N__14533),
            .I(rgb_c_5));
    InMux I__1231 (
            .O(N__14530),
            .I(N__14527));
    LocalMux I__1230 (
            .O(N__14527),
            .I(\this_ppu.oam_cache.N_561_0 ));
    InMux I__1229 (
            .O(N__14524),
            .I(N__14521));
    LocalMux I__1228 (
            .O(N__14521),
            .I(N__14518));
    Odrv4 I__1227 (
            .O(N__14518),
            .I(\this_ppu.oam_cache.mem_17 ));
    InMux I__1226 (
            .O(N__14515),
            .I(N__14512));
    LocalMux I__1225 (
            .O(N__14512),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_17 ));
    CascadeMux I__1224 (
            .O(N__14509),
            .I(N__14506));
    InMux I__1223 (
            .O(N__14506),
            .I(N__14503));
    LocalMux I__1222 (
            .O(N__14503),
            .I(\this_ppu.M_oam_cache_read_data_i_16 ));
    InMux I__1221 (
            .O(N__14500),
            .I(N__14497));
    LocalMux I__1220 (
            .O(N__14497),
            .I(\this_ppu.M_oam_cache_read_data_i_17 ));
    CascadeMux I__1219 (
            .O(N__14494),
            .I(N__14491));
    InMux I__1218 (
            .O(N__14491),
            .I(N__14487));
    CascadeMux I__1217 (
            .O(N__14490),
            .I(N__14484));
    LocalMux I__1216 (
            .O(N__14487),
            .I(N__14477));
    InMux I__1215 (
            .O(N__14484),
            .I(N__14474));
    CascadeMux I__1214 (
            .O(N__14483),
            .I(N__14471));
    CascadeMux I__1213 (
            .O(N__14482),
            .I(N__14467));
    CascadeMux I__1212 (
            .O(N__14481),
            .I(N__14463));
    CascadeMux I__1211 (
            .O(N__14480),
            .I(N__14460));
    Span4Mux_v I__1210 (
            .O(N__14477),
            .I(N__14453));
    LocalMux I__1209 (
            .O(N__14474),
            .I(N__14453));
    InMux I__1208 (
            .O(N__14471),
            .I(N__14450));
    CascadeMux I__1207 (
            .O(N__14470),
            .I(N__14447));
    InMux I__1206 (
            .O(N__14467),
            .I(N__14443));
    CascadeMux I__1205 (
            .O(N__14466),
            .I(N__14440));
    InMux I__1204 (
            .O(N__14463),
            .I(N__14437));
    InMux I__1203 (
            .O(N__14460),
            .I(N__14434));
    CascadeMux I__1202 (
            .O(N__14459),
            .I(N__14431));
    CascadeMux I__1201 (
            .O(N__14458),
            .I(N__14428));
    Span4Mux_h I__1200 (
            .O(N__14453),
            .I(N__14423));
    LocalMux I__1199 (
            .O(N__14450),
            .I(N__14423));
    InMux I__1198 (
            .O(N__14447),
            .I(N__14420));
    CascadeMux I__1197 (
            .O(N__14446),
            .I(N__14417));
    LocalMux I__1196 (
            .O(N__14443),
            .I(N__14413));
    InMux I__1195 (
            .O(N__14440),
            .I(N__14410));
    LocalMux I__1194 (
            .O(N__14437),
            .I(N__14404));
    LocalMux I__1193 (
            .O(N__14434),
            .I(N__14404));
    InMux I__1192 (
            .O(N__14431),
            .I(N__14401));
    InMux I__1191 (
            .O(N__14428),
            .I(N__14398));
    Span4Mux_v I__1190 (
            .O(N__14423),
            .I(N__14393));
    LocalMux I__1189 (
            .O(N__14420),
            .I(N__14393));
    InMux I__1188 (
            .O(N__14417),
            .I(N__14390));
    CascadeMux I__1187 (
            .O(N__14416),
            .I(N__14387));
    Span4Mux_s2_v I__1186 (
            .O(N__14413),
            .I(N__14380));
    LocalMux I__1185 (
            .O(N__14410),
            .I(N__14380));
    CascadeMux I__1184 (
            .O(N__14409),
            .I(N__14377));
    Span4Mux_v I__1183 (
            .O(N__14404),
            .I(N__14370));
    LocalMux I__1182 (
            .O(N__14401),
            .I(N__14370));
    LocalMux I__1181 (
            .O(N__14398),
            .I(N__14370));
    Span4Mux_h I__1180 (
            .O(N__14393),
            .I(N__14365));
    LocalMux I__1179 (
            .O(N__14390),
            .I(N__14365));
    InMux I__1178 (
            .O(N__14387),
            .I(N__14361));
    CascadeMux I__1177 (
            .O(N__14386),
            .I(N__14358));
    CascadeMux I__1176 (
            .O(N__14385),
            .I(N__14355));
    Span4Mux_v I__1175 (
            .O(N__14380),
            .I(N__14352));
    InMux I__1174 (
            .O(N__14377),
            .I(N__14349));
    Span4Mux_v I__1173 (
            .O(N__14370),
            .I(N__14344));
    Span4Mux_v I__1172 (
            .O(N__14365),
            .I(N__14344));
    CascadeMux I__1171 (
            .O(N__14364),
            .I(N__14341));
    LocalMux I__1170 (
            .O(N__14361),
            .I(N__14338));
    InMux I__1169 (
            .O(N__14358),
            .I(N__14335));
    InMux I__1168 (
            .O(N__14355),
            .I(N__14332));
    Sp12to4 I__1167 (
            .O(N__14352),
            .I(N__14327));
    LocalMux I__1166 (
            .O(N__14349),
            .I(N__14327));
    Sp12to4 I__1165 (
            .O(N__14344),
            .I(N__14324));
    InMux I__1164 (
            .O(N__14341),
            .I(N__14321));
    Span4Mux_s3_v I__1163 (
            .O(N__14338),
            .I(N__14314));
    LocalMux I__1162 (
            .O(N__14335),
            .I(N__14314));
    LocalMux I__1161 (
            .O(N__14332),
            .I(N__14314));
    Span12Mux_h I__1160 (
            .O(N__14327),
            .I(N__14311));
    Span12Mux_s6_h I__1159 (
            .O(N__14324),
            .I(N__14306));
    LocalMux I__1158 (
            .O(N__14321),
            .I(N__14306));
    Span4Mux_v I__1157 (
            .O(N__14314),
            .I(N__14303));
    Span12Mux_v I__1156 (
            .O(N__14311),
            .I(N__14298));
    Span12Mux_h I__1155 (
            .O(N__14306),
            .I(N__14298));
    Span4Mux_v I__1154 (
            .O(N__14303),
            .I(N__14295));
    Odrv12 I__1153 (
            .O(N__14298),
            .I(M_this_ppu_spr_addr_4));
    Odrv4 I__1152 (
            .O(N__14295),
            .I(M_this_ppu_spr_addr_4));
    InMux I__1151 (
            .O(N__14290),
            .I(\this_ppu.offset_y_cry_0 ));
    InMux I__1150 (
            .O(N__14287),
            .I(\this_ppu.offset_y_cry_1 ));
    CascadeMux I__1149 (
            .O(N__14284),
            .I(N__14277));
    CascadeMux I__1148 (
            .O(N__14283),
            .I(N__14273));
    CascadeMux I__1147 (
            .O(N__14282),
            .I(N__14270));
    CascadeMux I__1146 (
            .O(N__14281),
            .I(N__14259));
    CascadeMux I__1145 (
            .O(N__14280),
            .I(N__14254));
    InMux I__1144 (
            .O(N__14277),
            .I(N__14251));
    CascadeMux I__1143 (
            .O(N__14276),
            .I(N__14248));
    InMux I__1142 (
            .O(N__14273),
            .I(N__14245));
    InMux I__1141 (
            .O(N__14270),
            .I(N__14242));
    CascadeMux I__1140 (
            .O(N__14269),
            .I(N__14239));
    CascadeMux I__1139 (
            .O(N__14268),
            .I(N__14236));
    CascadeMux I__1138 (
            .O(N__14267),
            .I(N__14233));
    CascadeMux I__1137 (
            .O(N__14266),
            .I(N__14230));
    CascadeMux I__1136 (
            .O(N__14265),
            .I(N__14227));
    CascadeMux I__1135 (
            .O(N__14264),
            .I(N__14224));
    CascadeMux I__1134 (
            .O(N__14263),
            .I(N__14221));
    CascadeMux I__1133 (
            .O(N__14262),
            .I(N__14218));
    InMux I__1132 (
            .O(N__14259),
            .I(N__14215));
    CascadeMux I__1131 (
            .O(N__14258),
            .I(N__14212));
    CascadeMux I__1130 (
            .O(N__14257),
            .I(N__14209));
    InMux I__1129 (
            .O(N__14254),
            .I(N__14206));
    LocalMux I__1128 (
            .O(N__14251),
            .I(N__14203));
    InMux I__1127 (
            .O(N__14248),
            .I(N__14200));
    LocalMux I__1126 (
            .O(N__14245),
            .I(N__14197));
    LocalMux I__1125 (
            .O(N__14242),
            .I(N__14194));
    InMux I__1124 (
            .O(N__14239),
            .I(N__14191));
    InMux I__1123 (
            .O(N__14236),
            .I(N__14188));
    InMux I__1122 (
            .O(N__14233),
            .I(N__14185));
    InMux I__1121 (
            .O(N__14230),
            .I(N__14182));
    InMux I__1120 (
            .O(N__14227),
            .I(N__14179));
    InMux I__1119 (
            .O(N__14224),
            .I(N__14176));
    InMux I__1118 (
            .O(N__14221),
            .I(N__14173));
    InMux I__1117 (
            .O(N__14218),
            .I(N__14170));
    LocalMux I__1116 (
            .O(N__14215),
            .I(N__14167));
    InMux I__1115 (
            .O(N__14212),
            .I(N__14164));
    InMux I__1114 (
            .O(N__14209),
            .I(N__14161));
    LocalMux I__1113 (
            .O(N__14206),
            .I(N__14158));
    Span12Mux_h I__1112 (
            .O(N__14203),
            .I(N__14155));
    LocalMux I__1111 (
            .O(N__14200),
            .I(N__14152));
    Span12Mux_s6_v I__1110 (
            .O(N__14197),
            .I(N__14147));
    Span12Mux_s7_h I__1109 (
            .O(N__14194),
            .I(N__14147));
    LocalMux I__1108 (
            .O(N__14191),
            .I(N__14140));
    LocalMux I__1107 (
            .O(N__14188),
            .I(N__14140));
    LocalMux I__1106 (
            .O(N__14185),
            .I(N__14140));
    LocalMux I__1105 (
            .O(N__14182),
            .I(N__14131));
    LocalMux I__1104 (
            .O(N__14179),
            .I(N__14131));
    LocalMux I__1103 (
            .O(N__14176),
            .I(N__14131));
    LocalMux I__1102 (
            .O(N__14173),
            .I(N__14131));
    LocalMux I__1101 (
            .O(N__14170),
            .I(N__14128));
    Span4Mux_s2_v I__1100 (
            .O(N__14167),
            .I(N__14121));
    LocalMux I__1099 (
            .O(N__14164),
            .I(N__14121));
    LocalMux I__1098 (
            .O(N__14161),
            .I(N__14121));
    Span12Mux_h I__1097 (
            .O(N__14158),
            .I(N__14118));
    Span12Mux_h I__1096 (
            .O(N__14155),
            .I(N__14115));
    Span12Mux_h I__1095 (
            .O(N__14152),
            .I(N__14112));
    Span12Mux_h I__1094 (
            .O(N__14147),
            .I(N__14109));
    Span12Mux_v I__1093 (
            .O(N__14140),
            .I(N__14102));
    Span12Mux_v I__1092 (
            .O(N__14131),
            .I(N__14102));
    Span12Mux_s7_h I__1091 (
            .O(N__14128),
            .I(N__14102));
    Span4Mux_v I__1090 (
            .O(N__14121),
            .I(N__14099));
    Span12Mux_h I__1089 (
            .O(N__14118),
            .I(N__14096));
    Span12Mux_v I__1088 (
            .O(N__14115),
            .I(N__14091));
    Span12Mux_h I__1087 (
            .O(N__14112),
            .I(N__14091));
    Span12Mux_v I__1086 (
            .O(N__14109),
            .I(N__14086));
    Span12Mux_h I__1085 (
            .O(N__14102),
            .I(N__14086));
    Span4Mux_v I__1084 (
            .O(N__14099),
            .I(N__14083));
    Odrv12 I__1083 (
            .O(N__14096),
            .I(M_this_ppu_spr_addr_5));
    Odrv12 I__1082 (
            .O(N__14091),
            .I(M_this_ppu_spr_addr_5));
    Odrv12 I__1081 (
            .O(N__14086),
            .I(M_this_ppu_spr_addr_5));
    Odrv4 I__1080 (
            .O(N__14083),
            .I(M_this_ppu_spr_addr_5));
    InMux I__1079 (
            .O(N__14074),
            .I(N__14071));
    LocalMux I__1078 (
            .O(N__14071),
            .I(\this_ppu.oam_cache.mem_16 ));
    IoInMux I__1077 (
            .O(N__14068),
            .I(N__14065));
    LocalMux I__1076 (
            .O(N__14065),
            .I(\this_vga_signals.N_1307_0 ));
    IoInMux I__1075 (
            .O(N__14062),
            .I(N__14059));
    LocalMux I__1074 (
            .O(N__14059),
            .I(N_428));
    IoInMux I__1073 (
            .O(N__14056),
            .I(N__14053));
    LocalMux I__1072 (
            .O(N__14053),
            .I(N__14050));
    Span12Mux_s1_v I__1071 (
            .O(N__14050),
            .I(N__14047));
    Odrv12 I__1070 (
            .O(N__14047),
            .I(N_842));
    IoInMux I__1069 (
            .O(N__14044),
            .I(N__14041));
    LocalMux I__1068 (
            .O(N__14041),
            .I(N__14038));
    IoSpan4Mux I__1067 (
            .O(N__14038),
            .I(N__14035));
    Span4Mux_s3_v I__1066 (
            .O(N__14035),
            .I(N__14032));
    Span4Mux_v I__1065 (
            .O(N__14032),
            .I(N__14029));
    Span4Mux_v I__1064 (
            .O(N__14029),
            .I(N__14026));
    Span4Mux_v I__1063 (
            .O(N__14026),
            .I(N__14023));
    Odrv4 I__1062 (
            .O(N__14023),
            .I(rgb_c_4));
    IoInMux I__1061 (
            .O(N__14020),
            .I(N__14017));
    LocalMux I__1060 (
            .O(N__14017),
            .I(N__14014));
    IoSpan4Mux I__1059 (
            .O(N__14014),
            .I(N__14011));
    IoSpan4Mux I__1058 (
            .O(N__14011),
            .I(N__14008));
    Span4Mux_s3_h I__1057 (
            .O(N__14008),
            .I(N__14005));
    Odrv4 I__1056 (
            .O(N__14005),
            .I(M_vcounter_q_esr_RNIQ82H7_9));
    InMux I__1055 (
            .O(N__14002),
            .I(N__13999));
    LocalMux I__1054 (
            .O(N__13999),
            .I(N__13996));
    Span4Mux_v I__1053 (
            .O(N__13996),
            .I(N__13993));
    Odrv4 I__1052 (
            .O(N__13993),
            .I(M_this_oam_ram_read_data_13));
    InMux I__1051 (
            .O(N__13990),
            .I(N__13987));
    LocalMux I__1050 (
            .O(N__13987),
            .I(N__13984));
    Span4Mux_h I__1049 (
            .O(N__13984),
            .I(N__13981));
    Odrv4 I__1048 (
            .O(N__13981),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_13 ));
    IoInMux I__1047 (
            .O(N__13978),
            .I(N__13975));
    LocalMux I__1046 (
            .O(N__13975),
            .I(N__13972));
    IoSpan4Mux I__1045 (
            .O(N__13972),
            .I(N__13969));
    Span4Mux_s3_h I__1044 (
            .O(N__13969),
            .I(N__13966));
    Odrv4 I__1043 (
            .O(N__13966),
            .I(rgb_c_2));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\this_ppu.un1_M_surface_y_d_cry_6 ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(un1_M_this_warmup_d_cry_8),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(un1_M_this_warmup_d_cry_16),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(un1_M_this_warmup_d_cry_24),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_24_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_23_0_));
    defparam IN_MUX_bfv_24_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_24_0_ (
            .carryinitin(un1_M_this_map_address_q_cry_7),
            .carryinitout(bfn_24_24_0_));
    defparam IN_MUX_bfv_26_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_26_21_0_));
    defparam IN_MUX_bfv_26_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_22_0_ (
            .carryinitin(un1_M_this_ext_address_q_cry_7),
            .carryinitout(bfn_26_22_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(M_this_data_count_q_cry_7),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_18_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_21_0_));
    defparam IN_MUX_bfv_18_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_22_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_18_22_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\this_ppu.offset_x_cry_6_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_22_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_14_0_));
    defparam IN_MUX_bfv_22_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_15_0_ (
            .carryinitin(un1_M_this_spr_address_q_cry_7),
            .carryinitout(bfn_22_15_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNIFLF77_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__14068),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_1307_0_g ));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNI01JU6_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__25600),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_1637_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNI6VB7_3  (
            .USERSIGNALTOGLOBALBUFFER(N__26116),
            .GLOBALBUFFEROUTPUT(M_this_reset_cond_out_g_0));
    ICE_GB \this_reset_cond.M_stage_q_RNI6VB7_0_3  (
            .USERSIGNALTOGLOBALBUFFER(N__21778),
            .GLOBALBUFFEROUTPUT(N_620_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFLF77_9_LC_1_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFLF77_9_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFLF77_9_LC_1_17_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIFLF77_9_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__27343),
            .in2(_gnd_net_),
            .in3(N__34225),
            .lcout(\this_vga_signals.N_1307_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.port_data_rw_i_i_LC_1_22_3 .C_ON=1'b0;
    defparam \this_ppu.port_data_rw_i_i_LC_1_22_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.port_data_rw_i_i_LC_1_22_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \this_ppu.port_data_rw_i_i_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(N__37755),
            .in2(_gnd_net_),
            .in3(N__32877),
            .lcout(N_428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_4_17_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_17_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_17_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA65T2_0_9_LC_5_25_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA65T2_0_9_LC_5_25_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA65T2_0_9_LC_5_25_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIA65T2_0_9_LC_5_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39506),
            .lcout(N_842),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_6_17_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_6_17_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_6_17_6  (
            .in0(N__17218),
            .in1(N__18526),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQ82H7_9_LC_6_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQ82H7_9_LC_6_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQ82H7_9_LC_6_18_6 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIQ82H7_9_LC_6_18_6  (
            .in0(N__39505),
            .in1(N__37735),
            .in2(_gnd_net_),
            .in3(N__37813),
            .lcout(M_vcounter_q_esr_RNIQ82H7_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_6_21_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_6_21_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_6_21_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_6_21_3  (
            .in0(N__24136),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14002),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_7_16_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_7_16_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_7_16_2  (
            .in0(N__18127),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17216),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_7_16_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_7_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__17217),
            .in2(_gnd_net_),
            .in3(N__20272),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_7_17_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_7_17_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(N__24081),
            .in2(_gnd_net_),
            .in3(N__15924),
            .lcout(\this_ppu.oam_cache.N_561_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_17_LC_7_18_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_17_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_17_LC_7_18_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_17_LC_7_18_6  (
            .in0(N__14524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42083),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNID8M7_17_LC_7_18_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNID8M7_17_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNID8M7_17_LC_7_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNID8M7_17_LC_7_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14515),
            .lcout(\this_ppu.M_oam_cache_read_data_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_y_cry_0_c_inv_LC_7_19_0 .C_ON=1'b1;
    defparam \this_ppu.offset_y_cry_0_c_inv_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_y_cry_0_c_inv_LC_7_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.offset_y_cry_0_c_inv_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__21586),
            .in2(N__14509),
            .in3(N__20151),
            .lcout(\this_ppu.M_oam_cache_read_data_i_16 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\this_ppu.offset_y_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_y_cry_0_c_RNIVBJT1_LC_7_19_1 .C_ON=1'b1;
    defparam \this_ppu.offset_y_cry_0_c_RNIVBJT1_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_y_cry_0_c_RNIVBJT1_LC_7_19_1 .LUT_INIT=16'b1110000110110100;
    LogicCell40 \this_ppu.offset_y_cry_0_c_RNIVBJT1_LC_7_19_1  (
            .in0(N__38187),
            .in1(N__14500),
            .in2(N__21541),
            .in3(N__14290),
            .lcout(M_this_ppu_spr_addr_4),
            .ltout(),
            .carryin(\this_ppu.offset_y_cry_0 ),
            .carryout(\this_ppu.offset_y_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI2GKT1_18_LC_7_19_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI2GKT1_18_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI2GKT1_18_LC_7_19_2 .LUT_INIT=16'b1101001011100001;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI2GKT1_18_LC_7_19_2  (
            .in0(N__14644),
            .in1(N__38188),
            .in2(N__21508),
            .in3(N__14287),
            .lcout(M_this_ppu_spr_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_16_LC_7_19_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_16_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_16_LC_7_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_16_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14074),
            .lcout(\this_ppu.M_oam_cache_read_data_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42097),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_18_LC_7_19_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_18_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_18_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_18_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14650),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42097),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_7_20_3 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_7_20_3 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_7_20_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_7_20_3  (
            .in0(N__14638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42102),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_7_20_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_7_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14629),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42102),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_7_21_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_7_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__14623),
            .in2(_gnd_net_),
            .in3(N__24137),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_7_21_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_7_21_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_7_21_6  (
            .in0(N__16860),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24139),
            .lcout(\this_ppu.oam_cache.N_579_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_7_21_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_7_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(N__14590),
            .in2(_gnd_net_),
            .in3(N__24138),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_warmup_q_0_LC_7_22_0.C_ON=1'b0;
    defparam M_this_warmup_q_0_LC_7_22_0.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_0_LC_7_22_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 M_this_warmup_q_0_LC_7_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14945),
            .lcout(M_this_warmup_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42116),
            .ce(),
            .sr(N__43129));
    defparam M_this_warmup_q_1_LC_7_22_5.C_ON=1'b0;
    defparam M_this_warmup_q_1_LC_7_22_5.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_1_LC_7_22_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 M_this_warmup_q_1_LC_7_22_5 (
            .in0(N__14946),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14961),
            .lcout(M_this_warmup_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42116),
            .ce(),
            .sr(N__43129));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_7_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_7_24_2 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_7_24_2  (
            .in0(N__17941),
            .in1(N__17806),
            .in2(_gnd_net_),
            .in3(N__17874),
            .lcout(N_84),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_9_15_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_9_15_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__17194),
            .in2(_gnd_net_),
            .in3(N__18148),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_3_LC_9_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_3_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_3_LC_9_17_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.M_state_q_3_LC_9_17_0  (
            .in0(N__23254),
            .in1(N__15277),
            .in2(_gnd_net_),
            .in3(N__17515),
            .lcout(\this_ppu.M_state_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42049),
            .ce(),
            .sr(N__43112));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_9_17_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_9_17_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__14749),
            .in2(_gnd_net_),
            .in3(N__24016),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_9_17_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_9_17_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_9_17_2  (
            .in0(N__24008),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15025),
            .lcout(\this_ppu.oam_cache.N_577_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_9_17_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_9_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__24011),
            .in2(_gnd_net_),
            .in3(N__15007),
            .lcout(\this_ppu.oam_cache.N_567_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_9_17_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_9_17_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_9_17_4  (
            .in0(N__24009),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14719),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_9_17_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_9_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__14701),
            .in2(_gnd_net_),
            .in3(N__24017),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_9_17_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_9_17_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_9_17_6  (
            .in0(N__24010),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14683),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_9_17_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_9_17_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__24007),
            .in2(_gnd_net_),
            .in3(N__15999),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_1_3_LC_9_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_1_3_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_1_3_LC_9_18_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_1_3_LC_9_18_2  (
            .in0(N__15728),
            .in1(N__15671),
            .in2(N__15619),
            .in3(N__15439),
            .lcout(\this_ppu.m35_i_0_a3_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_18_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_18_3 .LUT_INIT=16'b0001110100100101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_18_3  (
            .in0(N__18342),
            .in1(N__18294),
            .in2(N__18394),
            .in3(N__18428),
            .lcout(\this_vga_ramdac.i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_4_LC_9_18_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_4_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_4_LC_9_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_4_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14830),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42062),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNI61SIV_1_LC_9_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNI61SIV_1_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNI61SIV_1_LC_9_19_0 .LUT_INIT=16'b1010000000101000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNI61SIV_1_LC_9_19_0  (
            .in0(N__14894),
            .in1(N__16609),
            .in2(N__15441),
            .in3(N__14857),
            .lcout(\this_ppu.N_985_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNIU85NV_2_LC_9_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNIU85NV_2_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNIU85NV_2_LC_9_19_1 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNIU85NV_2_LC_9_19_1  (
            .in0(N__15571),
            .in1(N__15678),
            .in2(_gnd_net_),
            .in3(N__14895),
            .lcout(\this_ppu.N_671_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIK7UCK_3_LC_9_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIK7UCK_3_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIK7UCK_3_LC_9_19_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_state_q_RNIK7UCK_3_LC_9_19_2  (
            .in0(N__16566),
            .in1(N__22117),
            .in2(N__24164),
            .in3(N__17497),
            .lcout(\this_ppu.N_426_0 ),
            .ltout(\this_ppu.N_426_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNI1KGLK_1_LC_9_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNI1KGLK_1_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNI1KGLK_1_LC_9_19_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNI1KGLK_1_LC_9_19_3  (
            .in0(N__16608),
            .in1(_gnd_net_),
            .in2(N__14794),
            .in3(N__15431),
            .lcout(\this_ppu.un1_M_oam_curr_q_1_c2 ),
            .ltout(\this_ppu.un1_M_oam_curr_q_1_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNINHERV_3_LC_9_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNINHERV_3_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNINHERV_3_LC_9_19_4 .LUT_INIT=16'b0100100010001000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNINHERV_3_LC_9_19_4  (
            .in0(N__15747),
            .in1(N__14896),
            .in2(N__14791),
            .in3(N__15676),
            .lcout(\this_ppu.N_986_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNII43UK_3_LC_9_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNII43UK_3_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNII43UK_3_LC_9_19_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNII43UK_3_LC_9_19_6  (
            .in0(N__15746),
            .in1(N__15675),
            .in2(_gnd_net_),
            .in3(N__15570),
            .lcout(\this_ppu.un1_M_oam_curr_q_1_c4 ),
            .ltout(\this_ppu.un1_M_oam_curr_q_1_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_4_LC_9_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_4_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_4_LC_9_19_7 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \this_ppu.M_oam_curr_q_4_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__15615),
            .in2(N__14773),
            .in3(N__15835),
            .lcout(M_this_ppu_oam_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42073),
            .ce(),
            .sr(N__41651));
    defparam \this_ppu.M_oam_curr_q_0_LC_9_20_0 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_0_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_0_LC_9_20_0 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \this_ppu.M_oam_curr_q_0_LC_9_20_0  (
            .in0(N__14855),
            .in1(N__16624),
            .in2(_gnd_net_),
            .in3(N__15845),
            .lcout(M_this_ppu_oam_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42086),
            .ce(),
            .sr(N__41648));
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_i_a3_LC_9_20_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_i_a3_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_i_a3_LC_9_20_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m13_0_i_a3_LC_9_20_1  (
            .in0(N__23112),
            .in1(N__24318),
            .in2(_gnd_net_),
            .in3(N__25906),
            .lcout(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0 ),
            .ltout(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIVDVLA_4_LC_9_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIVDVLA_4_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIVDVLA_4_LC_9_20_2 .LUT_INIT=16'b0000111100000011;
    LogicCell40 \this_ppu.M_state_q_RNIVDVLA_4_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__22185),
            .in2(N__14899),
            .in3(N__24429),
            .lcout(\this_ppu.M_oam_curr_qc_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI5DBTA_4_LC_9_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI5DBTA_4_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI5DBTA_4_LC_9_20_3 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \this_ppu.M_state_q_RNI5DBTA_4_LC_9_20_3  (
            .in0(N__24428),
            .in1(N__43223),
            .in2(N__22186),
            .in3(N__24569),
            .lcout(\this_ppu.N_841_0 ),
            .ltout(\this_ppu.N_841_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNIFQIEV_0_LC_9_20_4 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNIFQIEV_0_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNIFQIEV_0_LC_9_20_4 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNIFQIEV_0_LC_9_20_4  (
            .in0(N__14854),
            .in1(_gnd_net_),
            .in2(N__14878),
            .in3(N__16623),
            .lcout(\this_ppu.N_669_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_1_LC_9_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_1_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_1_LC_9_20_5 .LUT_INIT=16'b1010101000101010;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_o2_1_LC_9_20_5  (
            .in0(N__29791),
            .in1(N__35014),
            .in2(N__26236),
            .in3(N__30699),
            .lcout(),
            .ltout(\this_ppu.m18_i_o2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_LC_9_20_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_LC_9_20_6 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_o2_LC_9_20_6  (
            .in0(N__30700),
            .in1(N__26200),
            .in2(N__14860),
            .in3(N__34751),
            .lcout(N_792_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_1_LC_9_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_1_LC_9_20_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_1_LC_9_20_7 .LUT_INIT=16'b1000100000101000;
    LogicCell40 \this_ppu.M_oam_curr_q_1_LC_9_20_7  (
            .in0(N__15846),
            .in1(N__15435),
            .in2(N__16632),
            .in3(N__14856),
            .lcout(M_this_ppu_oam_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42086),
            .ce(),
            .sr(N__41648));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIK68L03_9_LC_9_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIK68L03_9_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIK68L03_9_LC_9_21_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIK68L03_9_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__18105),
            .in2(_gnd_net_),
            .in3(N__16090),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_2_LC_9_21_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_2_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_2_LC_9_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_2_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15049),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42098),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_9_21_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_9_21_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_9_21_2  (
            .in0(N__24114),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16408),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_9_21_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_9_21_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_9_21_4  (
            .in0(N__24115),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16135),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_4_LC_9_21_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_4_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_4_LC_9_21_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_4_LC_9_21_6  (
            .in0(N__15021),
            .in1(N__21636),
            .in2(N__15006),
            .in3(N__15324),
            .lcout(\this_ppu.m28_e_i_a3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_9_21_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_9_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__14986),
            .in2(_gnd_net_),
            .in3(N__24113),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_warmup_d_cry_1_c_LC_9_22_0.C_ON=1'b1;
    defparam un1_M_this_warmup_d_cry_1_c_LC_9_22_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_warmup_d_cry_1_c_LC_9_22_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_warmup_d_cry_1_c_LC_9_22_0 (
            .in0(_gnd_net_),
            .in1(N__14962),
            .in2(N__14947),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(un1_M_this_warmup_d_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_warmup_q_2_LC_9_22_1.C_ON=1'b1;
    defparam M_this_warmup_q_2_LC_9_22_1.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_2_LC_9_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_2_LC_9_22_1 (
            .in0(_gnd_net_),
            .in1(N__14926),
            .in2(_gnd_net_),
            .in3(N__14920),
            .lcout(M_this_warmup_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_1),
            .carryout(un1_M_this_warmup_d_cry_2),
            .clk(N__42105),
            .ce(),
            .sr(N__43123));
    defparam M_this_warmup_q_3_LC_9_22_2.C_ON=1'b1;
    defparam M_this_warmup_q_3_LC_9_22_2.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_3_LC_9_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_3_LC_9_22_2 (
            .in0(_gnd_net_),
            .in1(N__14917),
            .in2(_gnd_net_),
            .in3(N__14911),
            .lcout(M_this_warmup_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_2),
            .carryout(un1_M_this_warmup_d_cry_3),
            .clk(N__42105),
            .ce(),
            .sr(N__43123));
    defparam M_this_warmup_q_4_LC_9_22_3.C_ON=1'b1;
    defparam M_this_warmup_q_4_LC_9_22_3.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_4_LC_9_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_4_LC_9_22_3 (
            .in0(_gnd_net_),
            .in1(N__14908),
            .in2(_gnd_net_),
            .in3(N__14902),
            .lcout(M_this_warmup_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_3),
            .carryout(un1_M_this_warmup_d_cry_4),
            .clk(N__42105),
            .ce(),
            .sr(N__43123));
    defparam M_this_warmup_q_5_LC_9_22_4.C_ON=1'b1;
    defparam M_this_warmup_q_5_LC_9_22_4.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_5_LC_9_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_5_LC_9_22_4 (
            .in0(_gnd_net_),
            .in1(N__15121),
            .in2(_gnd_net_),
            .in3(N__15115),
            .lcout(M_this_warmup_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_4),
            .carryout(un1_M_this_warmup_d_cry_5),
            .clk(N__42105),
            .ce(),
            .sr(N__43123));
    defparam M_this_warmup_q_6_LC_9_22_5.C_ON=1'b1;
    defparam M_this_warmup_q_6_LC_9_22_5.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_6_LC_9_22_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_6_LC_9_22_5 (
            .in0(_gnd_net_),
            .in1(N__15112),
            .in2(_gnd_net_),
            .in3(N__15106),
            .lcout(M_this_warmup_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_5),
            .carryout(un1_M_this_warmup_d_cry_6),
            .clk(N__42105),
            .ce(),
            .sr(N__43123));
    defparam M_this_warmup_q_7_LC_9_22_6.C_ON=1'b1;
    defparam M_this_warmup_q_7_LC_9_22_6.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_7_LC_9_22_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_7_LC_9_22_6 (
            .in0(_gnd_net_),
            .in1(N__15103),
            .in2(_gnd_net_),
            .in3(N__15097),
            .lcout(M_this_warmup_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_6),
            .carryout(un1_M_this_warmup_d_cry_7),
            .clk(N__42105),
            .ce(),
            .sr(N__43123));
    defparam M_this_warmup_q_8_LC_9_22_7.C_ON=1'b1;
    defparam M_this_warmup_q_8_LC_9_22_7.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_8_LC_9_22_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_8_LC_9_22_7 (
            .in0(_gnd_net_),
            .in1(N__15094),
            .in2(_gnd_net_),
            .in3(N__15088),
            .lcout(M_this_warmup_qZ0Z_8),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_7),
            .carryout(un1_M_this_warmup_d_cry_8),
            .clk(N__42105),
            .ce(),
            .sr(N__43123));
    defparam M_this_warmup_q_9_LC_9_23_0.C_ON=1'b1;
    defparam M_this_warmup_q_9_LC_9_23_0.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_9_LC_9_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_9_LC_9_23_0 (
            .in0(_gnd_net_),
            .in1(N__15085),
            .in2(_gnd_net_),
            .in3(N__15079),
            .lcout(M_this_warmup_qZ0Z_9),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(un1_M_this_warmup_d_cry_9),
            .clk(N__42112),
            .ce(),
            .sr(N__43126));
    defparam M_this_warmup_q_10_LC_9_23_1.C_ON=1'b1;
    defparam M_this_warmup_q_10_LC_9_23_1.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_10_LC_9_23_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_10_LC_9_23_1 (
            .in0(_gnd_net_),
            .in1(N__15076),
            .in2(_gnd_net_),
            .in3(N__15070),
            .lcout(M_this_warmup_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_9),
            .carryout(un1_M_this_warmup_d_cry_10),
            .clk(N__42112),
            .ce(),
            .sr(N__43126));
    defparam M_this_warmup_q_11_LC_9_23_2.C_ON=1'b1;
    defparam M_this_warmup_q_11_LC_9_23_2.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_11_LC_9_23_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_11_LC_9_23_2 (
            .in0(_gnd_net_),
            .in1(N__15067),
            .in2(_gnd_net_),
            .in3(N__15061),
            .lcout(M_this_warmup_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_10),
            .carryout(un1_M_this_warmup_d_cry_11),
            .clk(N__42112),
            .ce(),
            .sr(N__43126));
    defparam M_this_warmup_q_12_LC_9_23_3.C_ON=1'b1;
    defparam M_this_warmup_q_12_LC_9_23_3.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_12_LC_9_23_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_12_LC_9_23_3 (
            .in0(_gnd_net_),
            .in1(N__15058),
            .in2(_gnd_net_),
            .in3(N__15052),
            .lcout(M_this_warmup_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_11),
            .carryout(un1_M_this_warmup_d_cry_12),
            .clk(N__42112),
            .ce(),
            .sr(N__43126));
    defparam M_this_warmup_q_13_LC_9_23_4.C_ON=1'b1;
    defparam M_this_warmup_q_13_LC_9_23_4.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_13_LC_9_23_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_13_LC_9_23_4 (
            .in0(_gnd_net_),
            .in1(N__15199),
            .in2(_gnd_net_),
            .in3(N__15193),
            .lcout(M_this_warmup_qZ0Z_13),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_12),
            .carryout(un1_M_this_warmup_d_cry_13),
            .clk(N__42112),
            .ce(),
            .sr(N__43126));
    defparam M_this_warmup_q_14_LC_9_23_5.C_ON=1'b1;
    defparam M_this_warmup_q_14_LC_9_23_5.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_14_LC_9_23_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_14_LC_9_23_5 (
            .in0(_gnd_net_),
            .in1(N__15190),
            .in2(_gnd_net_),
            .in3(N__15184),
            .lcout(M_this_warmup_qZ0Z_14),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_13),
            .carryout(un1_M_this_warmup_d_cry_14),
            .clk(N__42112),
            .ce(),
            .sr(N__43126));
    defparam M_this_warmup_q_15_LC_9_23_6.C_ON=1'b1;
    defparam M_this_warmup_q_15_LC_9_23_6.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_15_LC_9_23_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_15_LC_9_23_6 (
            .in0(_gnd_net_),
            .in1(N__15181),
            .in2(_gnd_net_),
            .in3(N__15175),
            .lcout(M_this_warmup_qZ0Z_15),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_14),
            .carryout(un1_M_this_warmup_d_cry_15),
            .clk(N__42112),
            .ce(),
            .sr(N__43126));
    defparam M_this_warmup_q_16_LC_9_23_7.C_ON=1'b1;
    defparam M_this_warmup_q_16_LC_9_23_7.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_16_LC_9_23_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_16_LC_9_23_7 (
            .in0(_gnd_net_),
            .in1(N__15172),
            .in2(_gnd_net_),
            .in3(N__15166),
            .lcout(M_this_warmup_qZ0Z_16),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_15),
            .carryout(un1_M_this_warmup_d_cry_16),
            .clk(N__42112),
            .ce(),
            .sr(N__43126));
    defparam M_this_warmup_q_17_LC_9_24_0.C_ON=1'b1;
    defparam M_this_warmup_q_17_LC_9_24_0.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_17_LC_9_24_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_17_LC_9_24_0 (
            .in0(_gnd_net_),
            .in1(N__15163),
            .in2(_gnd_net_),
            .in3(N__15157),
            .lcout(M_this_warmup_qZ0Z_17),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(un1_M_this_warmup_d_cry_17),
            .clk(N__42119),
            .ce(),
            .sr(N__43130));
    defparam M_this_warmup_q_18_LC_9_24_1.C_ON=1'b1;
    defparam M_this_warmup_q_18_LC_9_24_1.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_18_LC_9_24_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_18_LC_9_24_1 (
            .in0(_gnd_net_),
            .in1(N__15154),
            .in2(_gnd_net_),
            .in3(N__15148),
            .lcout(M_this_warmup_qZ0Z_18),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_17),
            .carryout(un1_M_this_warmup_d_cry_18),
            .clk(N__42119),
            .ce(),
            .sr(N__43130));
    defparam M_this_warmup_q_19_LC_9_24_2.C_ON=1'b1;
    defparam M_this_warmup_q_19_LC_9_24_2.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_19_LC_9_24_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_19_LC_9_24_2 (
            .in0(_gnd_net_),
            .in1(N__15145),
            .in2(_gnd_net_),
            .in3(N__15139),
            .lcout(M_this_warmup_qZ0Z_19),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_18),
            .carryout(un1_M_this_warmup_d_cry_19),
            .clk(N__42119),
            .ce(),
            .sr(N__43130));
    defparam M_this_warmup_q_20_LC_9_24_3.C_ON=1'b1;
    defparam M_this_warmup_q_20_LC_9_24_3.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_20_LC_9_24_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_20_LC_9_24_3 (
            .in0(_gnd_net_),
            .in1(N__15136),
            .in2(_gnd_net_),
            .in3(N__15130),
            .lcout(M_this_warmup_qZ0Z_20),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_19),
            .carryout(un1_M_this_warmup_d_cry_20),
            .clk(N__42119),
            .ce(),
            .sr(N__43130));
    defparam M_this_warmup_q_21_LC_9_24_4.C_ON=1'b1;
    defparam M_this_warmup_q_21_LC_9_24_4.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_21_LC_9_24_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_21_LC_9_24_4 (
            .in0(_gnd_net_),
            .in1(N__15127),
            .in2(_gnd_net_),
            .in3(N__15265),
            .lcout(M_this_warmup_qZ0Z_21),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_20),
            .carryout(un1_M_this_warmup_d_cry_21),
            .clk(N__42119),
            .ce(),
            .sr(N__43130));
    defparam M_this_warmup_q_22_LC_9_24_5.C_ON=1'b1;
    defparam M_this_warmup_q_22_LC_9_24_5.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_22_LC_9_24_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_22_LC_9_24_5 (
            .in0(_gnd_net_),
            .in1(N__15262),
            .in2(_gnd_net_),
            .in3(N__15256),
            .lcout(M_this_warmup_qZ0Z_22),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_21),
            .carryout(un1_M_this_warmup_d_cry_22),
            .clk(N__42119),
            .ce(),
            .sr(N__43130));
    defparam M_this_warmup_q_23_LC_9_24_6.C_ON=1'b1;
    defparam M_this_warmup_q_23_LC_9_24_6.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_23_LC_9_24_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_23_LC_9_24_6 (
            .in0(_gnd_net_),
            .in1(N__15253),
            .in2(_gnd_net_),
            .in3(N__15247),
            .lcout(M_this_warmup_qZ0Z_23),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_22),
            .carryout(un1_M_this_warmup_d_cry_23),
            .clk(N__42119),
            .ce(),
            .sr(N__43130));
    defparam M_this_warmup_q_24_LC_9_24_7.C_ON=1'b1;
    defparam M_this_warmup_q_24_LC_9_24_7.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_24_LC_9_24_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_24_LC_9_24_7 (
            .in0(_gnd_net_),
            .in1(N__15244),
            .in2(_gnd_net_),
            .in3(N__15238),
            .lcout(M_this_warmup_qZ0Z_24),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_23),
            .carryout(un1_M_this_warmup_d_cry_24),
            .clk(N__42119),
            .ce(),
            .sr(N__43130));
    defparam M_this_warmup_q_25_LC_9_25_0.C_ON=1'b1;
    defparam M_this_warmup_q_25_LC_9_25_0.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_25_LC_9_25_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_25_LC_9_25_0 (
            .in0(_gnd_net_),
            .in1(N__15235),
            .in2(_gnd_net_),
            .in3(N__15229),
            .lcout(M_this_warmup_qZ0Z_25),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(un1_M_this_warmup_d_cry_25),
            .clk(N__42123),
            .ce(),
            .sr(N__43131));
    defparam M_this_warmup_q_26_LC_9_25_1.C_ON=1'b1;
    defparam M_this_warmup_q_26_LC_9_25_1.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_26_LC_9_25_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_26_LC_9_25_1 (
            .in0(_gnd_net_),
            .in1(N__15226),
            .in2(_gnd_net_),
            .in3(N__15220),
            .lcout(M_this_warmup_qZ0Z_26),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_25),
            .carryout(un1_M_this_warmup_d_cry_26),
            .clk(N__42123),
            .ce(),
            .sr(N__43131));
    defparam M_this_warmup_q_27_LC_9_25_2.C_ON=1'b0;
    defparam M_this_warmup_q_27_LC_9_25_2.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_27_LC_9_25_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 M_this_warmup_q_27_LC_9_25_2 (
            .in0(_gnd_net_),
            .in1(N__15213),
            .in2(_gnd_net_),
            .in3(N__15217),
            .lcout(M_this_warmup_qZ0Z_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42123),
            .ce(),
            .sr(N__43131));
    defparam M_this_status_flags_q_0_LC_9_25_3.C_ON=1'b0;
    defparam M_this_status_flags_q_0_LC_9_25_3.SEQ_MODE=4'b1000;
    defparam M_this_status_flags_q_0_LC_9_25_3.LUT_INIT=16'b1111111110101010;
    LogicCell40 M_this_status_flags_q_0_LC_9_25_3 (
            .in0(N__15214),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21856),
            .lcout(M_this_status_flags_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42123),
            .ce(),
            .sr(N__43131));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_18_LC_9_26_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_18_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_18_LC_9_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_18_LC_9_26_0  (
            .in0(_gnd_net_),
            .in1(N__26731),
            .in2(_gnd_net_),
            .in3(N__17239),
            .lcout(M_this_oam_ram_write_data_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_23_LC_9_26_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_23_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_23_LC_9_26_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_23_LC_9_26_1  (
            .in0(N__26734),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18163),
            .lcout(M_this_oam_ram_write_data_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_20_LC_9_26_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_20_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_20_LC_9_26_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_20_LC_9_26_3  (
            .in0(N__26733),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17248),
            .lcout(M_this_oam_ram_write_data_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_19_LC_9_26_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_19_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_19_LC_9_26_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_19_LC_9_26_5  (
            .in0(N__26732),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17068),
            .lcout(M_this_oam_ram_write_data_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_17_LC_9_27_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_17_LC_9_27_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_17_LC_9_27_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_17_LC_9_27_6  (
            .in0(_gnd_net_),
            .in1(N__17080),
            .in2(_gnd_net_),
            .in3(N__26643),
            .lcout(M_this_oam_ram_write_data_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_10_16_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_10_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__18253),
            .in2(_gnd_net_),
            .in3(N__17206),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_10_16_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_10_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__24012),
            .in2(_gnd_net_),
            .in3(N__15331),
            .lcout(\this_ppu.oam_cache.N_586_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_10_LC_10_16_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_10_LC_10_16_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_10_LC_10_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_10_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15289),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42024),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o3_LC_10_16_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o3_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o3_LC_10_16_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m28_e_i_o3_LC_10_16_5  (
            .in0(N__16258),
            .in1(N__16240),
            .in2(_gnd_net_),
            .in3(N__16201),
            .lcout(\this_ppu.N_844_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI61M7_10_LC_10_16_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI61M7_10_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI61M7_10_LC_10_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI61M7_10_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15271),
            .lcout(\this_ppu.M_oam_cache_read_data_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_c_LC_10_17_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_c_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_c_LC_10_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_cnt_q_cry_0_c_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__23993),
            .in2(N__16053),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\this_ppu.un1_M_oam_cache_cnt_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_LUT4_0_LC_10_17_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_LUT4_0_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_LUT4_0_LC_10_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_LUT4_0_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__15794),
            .in2(_gnd_net_),
            .in3(N__15490),
            .lcout(\this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_cnt_q_cry_0 ),
            .carryout(\this_ppu.un1_M_oam_cache_cnt_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_LUT4_0_LC_10_17_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_LUT4_0_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_LUT4_0_LC_10_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_LUT4_0_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22643),
            .in3(N__15487),
            .lcout(\this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_cnt_q_cry_1 ),
            .carryout(\this_ppu.un1_M_oam_cache_cnt_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_LUT4_0_LC_10_17_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_LUT4_0_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_LUT4_0_LC_10_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_LUT4_0_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__15523),
            .in2(_gnd_net_),
            .in3(N__15484),
            .lcout(\this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_cnt_q_cry_2 ),
            .carryout(\this_ppu.un1_M_oam_cache_cnt_q_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_cache_cnt_q_4_LC_10_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_oam_cache_cnt_q_4_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_cache_cnt_q_4_LC_10_17_4 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \this_ppu.M_oam_cache_cnt_q_4_LC_10_17_4  (
            .in0(N__15394),
            .in1(N__43237),
            .in2(N__24679),
            .in3(N__15481),
            .lcout(\this_ppu.M_oam_cache_cnt_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42031),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_7_LC_10_17_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_7_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_7_LC_10_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_7_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15478),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42031),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIDR5V3_7_LC_10_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIDR5V3_7_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIDR5V3_7_LC_10_17_7 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIDR5V3_7_LC_10_17_7  (
            .in0(N__39508),
            .in1(N__17929),
            .in2(N__17716),
            .in3(N__16705),
            .lcout(N_41_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_0_LC_10_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_0_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_0_LC_10_18_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_0_LC_10_18_1  (
            .in0(N__15795),
            .in1(N__15672),
            .in2(N__22653),
            .in3(N__15440),
            .lcout(),
            .ltout(\this_ppu.m62_0_a2_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_LC_10_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_LC_10_18_2 .LUT_INIT=16'b1001000000000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_LC_10_18_2  (
            .in0(N__15393),
            .in1(N__15608),
            .in2(N__15376),
            .in3(N__15763),
            .lcout(\this_ppu.N_762_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_3_LC_10_18_3 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_3_LC_10_18_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_3_LC_10_18_3 .LUT_INIT=16'b0110000011000000;
    LogicCell40 \this_ppu.M_oam_curr_q_3_LC_10_18_3  (
            .in0(N__15574),
            .in1(N__15733),
            .in2(N__15853),
            .in3(N__15674),
            .lcout(M_this_ppu_oam_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42040),
            .ce(),
            .sr(N__41649));
    defparam \this_ppu.M_oam_curr_q_2_LC_10_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_2_LC_10_18_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_2_LC_10_18_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_oam_curr_q_2_LC_10_18_4  (
            .in0(N__15673),
            .in1(N__15847),
            .in2(_gnd_net_),
            .in3(N__15573),
            .lcout(M_this_ppu_oam_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42040),
            .ce(),
            .sr(N__41649));
    defparam \this_ppu.M_oam_curr_q_5_LC_10_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_5_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_5_LC_10_18_5 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \this_ppu.M_oam_curr_q_5_LC_10_18_5  (
            .in0(N__15851),
            .in1(N__16662),
            .in2(N__15620),
            .in3(N__15859),
            .lcout(M_this_ppu_oam_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42040),
            .ce(),
            .sr(N__41649));
    defparam \this_ppu.M_oam_curr_q_6_LC_10_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_6_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_6_LC_10_18_6 .LUT_INIT=16'b0100100011000000;
    LogicCell40 \this_ppu.M_oam_curr_q_6_LC_10_18_6  (
            .in0(N__16661),
            .in1(N__15852),
            .in2(N__18713),
            .in3(N__15550),
            .lcout(\this_ppu.M_oam_curr_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42040),
            .ce(),
            .sr(N__41649));
    defparam \this_ppu.M_surface_x_q_RNO_0_7_LC_10_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNO_0_7_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNO_0_7_LC_10_18_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNO_0_7_LC_10_18_7  (
            .in0(N__22904),
            .in1(N__21243),
            .in2(N__23004),
            .in3(N__23271),
            .lcout(\this_ppu.un1_M_surface_x_q_ac0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_cache_cnt_q_1_LC_10_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_oam_cache_cnt_q_1_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_cache_cnt_q_1_LC_10_19_0 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \this_ppu.M_oam_cache_cnt_q_1_LC_10_19_0  (
            .in0(N__15790),
            .in1(N__43238),
            .in2(N__15817),
            .in3(N__24581),
            .lcout(\this_ppu.M_oam_cache_cnt_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42051),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_1_LC_10_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_1_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_1_LC_10_19_2 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_1_LC_10_19_2  (
            .in0(N__15737),
            .in1(N__16607),
            .in2(N__15527),
            .in3(N__16048),
            .lcout(\this_ppu.m62_0_a2_0_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNO_0_6_LC_10_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNO_0_6_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNO_0_6_LC_10_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNO_0_6_LC_10_19_3  (
            .in0(N__15732),
            .in1(N__15677),
            .in2(N__15621),
            .in3(N__15572),
            .lcout(\this_ppu.un1_M_oam_curr_q_1_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_cache_cnt_q_3_LC_10_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_oam_cache_cnt_q_3_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_cache_cnt_q_3_LC_10_19_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \this_ppu.M_oam_cache_cnt_q_3_LC_10_19_4  (
            .in0(N__15544),
            .in1(N__43239),
            .in2(N__15528),
            .in3(N__24582),
            .lcout(\this_ppu.M_oam_cache_cnt_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42051),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_10_19_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_10_19_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_10_19_5  (
            .in0(N__24134),
            .in1(N__15961),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_10_19_6 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_10_19_6 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_10_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15937),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42051),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_3_LC_10_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_3_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_3_LC_10_19_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_3_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__15925),
            .in2(_gnd_net_),
            .in3(N__16752),
            .lcout(\this_ppu.m28_e_i_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_10_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_10_20_0 .LUT_INIT=16'b0111010010001011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_10_20_0  (
            .in0(N__17317),
            .in1(N__16098),
            .in2(N__18996),
            .in3(N__15867),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI8I4KS3_1_LC_10_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI8I4KS3_1_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI8I4KS3_1_LC_10_20_1 .LUT_INIT=16'b0111111010000001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI8I4KS3_1_LC_10_20_1  (
            .in0(N__17379),
            .in1(N__17319),
            .in2(N__15898),
            .in3(N__16066),
            .lcout(\this_vga_signals.haddress_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m1_LC_10_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m1_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m1_LC_10_20_2 .LUT_INIT=16'b0010000111011110;
    LogicCell40 \this_vga_signals.un4_haddress_if_m1_LC_10_20_2  (
            .in0(N__17318),
            .in1(N__16099),
            .in2(N__18997),
            .in3(N__15868),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_10_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_10_20_3 .LUT_INIT=16'b0011110100110100;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_m2_LC_10_20_3  (
            .in0(N__16921),
            .in1(N__17383),
            .in2(N__15895),
            .in3(N__17425),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un89_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI4NUA8C_1_LC_10_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI4NUA8C_1_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI4NUA8C_1_LC_10_20_4 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI4NUA8C_1_LC_10_20_4  (
            .in0(N__18091),
            .in1(N__16809),
            .in2(N__15892),
            .in3(N__15889),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0_LC_10_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0_LC_10_20_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__17605),
            .in2(_gnd_net_),
            .in3(N__16955),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_20_6 .LUT_INIT=16'b1101111000000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_20_6  (
            .in0(N__18553),
            .in1(N__19042),
            .in2(N__18061),
            .in3(N__16966),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m2_LC_10_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m2_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m2_LC_10_20_7 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \this_vga_signals.un4_haddress_if_m2_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16102),
            .in3(N__19120),
            .lcout(\this_vga_signals.if_m2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_a2_LC_10_21_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_a2_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_a2_LC_10_21_0 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_a2_LC_10_21_0  (
            .in0(N__16233),
            .in1(N__16254),
            .in2(N__23249),
            .in3(N__16194),
            .lcout(\this_ppu.N_1394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIDPGC47_9_LC_10_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIDPGC47_9_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIDPGC47_9_LC_10_21_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIDPGC47_9_LC_10_21_1  (
            .in0(N__18096),
            .in1(N__16089),
            .in2(_gnd_net_),
            .in3(N__16813),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_10_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_10_21_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__19126),
            .in2(_gnd_net_),
            .in3(N__16958),
            .lcout(\this_vga_signals.mult1_un75_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_cache_cnt_q_0_LC_10_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_oam_cache_cnt_q_0_LC_10_21_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_cache_cnt_q_0_LC_10_21_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \this_ppu.M_oam_cache_cnt_q_0_LC_10_21_5  (
            .in0(N__24135),
            .in1(N__43240),
            .in2(N__16049),
            .in3(N__24580),
            .lcout(\this_ppu.M_oam_cache_cnt_qZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42074),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1INF21_9_LC_10_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1INF21_9_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1INF21_9_LC_10_21_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI1INF21_9_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__18097),
            .in2(_gnd_net_),
            .in3(N__16959),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_0_c_inv_LC_10_22_0 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_0_c_inv_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_0_c_inv_LC_10_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_0_c_inv_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__15973),
            .in2(N__21585),
            .in3(N__16000),
            .lcout(\this_ppu.M_this_oam_ram_read_data_i_16 ),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\this_ppu.un1_oam_data_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_1_c_inv_LC_10_22_1 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_1_c_inv_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_1_c_inv_LC_10_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_1_c_inv_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__15967),
            .in2(N__21540),
            .in3(N__17010),
            .lcout(\this_ppu.M_this_oam_ram_read_data_i_17 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_0 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_2_c_inv_LC_10_22_2 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_2_c_inv_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_2_c_inv_LC_10_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_2_c_inv_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__16270),
            .in2(N__21504),
            .in3(N__16182),
            .lcout(\this_ppu.M_this_oam_ram_read_data_i_18 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_1 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_2_c_RNIR4HD_LC_10_22_3 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_2_c_RNIR4HD_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_2_c_RNIR4HD_LC_10_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_2_c_RNIR4HD_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__16324),
            .in2(N__21468),
            .in3(N__16264),
            .lcout(\this_ppu.un1_oam_data_1_cry_2_c_RNIR4HDZ0 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_2 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_3_c_RNIT7ID_LC_10_22_4 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_3_c_RNIT7ID_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_3_c_RNIT7ID_LC_10_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_3_c_RNIT7ID_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__16537),
            .in2(N__21423),
            .in3(N__16261),
            .lcout(\this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_3 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJD_LC_10_22_5 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJD_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJD_LC_10_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJD_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(N__21378),
            .in2(N__16384),
            .in3(N__16243),
            .lcout(\this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_4 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKD_LC_10_22_6 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKD_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKD_LC_10_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKD_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(N__21330),
            .in2(N__16111),
            .in3(N__16222),
            .lcout(\this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_5 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o3_2_LC_10_22_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o3_2_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o3_2_LC_10_22_7 .LUT_INIT=16'b0000001000000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m28_e_i_o3_2_LC_10_22_7  (
            .in0(N__17059),
            .in1(N__16219),
            .in2(N__16213),
            .in3(N__16204),
            .lcout(\this_ppu.m28_e_i_o3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_10_23_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_10_23_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__24172),
            .in2(_gnd_net_),
            .in3(N__16183),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_5_LC_10_23_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_5_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_5_LC_10_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_5_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(N__26761),
            .in2(_gnd_net_),
            .in3(N__17992),
            .lcout(M_this_oam_ram_write_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_10_23_2 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_10_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16134),
            .lcout(M_this_oam_ram_read_data_i_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_10_23_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_10_23_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_10_23_3  (
            .in0(N__24173),
            .in1(N__16432),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_10_23_4 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_10_23_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16407),
            .lcout(M_this_oam_ram_read_data_i_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_10_23_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_10_23_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_10_23_5  (
            .in0(N__24174),
            .in1(N__16375),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_10_23_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_10_23_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_10_23_6  (
            .in0(N__16339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24175),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_10_23_7 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_10_23_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16338),
            .lcout(M_this_oam_ram_read_data_i_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_10_LC_10_24_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_10_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_10_LC_10_24_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_10_LC_10_24_3  (
            .in0(_gnd_net_),
            .in1(N__16975),
            .in2(_gnd_net_),
            .in3(N__26747),
            .lcout(M_this_oam_ram_write_data_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIML464_9_LC_10_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIML464_9_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIML464_9_LC_10_24_4 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIML464_9_LC_10_24_4  (
            .in0(N__17875),
            .in1(N__16477),
            .in2(N__17805),
            .in3(N__17937),
            .lcout(N_260),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_10_24_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_10_24_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_10_24_6  (
            .in0(_gnd_net_),
            .in1(N__16294),
            .in2(_gnd_net_),
            .in3(N__24171),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_9_LC_10_24_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_9_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_9_LC_10_24_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_9_LC_10_24_7  (
            .in0(N__17137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26748),
            .lcout(M_this_oam_ram_write_data_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_10_25_0 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_10_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17583),
            .lcout(M_this_oam_ram_read_data_i_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_28_LC_10_25_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_28_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_28_LC_10_25_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_28_LC_10_25_1  (
            .in0(_gnd_net_),
            .in1(N__40783),
            .in2(_gnd_net_),
            .in3(N__26726),
            .lcout(M_this_oam_ram_write_data_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_8_LC_10_25_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_8_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_8_LC_10_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_8_LC_10_25_5  (
            .in0(_gnd_net_),
            .in1(N__17143),
            .in2(_gnd_net_),
            .in3(N__26728),
            .lcout(M_this_oam_ram_write_data_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_31_LC_10_25_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_31_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_31_LC_10_25_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_31_LC_10_25_6  (
            .in0(N__26727),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39870),
            .lcout(M_this_oam_ram_write_data_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_16_LC_10_26_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_16_LC_10_26_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_16_LC_10_26_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_16_LC_10_26_4  (
            .in0(N__26730),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17086),
            .lcout(M_this_oam_ram_write_data_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_24_LC_10_26_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_24_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_24_LC_10_26_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_24_LC_10_26_5  (
            .in0(_gnd_net_),
            .in1(N__42416),
            .in2(_gnd_net_),
            .in3(N__26729),
            .lcout(M_this_oam_ram_write_data_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIOC7D3_6_LC_11_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIOC7D3_6_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIOC7D3_6_LC_11_16_0 .LUT_INIT=16'b0101010111110011;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIOC7D3_6_LC_11_16_0  (
            .in0(N__17431),
            .in1(N__16438),
            .in2(N__19224),
            .in3(N__17707),
            .lcout(\this_vga_signals.hsync_1_i_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_11_16_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_11_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__16465),
            .in2(_gnd_net_),
            .in3(N__24140),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI69GD1_0_LC_11_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI69GD1_0_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI69GD1_0_LC_11_16_7 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI69GD1_0_LC_11_16_7  (
            .in0(N__17443),
            .in1(N__17358),
            .in2(N__18620),
            .in3(N__17417),
            .lcout(\this_vga_signals.hsync_1_i_0_0_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_11_17_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_11_17_2 .LUT_INIT=16'b0011000110010111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_11_17_2  (
            .in0(N__18353),
            .in1(N__18303),
            .in2(N__18404),
            .in3(N__18437),
            .lcout(\this_vga_ramdac.m16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_11_17_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_11_17_3 .LUT_INIT=16'b0001110110100011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_11_17_3  (
            .in0(N__18438),
            .in1(N__18354),
            .in2(N__18307),
            .in3(N__18398),
            .lcout(\this_vga_ramdac.m19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_11_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_11_17_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__17773),
            .in2(_gnd_net_),
            .in3(N__17855),
            .lcout(\this_vga_signals.N_811_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_11_17_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_11_17_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_11_17_7  (
            .in0(N__18211),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17207),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_1_LC_11_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_1_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_1_LC_11_18_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_1_LC_11_18_1  (
            .in0(N__16660),
            .in1(N__16631),
            .in2(_gnd_net_),
            .in3(N__16576),
            .lcout(\this_ppu.N_1196_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNITMA41_9_LC_11_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNITMA41_9_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNITMA41_9_LC_11_18_2 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNITMA41_9_LC_11_18_2  (
            .in0(N__17854),
            .in1(N__17915),
            .in2(N__30472),
            .in3(N__17769),
            .lcout(\this_vga_signals.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_1_LC_11_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_1_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_1_LC_11_18_4 .LUT_INIT=16'b0101010101010001;
    LogicCell40 \this_ppu.M_state_q_1_LC_11_18_4  (
            .in0(N__26135),
            .in1(N__16819),
            .in2(N__24183),
            .in3(N__16567),
            .lcout(\this_ppu.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42032),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_5_LC_11_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_5_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_5_LC_11_18_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIF4AR_5_LC_11_18_6  (
            .in0(N__17702),
            .in1(N__18594),
            .in2(_gnd_net_),
            .in3(N__17914),
            .lcout(\this_vga_signals.M_hcounter_d7_0_i_0_o3_0_o3_4_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_11_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_11_18_7 .LUT_INIT=16'b0110101000101000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_11_18_7  (
            .in0(N__17844),
            .in1(N__17905),
            .in2(N__17784),
            .in3(N__17701),
            .lcout(\this_vga_signals.N_291_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_LC_11_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_LC_11_19_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_LC_11_19_0  (
            .in0(N__16864),
            .in1(N__16840),
            .in2(N__16786),
            .in3(N__16828),
            .lcout(\this_ppu.N_1184_7 ),
            .ltout(\this_ppu.N_1184_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_1_LC_11_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_1_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_1_LC_11_19_1 .LUT_INIT=16'b0000000100110011;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_1_LC_11_19_1  (
            .in0(N__24270),
            .in1(N__16720),
            .in2(N__16822),
            .in3(N__23250),
            .lcout(\this_ppu.m18_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_2_LC_11_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_2_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_2_LC_11_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_2_LC_11_19_2  (
            .in0(N__16711),
            .in1(N__16930),
            .in2(N__17956),
            .in3(N__16960),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_12_LC_11_19_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_12_LC_11_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_12_LC_11_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_12_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16798),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42041),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_11_19_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_11_19_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_11_19_4  (
            .in0(N__16785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24095),
            .lcout(\this_ppu.oam_cache.N_569_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_11_19_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_11_19_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_11_19_5  (
            .in0(N__24094),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16753),
            .lcout(\this_ppu.oam_cache.N_575_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_a3_LC_11_20_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_a3_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_a3_LC_11_20_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_a3_LC_11_20_0  (
            .in0(N__23113),
            .in1(N__24319),
            .in2(N__21885),
            .in3(N__25916),
            .lcout(\this_ppu.N_1182 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_11_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_11_20_1 .LUT_INIT=16'b0001011100101011;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_11_20_1  (
            .in0(N__17635),
            .in1(N__17305),
            .in2(N__17378),
            .in3(N__17604),
            .lcout(),
            .ltout(\this_vga_signals.if_N_9_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_11_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_11_20_2 .LUT_INIT=16'b0000011010011111;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_11_20_2  (
            .in0(N__16957),
            .in1(N__19122),
            .in2(N__16714),
            .in3(N__17320),
            .lcout(\this_vga_signals.mult1_un82_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_11_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_11_20_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_11_20_3  (
            .in0(N__19225),
            .in1(N__19149),
            .in2(_gnd_net_),
            .in3(N__19030),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_2 ),
            .ltout(\this_vga_signals.mult1_un68_sum_ac0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_1_LC_11_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_1_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_1_LC_11_20_4 .LUT_INIT=16'b0011011100111111;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_1_LC_11_20_4  (
            .in0(N__19119),
            .in1(N__17616),
            .in2(N__16969),
            .in3(N__17634),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_11_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_11_20_5 .LUT_INIT=16'b0010001010111011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_11_20_5  (
            .in0(N__19121),
            .in1(N__17306),
            .in2(_gnd_net_),
            .in3(N__16956),
            .lcout(\this_vga_signals.mult1_un75_sum_c2_0 ),
            .ltout(\this_vga_signals.mult1_un75_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_LC_11_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_LC_11_20_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_x4_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__17952),
            .in2(N__16924),
            .in3(N__19123),
            .lcout(\this_vga_signals.if_N_8_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_11_21_0 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_11_21_0 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_11_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16915),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42063),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI8F2M3_9_LC_11_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI8F2M3_9_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI8F2M3_9_LC_11_21_2 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI8F2M3_9_LC_11_21_2  (
            .in0(N__17787),
            .in1(N__17870),
            .in2(N__39507),
            .in3(N__17930),
            .lcout(N_852_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_11_22_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_11_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__16903),
            .in2(_gnd_net_),
            .in3(N__24163),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_0_LC_11_22_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_0_LC_11_22_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_0_LC_11_22_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_ppu.oam_cache.read_data_0_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__16876),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42075),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_o2_1_LC_11_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_o2_1_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_o2_1_LC_11_22_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.IO_port_data_write_0_a2_i_o2_1_LC_11_22_3  (
            .in0(N__29248),
            .in1(N__27172),
            .in2(N__36358),
            .in3(N__29290),
            .lcout(\this_vga_signals.N_834_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_y_q_esr_RNICCL8_7_LC_11_22_5 .C_ON=1'b0;
    defparam \this_ppu.M_surface_y_q_esr_RNICCL8_7_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_y_q_esr_RNICCL8_7_LC_11_22_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_ppu.M_surface_y_q_esr_RNICCL8_7_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__21705),
            .in2(_gnd_net_),
            .in3(N__21672),
            .lcout(\this_ppu.un1_oam_data_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_6_LC_11_23_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_6_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_6_LC_11_23_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_6_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__17035),
            .in2(_gnd_net_),
            .in3(N__26759),
            .lcout(M_this_oam_ram_write_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_6_LC_11_23_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_6_LC_11_23_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_6_LC_11_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_6_LC_11_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40415),
            .lcout(M_this_data_tmp_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42087),
            .ce(N__25686),
            .sr(N__43119));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_7_LC_11_23_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_7_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_7_LC_11_23_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_7_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(N__17017),
            .in2(_gnd_net_),
            .in3(N__26760),
            .lcout(M_this_oam_ram_write_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_7_LC_11_23_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_7_LC_11_23_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_7_LC_11_23_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_7_LC_11_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39926),
            .lcout(M_this_data_tmp_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42087),
            .ce(N__25686),
            .sr(N__43119));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_11_23_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_11_23_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_11_23_7  (
            .in0(N__24177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17011),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_11_LC_11_24_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_11_LC_11_24_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_11_LC_11_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_11_LC_11_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41513),
            .lcout(M_this_data_tmp_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42099),
            .ce(N__26563),
            .sr(N__43122));
    defparam M_this_data_tmp_q_esr_10_LC_11_24_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_10_LC_11_24_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_10_LC_11_24_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_10_LC_11_24_4 (
            .in0(N__42796),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42099),
            .ce(N__26563),
            .sr(N__43122));
    defparam M_this_data_tmp_q_esr_15_LC_11_24_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_15_LC_11_24_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_15_LC_11_24_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_15_LC_11_24_5 (
            .in0(N__39927),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42099),
            .ce(N__26563),
            .sr(N__43122));
    defparam M_this_data_tmp_q_esr_8_LC_11_24_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_8_LC_11_24_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_8_LC_11_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_8_LC_11_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42429),
            .lcout(M_this_data_tmp_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42099),
            .ce(N__26563),
            .sr(N__43122));
    defparam M_this_data_tmp_q_esr_9_LC_11_24_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_9_LC_11_24_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_9_LC_11_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_9_LC_11_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39760),
            .lcout(M_this_data_tmp_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42099),
            .ce(N__26563),
            .sr(N__43122));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_26_LC_11_25_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_26_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_26_LC_11_25_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_26_LC_11_25_0  (
            .in0(N__42792),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26722),
            .lcout(M_this_oam_ram_write_data_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_27_LC_11_25_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_27_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_27_LC_11_25_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_27_LC_11_25_2  (
            .in0(N__41512),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26723),
            .lcout(M_this_oam_ram_write_data_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_30_LC_11_25_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_30_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_30_LC_11_25_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_30_LC_11_25_6  (
            .in0(_gnd_net_),
            .in1(N__40435),
            .in2(_gnd_net_),
            .in3(N__26724),
            .lcout(M_this_oam_ram_write_data_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_15_LC_11_25_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_15_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_15_LC_11_25_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_15_LC_11_25_7  (
            .in0(N__26725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17104),
            .lcout(M_this_oam_ram_write_data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_16_LC_11_26_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_16_LC_11_26_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_16_LC_11_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_16_LC_11_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42415),
            .lcout(M_this_data_tmp_qZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42113),
            .ce(N__25632),
            .sr(N__43127));
    defparam M_this_data_tmp_q_esr_17_LC_11_26_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_17_LC_11_26_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_17_LC_11_26_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_17_LC_11_26_1 (
            .in0(N__39728),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42113),
            .ce(N__25632),
            .sr(N__43127));
    defparam M_this_data_tmp_q_esr_19_LC_11_26_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_19_LC_11_26_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_19_LC_11_26_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_19_LC_11_26_2 (
            .in0(N__41511),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42113),
            .ce(N__25632),
            .sr(N__43127));
    defparam M_this_data_tmp_q_esr_20_LC_11_26_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_20_LC_11_26_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_20_LC_11_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_20_LC_11_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40782),
            .lcout(M_this_data_tmp_qZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42113),
            .ce(N__25632),
            .sr(N__43127));
    defparam M_this_data_tmp_q_esr_18_LC_11_26_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_18_LC_11_26_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_18_LC_11_26_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_18_LC_11_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42791),
            .lcout(M_this_data_tmp_qZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42113),
            .ce(N__25632),
            .sr(N__43127));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_0_LC_11_27_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_0_LC_11_27_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_0_LC_11_27_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_0_LC_11_27_3  (
            .in0(_gnd_net_),
            .in1(N__18154),
            .in2(_gnd_net_),
            .in3(N__26642),
            .lcout(M_this_oam_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_12_15_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_12_15_3 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_q_ret_LC_12_15_3  (
            .in0(N__20307),
            .in1(N__18109),
            .in2(N__17193),
            .in3(N__26136),
            .lcout(\this_vga_ramdac.N_852_i_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41998),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_12_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_12_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__17284),
            .in2(_gnd_net_),
            .in3(N__19072),
            .lcout(\this_vga_signals.N_298_0 ),
            .ltout(\this_vga_signals.N_298_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_12_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_12_16_1 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_12_16_1  (
            .in0(N__17345),
            .in1(N__17408),
            .in2(N__17158),
            .in3(N__19209),
            .lcout(),
            .ltout(\this_vga_signals.N_1044_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_12_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_12_16_2 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_12_16_2  (
            .in0(N__17155),
            .in1(N__17785),
            .in2(N__17146),
            .in3(N__17853),
            .lcout(\this_vga_signals.M_hcounter_d7_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_12_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_12_16_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_12_16_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_12_16_4  (
            .in0(N__27296),
            .in1(_gnd_net_),
            .in2(N__17418),
            .in3(N__17346),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42005),
            .ce(),
            .sr(N__18682));
    defparam \this_vga_signals.M_hcounter_q_0_LC_12_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_12_16_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__17409),
            .in2(_gnd_net_),
            .in3(N__27295),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42005),
            .ce(),
            .sr(N__18682));
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_1_LC_12_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_1_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_1_LC_12_16_7 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIADGD1_1_LC_12_16_7  (
            .in0(N__17347),
            .in1(N__17442),
            .in2(N__18619),
            .in3(N__19210),
            .lcout(\this_vga_signals.hsync_1_i_0_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_17_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__17416),
            .in2(N__17368),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_17_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_17_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_12_17_1  (
            .in0(N__27291),
            .in1(N__17304),
            .in2(_gnd_net_),
            .in3(N__17269),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__42016),
            .ce(),
            .sr(N__18681));
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_17_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_17_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_17_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_12_17_2  (
            .in0(N__27344),
            .in1(N__19118),
            .in2(_gnd_net_),
            .in3(N__17266),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__42016),
            .ce(),
            .sr(N__18681));
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_17_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_17_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_12_17_3  (
            .in0(N__27292),
            .in1(N__19211),
            .in2(_gnd_net_),
            .in3(N__17263),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__42016),
            .ce(),
            .sr(N__18681));
    defparam \this_vga_signals.M_hcounter_q_5_LC_12_17_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_12_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_12_17_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_12_17_4  (
            .in0(N__27345),
            .in1(N__18603),
            .in2(_gnd_net_),
            .in3(N__17260),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__42016),
            .ce(),
            .sr(N__18681));
    defparam \this_vga_signals.M_hcounter_q_6_LC_12_17_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_12_17_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_12_17_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_12_17_5  (
            .in0(N__27293),
            .in1(N__17706),
            .in2(_gnd_net_),
            .in3(N__17257),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__42016),
            .ce(),
            .sr(N__18681));
    defparam \this_vga_signals.M_hcounter_q_7_LC_12_17_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_12_17_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_12_17_6  (
            .in0(N__27346),
            .in1(N__17916),
            .in2(_gnd_net_),
            .in3(N__17254),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__42016),
            .ce(),
            .sr(N__18681));
    defparam \this_vga_signals.M_hcounter_q_8_LC_12_17_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_12_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_12_17_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_12_17_7  (
            .in0(N__27294),
            .in1(N__17856),
            .in2(_gnd_net_),
            .in3(N__17251),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__42016),
            .ce(),
            .sr(N__18681));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_12_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_12_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_12_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__17774),
            .in2(_gnd_net_),
            .in3(N__17527),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42025),
            .ce(N__18649),
            .sr(N__18674));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_1_0_LC_12_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_1_0_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_1_0_LC_12_19_0 .LUT_INIT=16'b0111111111010011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_1_0_LC_12_19_0  (
            .in0(N__19216),
            .in1(N__17649),
            .in2(N__18621),
            .in3(N__17709),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_LC_12_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_LC_12_19_1 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__17521),
            .in2(N__17524),
            .in3(N__17727),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_tz_LC_12_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_tz_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_tz_LC_12_19_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_tz_LC_12_19_2  (
            .in0(N__18610),
            .in1(N__19215),
            .in2(_gnd_net_),
            .in3(N__17708),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI42MR5_6_LC_12_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI42MR5_6_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI42MR5_6_LC_12_19_3 .LUT_INIT=16'b0111011100000111;
    LogicCell40 \this_ppu.M_state_q_RNI42MR5_6_LC_12_19_3  (
            .in0(N__17508),
            .in1(N__23222),
            .in2(N__23836),
            .in3(N__23786),
            .lcout(\this_ppu.un1_M_state_q_7_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_12_19_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_12_19_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_12_19_4  (
            .in0(N__24096),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17488),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI83M7_12_LC_12_19_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI83M7_12_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI83M7_12_LC_12_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI83M7_12_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17464),
            .lcout(\this_ppu.M_oam_cache_read_data_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_15_LC_12_19_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_15_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_15_LC_12_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_15_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17458),
            .lcout(\this_ppu.M_oam_cache_read_data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42033),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_0_LC_12_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_0_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_0_LC_12_20_0 .LUT_INIT=16'b1100100011101100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_0_LC_12_20_0  (
            .in0(N__17656),
            .in1(N__17728),
            .in2(N__18622),
            .in3(N__17712),
            .lcout(\this_vga_signals.mult1_un54_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb2_LC_12_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb2_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb2_LC_12_20_1 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb2_LC_12_20_1  (
            .in0(N__19028),
            .in1(N__18549),
            .in2(N__17959),
            .in3(N__19150),
            .lcout(\this_vga_signals.mult1_un68_sum_axb2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_12_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_12_20_2 .LUT_INIT=16'b0111100010000111;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_12_20_2  (
            .in0(N__19151),
            .in1(N__19029),
            .in2(N__19125),
            .in3(N__19222),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_12_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_12_20_4 .LUT_INIT=16'b1101101100100100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_12_20_4  (
            .in0(N__17920),
            .in1(N__17860),
            .in2(N__17786),
            .in3(N__17710),
            .lcout(\this_vga_signals.N_968 ),
            .ltout(\this_vga_signals.N_968_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_12_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_12_20_5 .LUT_INIT=16'b0011111111011111;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_12_20_5  (
            .in0(N__17711),
            .in1(N__18614),
            .in2(N__17659),
            .in3(N__17655),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_12_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_12_20_6 .LUT_INIT=16'b1100000000111111;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__19027),
            .in2(N__17638),
            .in3(N__19221),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_12_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_12_20_7 .LUT_INIT=16'b0001001111101100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_12_20_7  (
            .in0(N__19108),
            .in1(N__17626),
            .in2(N__17620),
            .in3(N__17617),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_12_21_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_12_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(N__24181),
            .in2(_gnd_net_),
            .in3(N__17590),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_13_LC_12_21_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_13_LC_12_21_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_13_LC_12_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_13_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17551),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42052),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNILTV6A_9_LC_12_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNILTV6A_9_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNILTV6A_9_LC_12_21_5 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNILTV6A_9_LC_12_21_5  (
            .in0(N__19041),
            .in1(_gnd_net_),
            .in2(N__18104),
            .in3(N__19153),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNINGAC6_9_LC_12_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNINGAC6_9_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNINGAC6_9_LC_12_21_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNINGAC6_9_LC_12_21_7  (
            .in0(N__18092),
            .in1(N__18057),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_0_LC_12_22_0 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_0_LC_12_22_0 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_0_LC_12_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clk.M_counter_q_0_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19256),
            .lcout(this_pixel_clk_M_counter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42064),
            .ce(),
            .sr(N__43116));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_3_LC_12_23_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_3_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_3_LC_12_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_3_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(N__18016),
            .in2(_gnd_net_),
            .in3(N__26739),
            .lcout(M_this_oam_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_3_LC_12_23_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_3_LC_12_23_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_3_LC_12_23_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_3_LC_12_23_4 (
            .in0(N__41515),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42076),
            .ce(N__25685),
            .sr(N__43117));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_4_LC_12_23_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_4_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_4_LC_12_23_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_4_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(N__17998),
            .in2(_gnd_net_),
            .in3(N__26740),
            .lcout(M_this_oam_ram_write_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_4_LC_12_23_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_4_LC_12_23_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_4_LC_12_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_4_LC_12_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40785),
            .lcout(M_this_data_tmp_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42076),
            .ce(N__25685),
            .sr(N__43117));
    defparam M_this_data_tmp_q_esr_5_LC_12_24_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_5_LC_12_24_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_5_LC_12_24_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_5_LC_12_24_3 (
            .in0(N__40058),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42088),
            .ce(N__25687),
            .sr(N__43120));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_29_LC_12_25_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_29_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_29_LC_12_25_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_29_LC_12_25_1  (
            .in0(N__40059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26719),
            .lcout(M_this_oam_ram_write_data_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_21_LC_12_25_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_21_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_21_LC_12_25_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_21_LC_12_25_3  (
            .in0(_gnd_net_),
            .in1(N__18169),
            .in2(_gnd_net_),
            .in3(N__26721),
            .lcout(M_this_oam_ram_write_data_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_1_LC_12_25_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_1_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_1_LC_12_25_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_1_LC_12_25_6  (
            .in0(N__26720),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20227),
            .lcout(M_this_oam_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_25_LC_12_25_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_25_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_25_LC_12_25_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_25_LC_12_25_7  (
            .in0(N__39729),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26718),
            .lcout(M_this_oam_ram_write_data_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_21_LC_12_26_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_21_LC_12_26_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_21_LC_12_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_21_LC_12_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40060),
            .lcout(M_this_data_tmp_qZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42106),
            .ce(N__25631),
            .sr(N__43124));
    defparam M_this_data_tmp_q_esr_23_LC_12_26_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_23_LC_12_26_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_23_LC_12_26_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_23_LC_12_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39931),
            .lcout(M_this_data_tmp_qZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42106),
            .ce(N__25631),
            .sr(N__43124));
    defparam M_this_data_tmp_q_esr_0_LC_12_27_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_0_LC_12_27_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_0_LC_12_27_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_0_LC_12_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42377),
            .lcout(M_this_data_tmp_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42114),
            .ce(N__25681),
            .sr(N__43128));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_13_15_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_13_15_5 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_13_15_5  (
            .in0(N__18454),
            .in1(N__20308),
            .in2(N__18147),
            .in3(N__26115),
            .lcout(\this_vga_ramdac.N_3856_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41992),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_13_16_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_13_16_0 .LUT_INIT=16'b0000011101100111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_13_16_0  (
            .in0(N__18301),
            .in1(N__18349),
            .in2(N__18409),
            .in3(N__18447),
            .lcout(),
            .ltout(\this_vga_ramdac.i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_13_16_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_13_16_1 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_13_16_1  (
            .in0(N__20304),
            .in1(N__26075),
            .in2(N__18130),
            .in3(N__18120),
            .lcout(\this_vga_ramdac.N_3858_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41999),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.G_535_LC_13_16_3 .C_ON=1'b0;
    defparam \this_ppu.G_535_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.G_535_LC_13_16_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_ppu.G_535_LC_13_16_3  (
            .in0(N__19240),
            .in1(N__19263),
            .in2(_gnd_net_),
            .in3(N__43217),
            .lcout(G_535),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_13_16_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_13_16_4 .LUT_INIT=16'b0011001101000100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_13_16_4  (
            .in0(N__18300),
            .in1(N__18348),
            .in2(_gnd_net_),
            .in3(N__18446),
            .lcout(\this_vga_ramdac.N_24_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_13_16_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_13_16_5 .LUT_INIT=16'b0011001000111111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_13_16_5  (
            .in0(N__18448),
            .in1(N__18408),
            .in2(N__18355),
            .in3(N__18302),
            .lcout(),
            .ltout(\this_vga_ramdac.m6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_13_16_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_13_16_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_13_16_6 .LUT_INIT=16'b0010001000101110;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_13_16_6  (
            .in0(N__18249),
            .in1(N__20303),
            .in2(N__18256),
            .in3(N__26077),
            .lcout(\this_vga_ramdac.N_3857_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41999),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_9_LC_13_17_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_9_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_9_LC_13_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_9_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18238),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42006),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_RNIB85C3_LC_13_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIB85C3_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIB85C3_LC_13_17_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_RNIB85C3_LC_13_17_1  (
            .in0(N__22686),
            .in1(N__20341),
            .in2(_gnd_net_),
            .in3(N__27061),
            .lcout(),
            .ltout(\this_vga_signals.M_pcounter_q_ret_RNIB85CZ0Z3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNILVU44_1_LC_13_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNILVU44_1_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNILVU44_1_LC_13_17_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNILVU44_1_LC_13_17_2  (
            .in0(N__27280),
            .in1(_gnd_net_),
            .in2(N__18229),
            .in3(N__19327),
            .lcout(\this_vga_signals.N_3_0 ),
            .ltout(\this_vga_signals.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIOILK7_LC_13_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIOILK7_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIOILK7_LC_13_17_3 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_RNIOILK7_LC_13_17_3  (
            .in0(N__20366),
            .in1(_gnd_net_),
            .in2(N__18226),
            .in3(N__18196),
            .lcout(M_pcounter_q_ret_1_RNIOILK7),
            .ltout(M_pcounter_q_ret_1_RNIOILK7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_13_17_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_13_17_4 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_13_17_4  (
            .in0(N__18223),
            .in1(N__18207),
            .in2(N__18214),
            .in3(N__26074),
            .lcout(\this_vga_ramdac.N_3859_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42006),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIAI4F3_LC_13_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIAI4F3_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIAI4F3_LC_13_17_5 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_RNIAI4F3_LC_13_17_5  (
            .in0(N__20342),
            .in1(N__27279),
            .in2(N__20370),
            .in3(N__27062),
            .lcout(\this_vga_signals.N_2_0 ),
            .ltout(\this_vga_signals.N_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_13_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_13_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_13_17_6 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18538),
            .in3(N__22707),
            .lcout(\this_vga_signals.N_1417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42006),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_13_17_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_13_17_7 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_13_17_7  (
            .in0(N__26073),
            .in1(N__18535),
            .in2(N__18525),
            .in3(N__20306),
            .lcout(\this_vga_ramdac.N_3860_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42006),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_14_LC_13_18_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_14_LC_13_18_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_14_LC_13_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_14_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18508),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42017),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_0_LC_13_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_0_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_0_LC_13_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_0_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__18714),
            .in2(_gnd_net_),
            .in3(N__21916),
            .lcout(),
            .ltout(\this_ppu.m35_i_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_4_LC_13_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_4_LC_13_18_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_4_LC_13_18_2 .LUT_INIT=16'b0000000010110011;
    LogicCell40 \this_ppu.M_state_q_4_LC_13_18_2  (
            .in0(N__18730),
            .in1(N__21967),
            .in2(N__18496),
            .in3(N__26086),
            .lcout(\this_ppu.M_state_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42017),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNIUU07_9_LC_13_18_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNIUU07_9_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNIUU07_9_LC_13_18_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \this_ppu.oam_cache.read_data_RNIUU07_9_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__18493),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_oam_cache_read_data_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_11_LC_13_18_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_11_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_11_LC_13_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_11_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18487),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42017),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_1_LC_13_18_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_1_LC_13_18_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_1_LC_13_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_1_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18472),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42017),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNIA5M7_14_LC_13_18_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNIA5M7_14_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNIA5M7_14_LC_13_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNIA5M7_14_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18460),
            .lcout(\this_ppu.M_oam_cache_read_data_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_2_LC_13_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_2_LC_13_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_2_LC_13_18_7 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \this_ppu.M_state_q_2_LC_13_18_7  (
            .in0(N__18729),
            .in1(N__18715),
            .in2(N__43252),
            .in3(N__21917),
            .lcout(\this_ppu.M_state_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42017),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI94M7_13_LC_13_19_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI94M7_13_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI94M7_13_LC_13_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI94M7_13_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18691),
            .lcout(\this_ppu.M_oam_cache_read_data_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIRSG13_9_LC_13_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIRSG13_9_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIRSG13_9_LC_13_19_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIRSG13_9_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__27082),
            .in2(_gnd_net_),
            .in3(N__27312),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9 ),
            .ltout(\this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_19_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_19_2  (
            .in0(N__27313),
            .in1(_gnd_net_),
            .in2(N__18652),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.N_1307_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_8_LC_13_19_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_8_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_8_LC_13_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_8_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18643),
            .lcout(\this_ppu.M_oam_cache_read_data_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42026),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI72M7_11_LC_13_19_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI72M7_11_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI72M7_11_LC_13_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI72M7_11_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18628),
            .lcout(\this_ppu.M_oam_cache_read_data_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_o2_LC_13_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_o2_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_o2_LC_13_19_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m68_0_o2_LC_13_19_6  (
            .in0(N__21208),
            .in1(N__21145),
            .in2(N__21277),
            .in3(N__20437),
            .lcout(\this_ppu.N_82_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_0_LC_13_20_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_0_LC_13_20_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_0_LC_13_20_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \this_ppu.M_state_q_0_LC_13_20_1  (
            .in0(N__21592),
            .in1(N__26118),
            .in2(_gnd_net_),
            .in3(N__24615),
            .lcout(\this_ppu.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42034),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_0_LC_13_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_0_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_0_LC_13_20_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_0_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(N__18618),
            .in2(_gnd_net_),
            .in3(N__19220),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_1_LC_13_20_3 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_1_LC_13_20_3 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_1_LC_13_20_3 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clk.M_counter_q_1_LC_13_20_3  (
            .in0(N__19239),
            .in1(N__19267),
            .in2(_gnd_net_),
            .in3(N__43248),
            .lcout(this_pixel_clk_M_counter_q_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42034),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNII1437_3_LC_13_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNII1437_3_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNII1437_3_LC_13_20_4 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNII1437_3_LC_13_20_4  (
            .in0(N__19223),
            .in1(N__19152),
            .in2(N__19124),
            .in3(N__19034),
            .lcout(\this_vga_signals.M_hcounter_q_RNII1437Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_a3_1_0_LC_13_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_a3_1_0_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_a3_1_0_LC_13_20_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_a3_1_0_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__24250),
            .in2(_gnd_net_),
            .in3(N__30468),
            .lcout(\this_ppu.N_1182_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_ctle_7_LC_13_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_ctle_7_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_ctle_7_LC_13_20_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_ppu.M_screen_y_q_esr_ctle_7_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__26117),
            .in2(_gnd_net_),
            .in3(N__24614),
            .lcout(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_13_21_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_13_21_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_13_21_0  (
            .in0(N__24182),
            .in1(N__18979),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_3_LC_13_21_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_3_LC_13_21_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_3_LC_13_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_3_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18949),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42042),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_RNI8FJF7_4_LC_13_21_7 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_RNI8FJF7_4_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_RNI8FJF7_4_LC_13_21_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_RNI8FJF7_4_LC_13_21_7  (
            .in0(N__37330),
            .in1(N__39485),
            .in2(N__22474),
            .in3(N__37747),
            .lcout(\this_ppu.M_screen_y_q_RNI8FJF7Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_4_LC_13_22_0 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_4_LC_13_22_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_4_LC_13_22_0 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \this_ppu.M_surface_x_q_4_LC_13_22_0  (
            .in0(N__24678),
            .in1(N__22967),
            .in2(N__25822),
            .in3(N__23275),
            .lcout(M_this_ppu_map_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42053),
            .ce(),
            .sr(N__43114));
    defparam \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_13_22_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_13_22_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_13_22_1  (
            .in0(N__20200),
            .in1(N__38177),
            .in2(_gnd_net_),
            .in3(N__18934),
            .lcout(read_data_RNI5QFJ1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI62LG1_16_LC_13_22_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI62LG1_16_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI62LG1_16_LC_13_22_2 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI62LG1_16_LC_13_22_2  (
            .in0(N__38176),
            .in1(N__21572),
            .in2(_gnd_net_),
            .in3(N__20158),
            .lcout(M_this_ppu_spr_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_13_22_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_13_22_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_13_22_3  (
            .in0(N__19951),
            .in1(N__38175),
            .in2(_gnd_net_),
            .in3(N__41374),
            .lcout(read_data_RNI6RFJ1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_22_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_22_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_22_4  (
            .in0(N__38178),
            .in1(N__19723),
            .in2(_gnd_net_),
            .in3(N__43612),
            .lcout(read_data_RNI7SFJ1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_22_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_22_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_22_7  (
            .in0(N__19537),
            .in1(N__38174),
            .in2(_gnd_net_),
            .in3(N__43747),
            .lcout(read_data_RNI9TFJ1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_13_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_13_23_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_13_23_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_1_LC_13_23_0  (
            .in0(N__22693),
            .in1(N__20350),
            .in2(_gnd_net_),
            .in3(N__27101),
            .lcout(\this_vga_signals.M_pcounter_q_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42065),
            .ce(N__27335),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_11_LC_13_23_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_11_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_11_LC_13_23_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_11_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__19315),
            .in2(_gnd_net_),
            .in3(N__26735),
            .lcout(M_this_oam_ram_write_data_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_12_LC_13_23_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_12_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_12_LC_13_23_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_12_LC_13_23_3  (
            .in0(N__26736),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20239),
            .lcout(M_this_oam_ram_write_data_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_13_LC_13_23_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_13_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_13_LC_13_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_13_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__21598),
            .in2(_gnd_net_),
            .in3(N__26737),
            .lcout(M_this_oam_ram_write_data_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_14_LC_13_23_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_14_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_14_LC_13_23_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_14_LC_13_23_5  (
            .in0(N__26738),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20233),
            .lcout(M_this_oam_ram_write_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_12_LC_13_24_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_12_LC_13_24_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_12_LC_13_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_12_LC_13_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40763),
            .lcout(M_this_data_tmp_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42077),
            .ce(N__26559),
            .sr(N__43118));
    defparam M_this_data_tmp_q_esr_14_LC_13_24_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_14_LC_13_24_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_14_LC_13_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_14_LC_13_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40443),
            .lcout(M_this_data_tmp_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42077),
            .ce(N__26559),
            .sr(N__43118));
    defparam M_this_data_tmp_q_esr_1_LC_13_25_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_1_LC_13_25_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_1_LC_13_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_1_LC_13_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39686),
            .lcout(M_this_data_tmp_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42089),
            .ce(N__25668),
            .sr(N__43121));
    defparam M_this_data_tmp_q_esr_2_LC_13_25_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_2_LC_13_25_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_2_LC_13_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_2_LC_13_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42764),
            .lcout(M_this_data_tmp_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42089),
            .ce(N__25668),
            .sr(N__43121));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_22_LC_13_27_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_22_LC_13_27_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_22_LC_13_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_22_LC_13_27_0  (
            .in0(_gnd_net_),
            .in1(N__20206),
            .in2(_gnd_net_),
            .in3(N__26641),
            .lcout(M_this_oam_ram_write_data_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_22_LC_13_27_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_22_LC_13_27_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_22_LC_13_27_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 M_this_data_tmp_q_esr_22_LC_13_27_1 (
            .in0(_gnd_net_),
            .in1(N__40444),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42107),
            .ce(N__25633),
            .sr(N__43125));
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_1_LC_13_30_4 .C_ON=1'b0;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_1_LC_13_30_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_1_LC_13_30_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.IO_port_data_write_0_a2_i_1_LC_13_30_4  (
            .in0(_gnd_net_),
            .in1(N__43665),
            .in2(_gnd_net_),
            .in3(N__20199),
            .lcout(N_724_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_14_16_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_14_16_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_14_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20420),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41993),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_14_16_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_14_16_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_14_16_6  (
            .in0(N__20421),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20164),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41993),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_14_16_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_14_16_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__20422),
            .in2(_gnd_net_),
            .in3(N__20428),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41993),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_8_LC_14_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_8_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_8_LC_14_17_1 .LUT_INIT=16'b1000000011000100;
    LogicCell40 \this_ppu.M_state_q_8_LC_14_17_1  (
            .in0(N__23081),
            .in1(N__22129),
            .in2(N__21991),
            .in3(N__24430),
            .lcout(\this_ppu.M_state_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42000),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_14_17_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_14_17_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_14_17_4  (
            .in0(N__20412),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20380),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42000),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_0_LC_14_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_0_LC_14_17_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_0_LC_14_17_5 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_0_LC_14_17_5  (
            .in0(N__20346),
            .in1(N__27297),
            .in2(N__20371),
            .in3(N__27103),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42000),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_14_17_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_14_17_6 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_14_17_6  (
            .in0(N__20320),
            .in1(N__20305),
            .in2(N__20265),
            .in3(N__26076),
            .lcout(\this_vga_ramdac.N_3861_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42000),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNII6H51_6_LC_14_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNII6H51_6_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNII6H51_6_LC_14_17_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_RNII6H51_6_LC_14_17_7  (
            .in0(N__23818),
            .in1(N__23614),
            .in2(N__23083),
            .in3(N__22160),
            .lcout(\this_ppu.N_785_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_4_LC_14_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_4_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_4_LC_14_18_0 .LUT_INIT=16'b0111110010001100;
    LogicCell40 \this_ppu.M_screen_y_q_4_LC_14_18_0  (
            .in0(N__37259),
            .in1(N__37318),
            .in2(N__24682),
            .in3(N__37289),
            .lcout(\this_ppu.M_screen_y_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42007),
            .ce(),
            .sr(N__43107));
    defparam \this_ppu.M_screen_y_q_0_LC_14_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_0_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_0_LC_14_18_1 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \this_ppu.M_screen_y_q_0_LC_14_18_1  (
            .in0(N__24677),
            .in1(N__22384),
            .in2(N__22401),
            .in3(N__37260),
            .lcout(M_this_ppu_vram_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42007),
            .ce(),
            .sr(N__43107));
    defparam \this_ppu.M_surface_x_q_7_LC_14_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_7_LC_14_18_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_7_LC_14_18_2 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \this_ppu.M_surface_x_q_7_LC_14_18_2  (
            .in0(N__24668),
            .in1(N__21167),
            .in2(N__25780),
            .in3(N__20248),
            .lcout(M_this_ppu_map_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42007),
            .ce(),
            .sr(N__43107));
    defparam \this_ppu.M_surface_x_q_1_LC_14_18_3 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_1_LC_14_18_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_1_LC_14_18_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \this_ppu.M_surface_x_q_1_LC_14_18_3  (
            .in0(N__25753),
            .in1(N__24669),
            .in2(N__23317),
            .in3(N__23425),
            .lcout(\this_ppu.M_surface_x_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42007),
            .ce(),
            .sr(N__43107));
    defparam \this_ppu.M_surface_x_q_6_LC_14_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_6_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_6_LC_14_18_4 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \this_ppu.M_surface_x_q_6_LC_14_18_4  (
            .in0(N__24667),
            .in1(N__21238),
            .in2(N__25795),
            .in3(N__21940),
            .lcout(M_this_ppu_map_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42007),
            .ce(),
            .sr(N__43107));
    defparam \this_ppu.M_surface_x_q_0_LC_14_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_0_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_0_LC_14_18_5 .LUT_INIT=16'b1111000010011001;
    LogicCell40 \this_ppu.M_surface_x_q_0_LC_14_18_5  (
            .in0(N__23455),
            .in1(N__21963),
            .in2(N__25765),
            .in3(N__24674),
            .lcout(\this_ppu.offset_x ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42007),
            .ce(),
            .sr(N__43107));
    defparam \this_ppu.oam_cache.read_data_RNIB6J72_8_LC_14_18_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNIB6J72_8_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNIB6J72_8_LC_14_18_6 .LUT_INIT=16'b1011111000010100;
    LogicCell40 \this_ppu.oam_cache.read_data_RNIB6J72_8_LC_14_18_6  (
            .in0(N__38151),
            .in1(N__23453),
            .in2(N__20905),
            .in3(N__23454),
            .lcout(M_this_ppu_spr_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_3_LC_14_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_3_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_3_LC_14_18_7 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \this_ppu.M_surface_x_q_3_LC_14_18_7  (
            .in0(N__21949),
            .in1(N__24670),
            .in2(N__23400),
            .in3(N__25831),
            .lcout(M_this_ppu_map_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42007),
            .ce(),
            .sr(N__43107));
    defparam \this_ppu.offset_x_cry_0_c_inv_LC_14_19_0 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_0_c_inv_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_0_c_inv_LC_14_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.offset_x_cry_0_c_inv_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__20890),
            .in2(N__23467),
            .in3(N__20901),
            .lcout(\this_ppu.M_oam_cache_read_data_i_8 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\this_ppu.offset_x_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_0_c_RNI5N4U1_LC_14_19_1 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_0_c_RNI5N4U1_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_0_c_RNI5N4U1_LC_14_19_1 .LUT_INIT=16'b1110000110110100;
    LogicCell40 \this_ppu.offset_x_cry_0_c_RNI5N4U1_LC_14_19_1  (
            .in0(N__38150),
            .in1(N__20884),
            .in2(N__23316),
            .in3(N__20680),
            .lcout(M_this_ppu_spr_addr_1),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_0 ),
            .carryout(\this_ppu.offset_x_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_1_c_RNIFSQU1_LC_14_19_2 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_1_c_RNIFSQU1_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_1_c_RNIFSQU1_LC_14_19_2 .LUT_INIT=16'b1110000110110100;
    LogicCell40 \this_ppu.offset_x_cry_1_c_RNIFSQU1_LC_14_19_2  (
            .in0(N__38163),
            .in1(N__20677),
            .in2(N__23353),
            .in3(N__20446),
            .lcout(M_this_ppu_spr_addr_2),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_1 ),
            .carryout(\this_ppu.offset_x_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_o2_0_LC_14_19_3 .C_ON=1'b1;
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_o2_0_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_o2_0_LC_14_19_3 .LUT_INIT=16'b0001010001000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m68_0_o2_0_LC_14_19_3  (
            .in0(N__21292),
            .in1(N__20443),
            .in2(N__23397),
            .in3(N__20431),
            .lcout(\this_ppu.m68_0_o2_0 ),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_2 ),
            .carryout(\this_ppu.offset_x_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_3_c_RNI3UBP_LC_14_19_4 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_3_c_RNI3UBP_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_3_c_RNI3UBP_LC_14_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.offset_x_cry_3_c_RNI3UBP_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__21301),
            .in2(N__22997),
            .in3(N__21286),
            .lcout(\this_ppu.offset_x_4 ),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_3 ),
            .carryout(\this_ppu.offset_x_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_4_c_RNI62DP_LC_14_19_5 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_4_c_RNI62DP_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_4_c_RNI62DP_LC_14_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.offset_x_cry_4_c_RNI62DP_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__21283),
            .in2(N__22914),
            .in3(N__21268),
            .lcout(\this_ppu.offset_x_5 ),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_4 ),
            .carryout(\this_ppu.offset_x_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_5_c_RNI96EP_LC_14_19_6 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_5_c_RNI96EP_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_5_c_RNI96EP_LC_14_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.offset_x_cry_5_c_RNI96EP_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__21265),
            .in2(N__21242),
            .in3(N__21202),
            .lcout(\this_ppu.offset_x_6 ),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_5 ),
            .carryout(\this_ppu.offset_x_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_6_c_THRU_CRY_0_LC_14_19_7 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_6_c_THRU_CRY_0_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_6_c_THRU_CRY_0_LC_14_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.offset_x_cry_6_c_THRU_CRY_0_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__24933),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_6 ),
            .carryout(\this_ppu.offset_x_cry_6_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_6_c_RNICAFP_LC_14_20_0 .C_ON=1'b0;
    defparam \this_ppu.offset_x_cry_6_c_RNICAFP_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_6_c_RNICAFP_LC_14_20_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_ppu.offset_x_cry_6_c_RNICAFP_LC_14_20_0  (
            .in0(N__21199),
            .in1(N__21171),
            .in2(_gnd_net_),
            .in3(N__21148),
            .lcout(\this_ppu.offset_x_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNI453Q6_1_LC_14_20_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNI453Q6_1_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNI453Q6_1_LC_14_20_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNI453Q6_1_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__22079),
            .in2(_gnd_net_),
            .in3(N__37237),
            .lcout(\this_ppu.M_screen_y_q_esr_RNI453Q6Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNII6H51_1_LC_14_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNII6H51_1_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNII6H51_1_LC_14_20_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_RNII6H51_1_LC_14_20_3  (
            .in0(N__23064),
            .in1(N__21918),
            .in2(N__23671),
            .in3(N__23610),
            .lcout(\this_ppu.un30_0_a2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIJ1SE_10_LC_14_20_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIJ1SE_10_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIJ1SE_10_LC_14_20_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_state_q_RNIJ1SE_10_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__23200),
            .in2(_gnd_net_),
            .in3(N__22164),
            .lcout(\this_ppu.N_999_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_i_1_LC_14_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_i_1_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_i_1_LC_14_20_7 .LUT_INIT=16'b0001011000010000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m13_0_i_1_LC_14_20_7  (
            .in0(N__22165),
            .in1(N__23202),
            .in2(N__24263),
            .in3(N__24422),
            .lcout(\this_ppu.m13_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CRY_0_LC_14_21_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CRY_0_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CRY_0_LC_14_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CRY_0_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__37238),
            .in2(N__37255),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_y_q_esr_0_LC_14_21_1 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_0_LC_14_21_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_0_LC_14_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_0_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__22345),
            .in2(N__22207),
            .in3(N__21550),
            .lcout(\this_ppu.offset_y ),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_0 ),
            .clk(N__42035),
            .ce(N__37169),
            .sr(N__43110));
    defparam \this_ppu.M_surface_y_q_esr_1_LC_14_21_2 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_1_LC_14_21_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_1_LC_14_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_1_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__21547),
            .in2(N__22198),
            .in3(N__21511),
            .lcout(\this_ppu.M_surface_y_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_0 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_1 ),
            .clk(N__42035),
            .ce(N__37169),
            .sr(N__43110));
    defparam \this_ppu.M_surface_y_q_esr_2_LC_14_21_3 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_2_LC_14_21_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_2_LC_14_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_2_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__21685),
            .in2(N__22483),
            .in3(N__21478),
            .lcout(\this_ppu.M_surface_y_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_1 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_2 ),
            .clk(N__42035),
            .ce(N__37169),
            .sr(N__43110));
    defparam \this_ppu.M_surface_y_q_esr_3_LC_14_21_4 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_3_LC_14_21_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_3_LC_14_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_3_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__23680),
            .in2(N__23697),
            .in3(N__21436),
            .lcout(M_this_ppu_map_addr_5),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_2 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_3 ),
            .clk(N__42035),
            .ce(N__37169),
            .sr(N__43110));
    defparam \this_ppu.M_surface_y_q_esr_4_LC_14_21_5 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_4_LC_14_21_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_4_LC_14_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_4_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__21433),
            .in2(N__22470),
            .in3(N__21391),
            .lcout(M_this_ppu_map_addr_6),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_3 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_4 ),
            .clk(N__42035),
            .ce(N__37169),
            .sr(N__43110));
    defparam \this_ppu.M_surface_y_q_esr_5_LC_14_21_6 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_5_LC_14_21_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_5_LC_14_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_5_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__37060),
            .in2(N__37086),
            .in3(N__21346),
            .lcout(M_this_ppu_map_addr_7),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_4 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_5 ),
            .clk(N__42035),
            .ce(N__37169),
            .sr(N__43110));
    defparam \this_ppu.M_surface_y_q_esr_6_LC_14_21_7 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_6_LC_14_21_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_6_LC_14_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_6_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__34597),
            .in2(N__34614),
            .in3(N__21304),
            .lcout(M_this_ppu_map_addr_8),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_5 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_6 ),
            .clk(N__42035),
            .ce(N__37169),
            .sr(N__43110));
    defparam \this_ppu.M_surface_y_q_esr_7_LC_14_22_0 .C_ON=1'b0;
    defparam \this_ppu.M_surface_y_q_esr_7_LC_14_22_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_7_LC_14_22_0 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \this_ppu.M_surface_y_q_esr_7_LC_14_22_0  (
            .in0(N__22447),
            .in1(N__37254),
            .in2(N__22102),
            .in3(N__21727),
            .lcout(M_this_ppu_map_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42043),
            .ce(N__37176),
            .sr(N__43113));
    defparam \this_ppu.M_screen_y_q_esr_1_LC_14_22_2 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_1_LC_14_22_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_1_LC_14_22_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_1_LC_14_22_2  (
            .in0(N__22080),
            .in1(N__22403),
            .in2(_gnd_net_),
            .in3(N__37253),
            .lcout(\this_ppu.M_screen_y_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42043),
            .ce(N__37176),
            .sr(N__43113));
    defparam \this_ppu.M_screen_y_q_esr_2_LC_14_22_3 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_2_LC_14_22_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_2_LC_14_22_3 .LUT_INIT=16'b0010100010100000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_2_LC_14_22_3  (
            .in0(N__37251),
            .in1(N__22081),
            .in2(N__22030),
            .in3(N__22404),
            .lcout(\this_ppu.M_screen_y_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42043),
            .ce(N__37176),
            .sr(N__43113));
    defparam \this_ppu.M_screen_y_q_esr_RNI563Q6_2_LC_14_22_4 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNI563Q6_2_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNI563Q6_2_LC_14_22_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNI563Q6_2_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__22025),
            .in2(_gnd_net_),
            .in3(N__37250),
            .lcout(\this_ppu.M_screen_y_q_esr_RNI563Q6Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_3_LC_14_22_5 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_3_LC_14_22_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_3_LC_14_22_5 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_3_LC_14_22_5  (
            .in0(N__37252),
            .in1(N__23736),
            .in2(N__22009),
            .in3(N__22054),
            .lcout(\this_ppu.M_screen_y_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42043),
            .ce(N__37176),
            .sr(N__43113));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_14_22_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_14_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_14_22_6  (
            .in0(N__24179),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21676),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_14_22_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_14_22_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(N__24178),
            .in2(_gnd_net_),
            .in3(N__21640),
            .lcout(\this_ppu.oam_cache.N_581_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_13_LC_14_23_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_13_LC_14_23_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_13_LC_14_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_13_LC_14_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40069),
            .lcout(M_this_data_tmp_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42054),
            .ce(N__26558),
            .sr(N__43115));
    defparam M_this_data_count_q_cry_c_0_LC_14_24_0.C_ON=1'b1;
    defparam M_this_data_count_q_cry_c_0_LC_14_24_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_c_0_LC_14_24_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 M_this_data_count_q_cry_c_0_LC_14_24_0 (
            .in0(_gnd_net_),
            .in1(N__22426),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(M_this_data_count_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_14_24_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_14_24_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_14_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_0_THRU_LUT4_0_LC_14_24_1 (
            .in0(_gnd_net_),
            .in1(N__22588),
            .in2(N__25018),
            .in3(N__21754),
            .lcout(M_this_data_count_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_0),
            .carryout(M_this_data_count_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_14_24_2.C_ON=1'b1;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_14_24_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_14_24_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_1_THRU_LUT4_0_LC_14_24_2 (
            .in0(_gnd_net_),
            .in1(N__24950),
            .in2(N__22567),
            .in3(N__21751),
            .lcout(M_this_data_count_q_cry_1_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_1),
            .carryout(M_this_data_count_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_14_24_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_14_24_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_14_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_2_THRU_LUT4_0_LC_14_24_3 (
            .in0(_gnd_net_),
            .in1(N__22541),
            .in2(N__25019),
            .in3(N__21748),
            .lcout(M_this_data_count_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_2),
            .carryout(M_this_data_count_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_14_24_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_14_24_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_14_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_3_THRU_LUT4_0_LC_14_24_4 (
            .in0(_gnd_net_),
            .in1(N__24954),
            .in2(N__22747),
            .in3(N__21745),
            .lcout(M_this_data_count_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_3),
            .carryout(M_this_data_count_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_14_24_5.C_ON=1'b1;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_14_24_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_14_24_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_4_THRU_LUT4_0_LC_14_24_5 (
            .in0(_gnd_net_),
            .in1(N__22764),
            .in2(N__25020),
            .in3(N__21742),
            .lcout(M_this_data_count_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_4),
            .carryout(M_this_data_count_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_14_24_6.C_ON=1'b1;
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_14_24_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_14_24_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_5_THRU_LUT4_0_LC_14_24_6 (
            .in0(_gnd_net_),
            .in1(N__24958),
            .in2(N__25717),
            .in3(N__21739),
            .lcout(M_this_data_count_q_cry_5_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_5),
            .carryout(M_this_data_count_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_14_24_7.C_ON=1'b1;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_14_24_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_14_24_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_6_THRU_LUT4_0_LC_14_24_7 (
            .in0(_gnd_net_),
            .in1(N__25741),
            .in2(N__25021),
            .in3(N__21736),
            .lcout(M_this_data_count_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_6),
            .carryout(M_this_data_count_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_8_LC_14_25_0.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_8_LC_14_25_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_8_LC_14_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_8_LC_14_25_0 (
            .in0(_gnd_net_),
            .in1(N__22777),
            .in2(N__24887),
            .in3(N__21733),
            .lcout(M_this_data_count_q_s_8),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(M_this_data_count_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_14_25_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_14_25_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_14_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_8_THRU_LUT4_0_LC_14_25_1 (
            .in0(_gnd_net_),
            .in1(N__25390),
            .in2(N__24890),
            .in3(N__21730),
            .lcout(M_this_data_count_q_cry_8_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_8),
            .carryout(M_this_data_count_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_10_LC_14_25_2.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_10_LC_14_25_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_10_LC_14_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_10_LC_14_25_2 (
            .in0(_gnd_net_),
            .in1(N__22795),
            .in2(N__24886),
            .in3(N__21826),
            .lcout(M_this_data_count_q_s_10),
            .ltout(),
            .carryin(M_this_data_count_q_cry_9),
            .carryout(M_this_data_count_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_14_25_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_14_25_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_14_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_10_THRU_LUT4_0_LC_14_25_3 (
            .in0(_gnd_net_),
            .in1(N__22825),
            .in2(N__24889),
            .in3(N__21823),
            .lcout(M_this_data_count_q_cry_10_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_10),
            .carryout(M_this_data_count_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_14_25_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_14_25_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_14_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_11_THRU_LUT4_0_LC_14_25_4 (
            .in0(_gnd_net_),
            .in1(N__22842),
            .in2(N__24888),
            .in3(N__21820),
            .lcout(M_this_data_count_q_cry_11_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_11),
            .carryout(M_this_data_count_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_13_LC_14_25_5.C_ON=1'b0;
    defparam M_this_data_count_q_RNO_0_13_LC_14_25_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_13_LC_14_25_5.LUT_INIT=16'b1100110000110011;
    LogicCell40 M_this_data_count_q_RNO_0_13_LC_14_25_5 (
            .in0(_gnd_net_),
            .in1(N__22809),
            .in2(_gnd_net_),
            .in3(N__21817),
            .lcout(M_this_data_count_q_s_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_7_LC_14_26_5.C_ON=1'b0;
    defparam M_this_oam_address_q_7_LC_14_26_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_7_LC_14_26_5.LUT_INIT=16'b0001001000110000;
    LogicCell40 M_this_oam_address_q_7_LC_14_26_5 (
            .in0(N__26457),
            .in1(N__27489),
            .in2(N__21807),
            .in3(N__22726),
            .lcout(M_this_oam_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42090),
            .ce(),
            .sr(N__41640));
    defparam \this_vga_signals.IO_port_data_write_i_m2_i_m2_0_LC_14_27_0 .C_ON=1'b0;
    defparam \this_vga_signals.IO_port_data_write_i_m2_i_m2_0_LC_14_27_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.IO_port_data_write_i_m2_i_m2_0_LC_14_27_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vga_signals.IO_port_data_write_i_m2_i_m2_0_LC_14_27_0  (
            .in0(N__38233),
            .in1(N__43664),
            .in2(_gnd_net_),
            .in3(N__21878),
            .lcout(IO_port_data_write_i_m2_i_m2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_15_15_5.C_ON=1'b0;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_15_15_5.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_15_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_15_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43218),
            .lcout(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m48_i_0_a3_0_LC_15_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m48_i_0_a3_0_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m48_i_0_a3_0_LC_15_17_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m48_i_0_a3_0_LC_15_17_2  (
            .in0(N__40479),
            .in1(N__22180),
            .in2(_gnd_net_),
            .in3(N__24423),
            .lcout(\this_ppu.N_1202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_9_LC_15_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_9_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_9_LC_15_17_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_state_q_9_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__21760),
            .in2(_gnd_net_),
            .in3(N__43242),
            .lcout(\this_ppu.M_state_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41994),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIU3I91_3_LC_15_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIU3I91_3_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIU3I91_3_LC_15_18_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIU3I91_3_LC_15_18_2  (
            .in0(N__23172),
            .in1(N__23751),
            .in2(_gnd_net_),
            .in3(N__34454),
            .lcout(\this_ppu.N_1426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_6_LC_15_18_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_6_LC_15_18_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_6_LC_15_18_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_ppu.M_state_q_6_LC_15_18_3  (
            .in0(N__21987),
            .in1(N__23074),
            .in2(_gnd_net_),
            .in3(N__43244),
            .lcout(\this_ppu.M_state_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42001),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_o3_LC_15_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_o3_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_0_o3_LC_15_18_4 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m35_i_0_o3_LC_15_18_4  (
            .in0(N__23609),
            .in1(N__34368),
            .in2(_gnd_net_),
            .in3(N__23653),
            .lcout(\this_ppu.N_91_0 ),
            .ltout(\this_ppu.N_91_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_RNIN4DCD_1_LC_15_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNIN4DCD_1_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNIN4DCD_1_LC_15_18_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNIN4DCD_1_LC_15_18_5  (
            .in0(N__23346),
            .in1(N__23312),
            .in2(N__21952),
            .in3(N__23461),
            .lcout(\this_ppu.un1_M_surface_x_q_c3 ),
            .ltout(\this_ppu.un1_M_surface_x_q_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_RNO_0_6_LC_15_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNO_0_6_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNO_0_6_LC_15_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNO_0_6_LC_15_18_6  (
            .in0(N__22887),
            .in1(N__22986),
            .in2(N__21943),
            .in3(N__23390),
            .lcout(\this_ppu.un1_M_surface_x_q_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_5_LC_15_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_5_LC_15_19_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_5_LC_15_19_0 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \this_ppu.M_state_q_5_LC_15_19_0  (
            .in0(N__26129),
            .in1(N__21832),
            .in2(N__21934),
            .in3(N__22116),
            .lcout(\this_ppu.M_state_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42008),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIRJK11_1_LC_15_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIRJK11_1_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIRJK11_1_LC_15_19_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_RNIRJK11_1_LC_15_19_2  (
            .in0(N__21922),
            .in1(N__23665),
            .in2(N__24176),
            .in3(N__24218),
            .lcout(\this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_10_LC_15_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_10_LC_15_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_10_LC_15_19_3 .LUT_INIT=16'b0010001100100010;
    LogicCell40 \this_ppu.M_state_q_10_LC_15_19_3  (
            .in0(N__24219),
            .in1(N__26130),
            .in2(N__21889),
            .in3(N__24681),
            .lcout(\this_ppu.M_state_qZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42008),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m48_i_0_a3_LC_15_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m48_i_0_a3_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m48_i_0_a3_LC_15_19_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m48_i_0_a3_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__23822),
            .in2(_gnd_net_),
            .in3(N__23793),
            .lcout(\this_ppu.N_1201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_8_LC_15_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_8_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_8_LC_15_19_6 .LUT_INIT=16'b0000000000100110;
    LogicCell40 \this_ppu.M_state_q_RNO_0_8_LC_15_19_6  (
            .in0(N__23073),
            .in1(N__22181),
            .in2(N__40480),
            .in3(N__43233),
            .lcout(\this_ppu.M_state_q_srsts_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNII1FQB_7_LC_15_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNII1FQB_7_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNII1FQB_7_LC_15_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_state_q_RNII1FQB_7_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__23596),
            .in2(_gnd_net_),
            .in3(N__34374),
            .lcout(\this_ppu.N_1145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_7_LC_15_20_0 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_7_LC_15_20_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_7_LC_15_20_0 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_7_LC_15_20_0  (
            .in0(N__37236),
            .in1(N__36594),
            .in2(N__22098),
            .in3(N__22039),
            .lcout(\this_ppu.M_screen_y_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42018),
            .ce(N__37165),
            .sr(N__43108));
    defparam \this_ppu.M_screen_y_q_esr_RNIQ8BT6_1_LC_15_20_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIQ8BT6_1_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIQ8BT6_1_LC_15_20_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIQ8BT6_1_LC_15_20_1  (
            .in0(N__22078),
            .in1(N__22394),
            .in2(_gnd_net_),
            .in3(N__37234),
            .lcout(\this_ppu.un3_M_screen_y_d_0_c2 ),
            .ltout(\this_ppu.un3_M_screen_y_d_0_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNI5MHHK_3_LC_15_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNI5MHHK_3_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNI5MHHK_3_LC_15_20_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNI5MHHK_3_LC_15_20_2  (
            .in0(N__37235),
            .in1(N__23750),
            .in2(N__22045),
            .in3(N__22002),
            .lcout(\this_ppu.un3_M_screen_y_d_0_c4 ),
            .ltout(\this_ppu.un3_M_screen_y_d_0_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNO_0_7_LC_15_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNO_0_7_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNO_0_7_LC_15_20_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNO_0_7_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__37135),
            .in2(N__22042),
            .in3(N__37329),
            .lcout(\this_ppu.un3_M_screen_y_d_0_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI467N6_8_LC_15_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI467N6_8_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI467N6_8_LC_15_20_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI467N6_8_LC_15_20_4  (
            .in0(N__26368),
            .in1(N__37730),
            .in2(_gnd_net_),
            .in3(N__28038),
            .lcout(N_861_0),
            .ltout(N_861_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNI563Q6_0_2_LC_15_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNI563Q6_0_2_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNI563Q6_0_2_LC_15_20_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNI563Q6_0_2_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22033),
            .in3(N__22029),
            .lcout(\this_ppu.un3_M_screen_y_d_a_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_2_LC_15_21_0 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_2_LC_15_21_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_2_LC_15_21_0 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \this_ppu.M_screen_x_q_2_LC_15_21_0  (
            .in0(N__24665),
            .in1(N__26131),
            .in2(N__22233),
            .in3(N__23481),
            .lcout(M_this_ppu_vram_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42027),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_RNIQ9FQ6_0_LC_15_21_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_RNIQ9FQ6_0_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_RNIQ9FQ6_0_LC_15_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_screen_y_q_RNIQ9FQ6_0_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__22402),
            .in2(_gnd_net_),
            .in3(N__37233),
            .lcout(\this_ppu.M_screen_y_q_RNIQ9FQ6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_RNI5A3DD_2_LC_15_21_2 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_RNI5A3DD_2_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_x_q_RNI5A3DD_2_LC_15_21_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_screen_x_q_RNI5A3DD_2_LC_15_21_2  (
            .in0(N__22224),
            .in1(N__23156),
            .in2(_gnd_net_),
            .in3(N__23479),
            .lcout(\this_ppu.un1_M_screen_x_q_c4 ),
            .ltout(\this_ppu.un1_M_screen_x_q_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_4_LC_15_21_3 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_4_LC_15_21_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_4_LC_15_21_3 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \this_ppu.M_screen_x_q_4_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__22313),
            .in2(N__22339),
            .in3(N__23769),
            .lcout(M_this_ppu_vram_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42027),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_5_LC_15_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_5_LC_15_21_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_5_LC_15_21_4 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \this_ppu.M_screen_x_q_5_LC_15_21_4  (
            .in0(N__23771),
            .in1(N__22281),
            .in2(N__22320),
            .in3(N__22336),
            .lcout(M_this_ppu_vram_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42027),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_RNO_0_6_LC_15_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_RNO_0_6_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_x_q_RNO_0_6_LC_15_21_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_screen_x_q_RNO_0_6_LC_15_21_5  (
            .in0(N__23480),
            .in1(N__22225),
            .in2(N__23170),
            .in3(N__22312),
            .lcout(),
            .ltout(\this_ppu.un1_M_screen_x_q_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_6_LC_15_21_6 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_6_LC_15_21_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_6_LC_15_21_6 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \this_ppu.M_screen_x_q_6_LC_15_21_6  (
            .in0(N__23772),
            .in1(N__22254),
            .in2(N__22297),
            .in3(N__22280),
            .lcout(M_this_ppu_vram_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42027),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_3_LC_15_21_7 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_3_LC_15_21_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_3_LC_15_21_7 .LUT_INIT=16'b0111100000000000;
    LogicCell40 \this_ppu.M_screen_x_q_3_LC_15_21_7  (
            .in0(N__23482),
            .in1(N__22229),
            .in2(N__23171),
            .in3(N__23770),
            .lcout(M_this_ppu_vram_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42027),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_scroll_q_esr_0_LC_15_22_0.C_ON=1'b0;
    defparam M_this_scroll_q_esr_0_LC_15_22_0.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_0_LC_15_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_0_LC_15_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42439),
            .lcout(M_this_scroll_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42036),
            .ce(N__26341),
            .sr(N__43111));
    defparam M_this_scroll_q_esr_1_LC_15_22_1.C_ON=1'b0;
    defparam M_this_scroll_q_esr_1_LC_15_22_1.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_1_LC_15_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_1_LC_15_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39753),
            .lcout(M_this_scroll_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42036),
            .ce(N__26341),
            .sr(N__43111));
    defparam M_this_scroll_q_esr_2_LC_15_22_2.C_ON=1'b0;
    defparam M_this_scroll_q_esr_2_LC_15_22_2.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_2_LC_15_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_2_LC_15_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42765),
            .lcout(M_this_scroll_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42036),
            .ce(N__26341),
            .sr(N__43111));
    defparam M_this_scroll_q_esr_3_LC_15_22_3.C_ON=1'b0;
    defparam M_this_scroll_q_esr_3_LC_15_22_3.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_3_LC_15_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_3_LC_15_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41514),
            .lcout(M_this_scroll_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42036),
            .ce(N__26341),
            .sr(N__43111));
    defparam M_this_scroll_q_esr_4_LC_15_22_4.C_ON=1'b0;
    defparam M_this_scroll_q_esr_4_LC_15_22_4.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_4_LC_15_22_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_4_LC_15_22_4 (
            .in0(N__40784),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42036),
            .ce(N__26341),
            .sr(N__43111));
    defparam M_this_scroll_q_esr_5_LC_15_22_5.C_ON=1'b0;
    defparam M_this_scroll_q_esr_5_LC_15_22_5.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_5_LC_15_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_5_LC_15_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40068),
            .lcout(M_this_scroll_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42036),
            .ce(N__26341),
            .sr(N__43111));
    defparam M_this_scroll_q_esr_6_LC_15_22_6.C_ON=1'b0;
    defparam M_this_scroll_q_esr_6_LC_15_22_6.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_6_LC_15_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_6_LC_15_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40411),
            .lcout(M_this_scroll_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42036),
            .ce(N__26341),
            .sr(N__43111));
    defparam M_this_scroll_q_esr_7_LC_15_22_7.C_ON=1'b0;
    defparam M_this_scroll_q_esr_7_LC_15_22_7.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_7_LC_15_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_7_LC_15_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39856),
            .lcout(M_this_scroll_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42036),
            .ce(N__26341),
            .sr(N__43111));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_15_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_15_23_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_15_23_0  (
            .in0(N__27853),
            .in1(N__27397),
            .in2(N__34768),
            .in3(N__35012),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_12_LC_15_23_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_12_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_12_LC_15_23_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_o2_12_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__43470),
            .in2(_gnd_net_),
            .in3(N__29285),
            .lcout(N_1005_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_9_16_LC_15_24_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_9_16_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_9_16_LC_15_24_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_9_16_LC_15_24_0  (
            .in0(N__22562),
            .in1(N__22586),
            .in2(N__22542),
            .in3(N__22424),
            .lcout(\this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_0_LC_15_24_1.C_ON=1'b0;
    defparam M_this_data_count_q_0_LC_15_24_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_15_24_1.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_0_LC_15_24_1 (
            .in0(N__22425),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27537),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42055),
            .ce(N__25358),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_1_LC_15_24_2.C_ON=1'b0;
    defparam M_this_data_count_q_1_LC_15_24_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_15_24_2.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_1_LC_15_24_2 (
            .in0(N__27538),
            .in1(N__22594),
            .in2(_gnd_net_),
            .in3(N__22587),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42055),
            .ce(N__25358),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_2_LC_15_24_3.C_ON=1'b0;
    defparam M_this_data_count_q_2_LC_15_24_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_15_24_3.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_2_LC_15_24_3 (
            .in0(N__22573),
            .in1(N__22563),
            .in2(_gnd_net_),
            .in3(N__27539),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42055),
            .ce(N__25358),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_3_LC_15_24_4.C_ON=1'b0;
    defparam M_this_data_count_q_3_LC_15_24_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_15_24_4.LUT_INIT=16'b0101000000000101;
    LogicCell40 M_this_data_count_q_3_LC_15_24_4 (
            .in0(N__27540),
            .in1(_gnd_net_),
            .in2(N__22543),
            .in3(N__22549),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42055),
            .ce(N__25358),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_4_LC_15_24_5.C_ON=1'b0;
    defparam M_this_data_count_q_4_LC_15_24_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_15_24_5.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_4_LC_15_24_5 (
            .in0(N__22522),
            .in1(N__27541),
            .in2(_gnd_net_),
            .in3(N__22746),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42055),
            .ce(N__25358),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_5_LC_15_24_6.C_ON=1'b0;
    defparam M_this_data_count_q_5_LC_15_24_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_15_24_6.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_5_LC_15_24_6 (
            .in0(N__27542),
            .in1(N__22516),
            .in2(_gnd_net_),
            .in3(N__22765),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42055),
            .ce(N__25358),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_6_LC_15_24_7.C_ON=1'b0;
    defparam M_this_data_count_q_6_LC_15_24_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_15_24_7.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_6_LC_15_24_7 (
            .in0(N__22510),
            .in1(N__25715),
            .in2(_gnd_net_),
            .in3(N__27543),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42055),
            .ce(N__25358),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_11_LC_15_25_1.C_ON=1'b0;
    defparam M_this_data_count_q_11_LC_15_25_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_15_25_1.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_11_LC_15_25_1 (
            .in0(N__27545),
            .in1(N__22504),
            .in2(_gnd_net_),
            .in3(N__22824),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42066),
            .ce(N__25366),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_10_LC_15_25_2.C_ON=1'b0;
    defparam M_this_data_count_q_10_LC_15_25_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_15_25_2.LUT_INIT=16'b1110001000100010;
    LogicCell40 M_this_data_count_q_10_LC_15_25_2 (
            .in0(N__22498),
            .in1(N__27544),
            .in2(N__43529),
            .in3(N__28138),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42066),
            .ce(N__25366),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_12_LC_15_25_3.C_ON=1'b0;
    defparam M_this_data_count_q_12_LC_15_25_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_15_25_3.LUT_INIT=16'b0101000000000101;
    LogicCell40 M_this_data_count_q_12_LC_15_25_3 (
            .in0(N__27546),
            .in1(_gnd_net_),
            .in2(N__22843),
            .in3(N__22489),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42066),
            .ce(N__25366),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_15_25_4.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_15_25_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_15_25_4.LUT_INIT=16'b0010001011100010;
    LogicCell40 M_this_data_count_q_13_LC_15_25_4 (
            .in0(N__22852),
            .in1(N__27547),
            .in2(N__33170),
            .in3(N__43249),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42066),
            .ce(N__25366),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_16_LC_15_25_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_16_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_16_LC_15_25_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_8_16_LC_15_25_5  (
            .in0(N__22838),
            .in1(N__22823),
            .in2(N__22810),
            .in3(N__22794),
            .lcout(\this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_8_LC_15_25_6.C_ON=1'b0;
    defparam M_this_data_count_q_8_LC_15_25_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_15_25_6.LUT_INIT=16'b0010001011100010;
    LogicCell40 M_this_data_count_q_8_LC_15_25_6 (
            .in0(N__22783),
            .in1(N__27548),
            .in2(N__27490),
            .in3(N__43250),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42066),
            .ce(N__25366),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_7_16_LC_15_25_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_7_16_LC_15_25_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_7_16_LC_15_25_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_7_16_LC_15_25_7  (
            .in0(N__22776),
            .in1(N__22763),
            .in2(N__25389),
            .in3(N__22742),
            .lcout(\this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNO_0_7_LC_15_26_2.C_ON=1'b0;
    defparam M_this_oam_address_q_RNO_0_7_LC_15_26_2.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNO_0_7_LC_15_26_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_oam_address_q_RNO_0_7_LC_15_26_2 (
            .in0(N__26923),
            .in1(N__26988),
            .in2(N__26514),
            .in3(N__26943),
            .lcout(un1_M_this_oam_address_q_c6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3SF72_9_LC_16_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3SF72_9_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3SF72_9_LC_16_16_5 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3SF72_9_LC_16_16_5  (
            .in0(N__30541),
            .in1(N__22720),
            .in2(_gnd_net_),
            .in3(N__30589),
            .lcout(\this_vga_signals.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_LC_16_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_16_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_16_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22708),
            .lcout(\this_vga_signals.M_pcounter_q_i_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41990),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_cache_cnt_q_2_LC_16_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_oam_cache_cnt_q_2_LC_16_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_cache_cnt_q_2_LC_16_17_2 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \this_ppu.M_oam_cache_cnt_q_2_LC_16_17_2  (
            .in0(N__22669),
            .in1(N__43236),
            .in2(N__22636),
            .in3(N__24666),
            .lcout(\this_ppu.M_oam_cache_cnt_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41990),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_16_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_16_17_3 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_0_LC_16_17_3  (
            .in0(N__30467),
            .in1(_gnd_net_),
            .in2(N__25891),
            .in3(N__25968),
            .lcout(),
            .ltout(\this_vga_signals.M_lcounter_q_e_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_0_LC_16_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_0_LC_16_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_0_LC_16_17_4 .LUT_INIT=16'b0110001010101010;
    LogicCell40 \this_vga_signals.M_lcounter_q_0_LC_16_17_4  (
            .in0(N__25932),
            .in1(N__27334),
            .in2(N__23038),
            .in3(N__27102),
            .lcout(this_vga_signals_M_lcounter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41990),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_2_LC_16_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_2_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_2_LC_16_17_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_o2_2_LC_16_17_7  (
            .in0(N__25887),
            .in1(N__25931),
            .in2(_gnd_net_),
            .in3(N__25855),
            .lcout(\this_ppu.N_838_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNICH7OC_11_LC_16_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNICH7OC_11_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNICH7OC_11_LC_16_18_0 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \this_ppu.M_state_q_RNICH7OC_11_LC_16_18_0  (
            .in0(N__24220),
            .in1(N__23658),
            .in2(N__39952),
            .in3(N__23017),
            .lcout(N_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNII1FQB_0_7_LC_16_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNII1FQB_0_7_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNII1FQB_0_7_LC_16_18_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_ppu.M_state_q_RNII1FQB_0_7_LC_16_18_1  (
            .in0(N__23611),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34369),
            .lcout(\this_ppu.N_1198 ),
            .ltout(\this_ppu.N_1198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_RNINHSUC_1_LC_16_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNINHSUC_1_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNINHSUC_1_LC_16_18_2 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNINHSUC_1_LC_16_18_2  (
            .in0(N__23311),
            .in1(N__23657),
            .in2(N__23011),
            .in3(N__23466),
            .lcout(\this_ppu.un1_M_surface_x_q_c2 ),
            .ltout(\this_ppu.un1_M_surface_x_q_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_RNO_0_5_LC_16_18_3 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNO_0_5_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNO_0_5_LC_16_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNO_0_5_LC_16_18_3  (
            .in0(N__23399),
            .in1(N__22987),
            .in2(N__22930),
            .in3(N__23344),
            .lcout(),
            .ltout(\this_ppu.un1_M_surface_x_q_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_5_LC_16_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_5_LC_16_18_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_5_LC_16_18_4 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \this_ppu.M_surface_x_q_5_LC_16_18_4  (
            .in0(N__24675),
            .in1(N__25804),
            .in2(N__22927),
            .in3(N__22888),
            .lcout(M_this_ppu_map_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41991),
            .ce(),
            .sr(N__43105));
    defparam \this_ppu.M_surface_x_q_2_LC_16_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_2_LC_16_18_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_2_LC_16_18_5 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \this_ppu.M_surface_x_q_2_LC_16_18_5  (
            .in0(N__22858),
            .in1(N__24676),
            .in2(N__25840),
            .in3(N__23345),
            .lcout(\this_ppu.M_surface_x_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41991),
            .ce(),
            .sr(N__43105));
    defparam \this_ppu.M_state_q_RNIOVBHC_9_LC_16_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIOVBHC_9_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIOVBHC_9_LC_16_18_6 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \this_ppu.M_state_q_RNIOVBHC_9_LC_16_18_6  (
            .in0(N__34370),
            .in1(N__23612),
            .in2(N__23666),
            .in3(N__23465),
            .lcout(\this_ppu.un1_M_surface_x_q_c1 ),
            .ltout(\this_ppu.un1_M_surface_x_q_c1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_RNIOOTPD_1_LC_16_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNIOOTPD_1_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNIOOTPD_1_LC_16_18_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNIOOTPD_1_LC_16_18_7  (
            .in0(N__23398),
            .in1(N__23343),
            .in2(N__23320),
            .in3(N__23310),
            .lcout(\this_ppu.un1_M_surface_x_q_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_11_LC_16_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_11_LC_16_19_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_11_LC_16_19_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_ppu.M_state_q_11_LC_16_19_0  (
            .in0(N__23203),
            .in1(N__24424),
            .in2(_gnd_net_),
            .in3(N__43243),
            .lcout(\this_ppu.M_state_qZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41997),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI41OT_10_LC_16_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI41OT_10_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI41OT_10_LC_16_19_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_RNI41OT_10_LC_16_19_2  (
            .in0(N__24142),
            .in1(N__23242),
            .in2(N__24223),
            .in3(N__23201),
            .lcout(\this_ppu.N_798_0 ),
            .ltout(\this_ppu.N_798_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIDPQ54_3_LC_16_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIDPQ54_3_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIDPQ54_3_LC_16_19_3 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIDPQ54_3_LC_16_19_3  (
            .in0(N__23166),
            .in1(N__23752),
            .in2(N__23128),
            .in3(N__34306),
            .lcout(M_this_ppu_vram_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_3_LC_16_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_3_LC_16_19_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_3_LC_16_19_6 .LUT_INIT=16'b1000010010001000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_3_LC_16_19_6  (
            .in0(N__25310),
            .in1(N__25528),
            .in2(N__25288),
            .in3(N__25483),
            .lcout(\this_ppu.M_pixel_cnt_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41997),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_595_LC_16_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_595_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_x_q_595_LC_16_20_2 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \this_ppu.M_screen_x_q_595_LC_16_20_2  (
            .in0(N__24311),
            .in1(N__23111),
            .in2(N__26141),
            .in3(N__25917),
            .lcout(\this_ppu.N_1659_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIPR8F3_5_LC_16_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIPR8F3_5_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIPR8F3_5_LC_16_20_3 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \this_ppu.M_state_q_RNIPR8F3_5_LC_16_20_3  (
            .in0(N__24341),
            .in1(N__23602),
            .in2(N__23082),
            .in3(N__24401),
            .lcout(\this_ppu.M_pixel_cnt_q_600_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_16_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_16_20_5 .LUT_INIT=16'b0011000100111011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_m2_LC_16_20_5  (
            .in0(N__26170),
            .in1(N__28483),
            .in2(N__25990),
            .in3(N__25975),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKTRBBJ2_6_LC_16_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKTRBBJ2_6_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKTRBBJ2_6_LC_16_20_6 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIKTRBBJ2_6_LC_16_20_6  (
            .in0(N__23866),
            .in1(N__28363),
            .in2(N__23857),
            .in3(N__27796),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_7_LC_16_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_7_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_7_LC_16_20_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_ppu.M_state_q_7_LC_16_20_7  (
            .in0(N__23835),
            .in1(N__26128),
            .in2(_gnd_net_),
            .in3(N__23797),
            .lcout(\this_ppu.M_state_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42004),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_0_LC_16_21_1 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_0_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_0_LC_16_21_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_0_LC_16_21_1  (
            .in0(N__23886),
            .in1(N__25508),
            .in2(_gnd_net_),
            .in3(N__25463),
            .lcout(\this_ppu.M_pixel_cnt_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42015),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNIF1DJ_7_LC_16_21_2 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_RNIF1DJ_7_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNIF1DJ_7_LC_16_21_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNIF1DJ_7_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(N__24693),
            .in2(_gnd_net_),
            .in3(N__23885),
            .lcout(\this_ppu.M_state_d30_i_i_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_0_LC_16_21_3 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_0_LC_16_21_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_0_LC_16_21_3 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \this_ppu.M_screen_x_q_0_LC_16_21_3  (
            .in0(N__23553),
            .in1(N__23498),
            .in2(N__26142),
            .in3(N__24664),
            .lcout(M_this_ppu_vram_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42015),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_1_LC_16_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_1_LC_16_21_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_1_LC_16_21_4 .LUT_INIT=16'b0100100011000000;
    LogicCell40 \this_ppu.M_screen_x_q_1_LC_16_21_4  (
            .in0(N__23499),
            .in1(N__23773),
            .in2(N__23535),
            .in3(N__23554),
            .lcout(M_this_ppu_vram_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42015),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIF77F7_3_LC_16_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIF77F7_3_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIF77F7_3_LC_16_21_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIF77F7_3_LC_16_21_5  (
            .in0(N__23749),
            .in1(N__39459),
            .in2(N__23698),
            .in3(N__37740),
            .lcout(\this_ppu.M_screen_y_q_esr_RNIF77F7Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIB9B9C_11_LC_16_21_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIB9B9C_11_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIB9B9C_11_LC_16_21_6 .LUT_INIT=16'b0000111011111110;
    LogicCell40 \this_ppu.M_state_q_RNIB9B9C_11_LC_16_21_6  (
            .in0(N__23667),
            .in1(N__24221),
            .in2(N__23613),
            .in3(N__34375),
            .lcout(\this_ppu.N_61_0 ),
            .ltout(\this_ppu.N_61_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_RNIM77RC_1_LC_16_21_7 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_RNIM77RC_1_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_x_q_RNIM77RC_1_LC_16_21_7 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \this_ppu.M_screen_x_q_RNIM77RC_1_LC_16_21_7  (
            .in0(_gnd_net_),
            .in1(N__23528),
            .in2(N__23515),
            .in3(N__23497),
            .lcout(\this_ppu.un1_M_screen_x_q_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNIS5KD2_3_LC_16_22_0 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_RNIS5KD2_3_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNIS5KD2_3_LC_16_22_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNIS5KD2_3_LC_16_22_0  (
            .in0(N__25311),
            .in1(N__24520),
            .in2(N__25441),
            .in3(N__24436),
            .lcout(\this_ppu.N_79_0 ),
            .ltout(\this_ppu.N_79_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_7_LC_16_22_1 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_7_LC_16_22_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_7_LC_16_22_1 .LUT_INIT=16'b0000000010101111;
    LogicCell40 \this_ppu.M_pixel_cnt_q_7_LC_16_22_1  (
            .in0(N__24343),
            .in1(_gnd_net_),
            .in2(N__24367),
            .in3(N__24526),
            .lcout(\this_ppu.M_pixel_cnt_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42023),
            .ce(),
            .sr(N__43109));
    defparam \this_ppu.M_state_q_RNIKF0ID_1_LC_16_22_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIKF0ID_1_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIKF0ID_1_LC_16_22_2 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \this_ppu.M_state_q_RNIKF0ID_1_LC_16_22_2  (
            .in0(N__24364),
            .in1(N__24229),
            .in2(N__24355),
            .in3(N__26137),
            .lcout(\this_ppu.N_1730_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIQ0NP8_0_LC_16_22_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIQ0NP8_0_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIQ0NP8_0_LC_16_22_5 .LUT_INIT=16'b1100010100000101;
    LogicCell40 \this_ppu.M_state_q_RNIQ0NP8_0_LC_16_22_5  (
            .in0(N__24342),
            .in1(N__24301),
            .in2(N__24271),
            .in3(N__25585),
            .lcout(\this_ppu.N_1042_0 ),
            .ltout(\this_ppu.N_1042_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIV84EA_11_LC_16_22_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIV84EA_11_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIV84EA_11_LC_16_22_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_ppu.M_state_q_RNIV84EA_11_LC_16_22_6  (
            .in0(N__24222),
            .in1(N__24180),
            .in2(N__23908),
            .in3(N__23905),
            .lcout(\this_ppu.N_677_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_c_LC_16_23_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_c_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_c_LC_16_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_c_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(N__23890),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_LUT4_0_LC_16_23_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_LUT4_0_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_LUT4_0_LC_16_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_LUT4_0_LC_16_23_1  (
            .in0(_gnd_net_),
            .in1(N__24504),
            .in2(N__25073),
            .in3(N__23872),
            .lcout(\this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_LUT4_0_LC_16_23_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_LUT4_0_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_LUT4_0_LC_16_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_LUT4_0_LC_16_23_2  (
            .in0(_gnd_net_),
            .in1(N__25009),
            .in2(N__24478),
            .in3(N__23869),
            .lcout(\this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_LUT4_0_LC_16_23_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_LUT4_0_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_LUT4_0_LC_16_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_LUT4_0_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(N__25312),
            .in2(N__25074),
            .in3(N__25273),
            .lcout(\this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_LUT4_0_LC_16_23_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_LUT4_0_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_LUT4_0_LC_16_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_LUT4_0_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(N__25013),
            .in2(N__25439),
            .in3(N__25270),
            .lcout(\this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_LUT4_0_LC_16_23_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_LUT4_0_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_LUT4_0_LC_16_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_LUT4_0_LC_16_23_5  (
            .in0(_gnd_net_),
            .in1(N__24451),
            .in2(N__25075),
            .in3(N__25267),
            .lcout(\this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_LUT4_0_LC_16_23_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_LUT4_0_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_LUT4_0_LC_16_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_LUT4_0_LC_16_23_6  (
            .in0(_gnd_net_),
            .in1(N__25017),
            .in2(N__25555),
            .in3(N__24697),
            .lcout(\this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_7_LC_16_23_7 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_7_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_7_LC_16_23_7 .LUT_INIT=16'b0000010100001001;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNO_0_7_LC_16_23_7  (
            .in0(N__24694),
            .in1(N__25462),
            .in2(N__24680),
            .in3(N__24529),
            .lcout(\this_ppu.N_1205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNIU2Q61_1_LC_16_24_0 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_RNIU2Q61_1_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNIU2Q61_1_LC_16_24_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNIU2Q61_1_LC_16_24_0  (
            .in0(N__24449),
            .in1(N__24473),
            .in2(N__25550),
            .in3(N__24500),
            .lcout(\this_ppu.M_state_d30_i_i_o2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_1_LC_16_24_1 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_1_LC_16_24_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_1_LC_16_24_1 .LUT_INIT=16'b1000001010100000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_1_LC_16_24_1  (
            .in0(N__25523),
            .in1(N__24511),
            .in2(N__24505),
            .in3(N__25478),
            .lcout(\this_ppu.M_pixel_cnt_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42039),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_2_LC_16_24_2 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_2_LC_16_24_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_2_LC_16_24_2 .LUT_INIT=16'b1100011000000000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_2_LC_16_24_2  (
            .in0(N__25479),
            .in1(N__24474),
            .in2(N__24487),
            .in3(N__25524),
            .lcout(\this_ppu.M_pixel_cnt_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42039),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_5_LC_16_24_3 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_5_LC_16_24_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_5_LC_16_24_3 .LUT_INIT=16'b1000001010001000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_5_LC_16_24_3  (
            .in0(N__25526),
            .in1(N__24450),
            .in2(N__24460),
            .in3(N__25481),
            .lcout(\this_ppu.M_pixel_cnt_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42039),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_16_LC_16_24_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_16_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_16_LC_16_24_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_16_LC_16_24_4  (
            .in0(N__26265),
            .in1(N__26283),
            .in2(_gnd_net_),
            .in3(N__26253),
            .lcout(\this_ppu.N_1301 ),
            .ltout(\this_ppu.N_1301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_data_count_qlde_i_0_i_LC_16_24_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_data_count_qlde_i_0_i_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_data_count_qlde_i_0_i_LC_16_24_5 .LUT_INIT=16'b0101010111111101;
    LogicCell40 \this_ppu.M_this_data_count_qlde_i_0_i_LC_16_24_5  (
            .in0(N__27562),
            .in1(N__35785),
            .in2(N__25564),
            .in3(N__37438),
            .lcout(N_231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_6_LC_16_24_6 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_6_LC_16_24_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_6_LC_16_24_6 .LUT_INIT=16'b1101001000000000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_6_LC_16_24_6  (
            .in0(N__25482),
            .in1(N__25561),
            .in2(N__25551),
            .in3(N__25527),
            .lcout(\this_ppu.M_pixel_cnt_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42039),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_4_LC_16_24_7 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_4_LC_16_24_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_4_LC_16_24_7 .LUT_INIT=16'b1000001010100000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_4_LC_16_24_7  (
            .in0(N__25525),
            .in1(N__25492),
            .in2(N__25440),
            .in3(N__25480),
            .lcout(\this_ppu.M_pixel_cnt_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42039),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_7_LC_16_25_0.C_ON=1'b0;
    defparam M_this_data_count_q_7_LC_16_25_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_16_25_0.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_7_LC_16_25_0 (
            .in0(N__25411),
            .in1(N__25737),
            .in2(_gnd_net_),
            .in3(N__27549),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42050),
            .ce(N__25365),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_9_LC_16_25_1.C_ON=1'b0;
    defparam M_this_data_count_q_9_LC_16_25_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_16_25_1.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_9_LC_16_25_1 (
            .in0(N__27550),
            .in1(N__25399),
            .in2(_gnd_net_),
            .in3(N__25388),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42050),
            .ce(N__25365),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_2_LC_16_25_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_2_LC_16_25_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_2_LC_16_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_2_LC_16_25_5  (
            .in0(N__26674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25339),
            .lcout(M_this_oam_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNIQFR31_2_LC_16_26_2.C_ON=1'b0;
    defparam M_this_oam_address_q_RNIQFR31_2_LC_16_26_2.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNIQFR31_2_LC_16_26_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_oam_address_q_RNIQFR31_2_LC_16_26_2 (
            .in0(N__26876),
            .in1(N__26838),
            .in2(N__26403),
            .in3(N__26791),
            .lcout(un1_M_this_oam_address_q_c3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_10_16_LC_16_26_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_10_16_LC_16_26_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_10_16_LC_16_26_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_10_16_LC_16_26_3  (
            .in0(N__25733),
            .in1(N__25716),
            .in2(_gnd_net_),
            .in3(N__25693),
            .lcout(\this_ppu.M_this_state_q_srsts_i_a2_10Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI13IA1_1_1_LC_16_26_4.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI13IA1_1_1_LC_16_26_4.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI13IA1_1_1_LC_16_26_4.LUT_INIT=16'b1111111100000100;
    LogicCell40 M_this_oam_address_q_RNI13IA1_1_1_LC_16_26_4 (
            .in0(N__26839),
            .in1(N__26792),
            .in2(N__26888),
            .in3(N__43226),
            .lcout(N_1709_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI13IA1_1_LC_16_26_7.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI13IA1_1_LC_16_26_7.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI13IA1_1_LC_16_26_7.LUT_INIT=16'b1010101011101010;
    LogicCell40 M_this_oam_address_q_RNI13IA1_1_LC_16_26_7 (
            .in0(N__43227),
            .in1(N__26880),
            .in2(N__26797),
            .in3(N__26840),
            .lcout(N_1693_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI01JU6_9_LC_17_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI01JU6_9_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI01JU6_9_LC_17_16_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI01JU6_9_LC_17_16_2  (
            .in0(N__27298),
            .in1(N__27074),
            .in2(N__25969),
            .in3(N__30466),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNI01JU6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un30_0_a2_i_a2_1_LC_17_17_0 .C_ON=1'b0;
    defparam \this_ppu.un30_0_a2_i_a2_1_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un30_0_a2_i_a2_1_LC_17_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.un30_0_a2_i_a2_1_LC_17_17_0  (
            .in0(N__35142),
            .in1(N__35004),
            .in2(N__26235),
            .in3(N__30687),
            .lcout(),
            .ltout(\this_ppu.N_1269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un30_0_a2_i_o2_LC_17_17_1 .C_ON=1'b0;
    defparam \this_ppu.un30_0_a2_i_o2_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un30_0_a2_i_o2_LC_17_17_1 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \this_ppu.un30_0_a2_i_o2_LC_17_17_1  (
            .in0(N__26357),
            .in1(N__26199),
            .in2(N__25588),
            .in3(N__30588),
            .lcout(\this_ppu.N_1006_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_8_LC_17_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_8_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_8_LC_17_17_2 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_8_LC_17_17_2  (
            .in0(N__35141),
            .in1(N__30686),
            .in2(N__30451),
            .in3(N__30173),
            .lcout(N_782_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_6_LC_17_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_6_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_6_LC_17_17_4 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_6_LC_17_17_4  (
            .in0(N__29760),
            .in1(_gnd_net_),
            .in2(N__29718),
            .in3(N__28261),
            .lcout(\this_vga_signals.N_1264 ),
            .ltout(\this_vga_signals.N_1264_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_ns_LC_17_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_ns_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_ns_LC_17_17_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_ns_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__25846),
            .in2(N__25573),
            .in3(N__25570),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_4_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_x0_LC_17_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_x0_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_x0_LC_17_17_6 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_x0_LC_17_17_6  (
            .in0(N__29706),
            .in1(N__29838),
            .in2(N__29766),
            .in3(N__29619),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_x1_LC_17_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_x1_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_x1_LC_17_17_7 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_x1_LC_17_17_7  (
            .in0(N__29618),
            .in1(N__29756),
            .in2(N__29849),
            .in3(N__29707),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_scroll_q_esr_10_LC_17_18_0.C_ON=1'b0;
    defparam M_this_scroll_q_esr_10_LC_17_18_0.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_10_LC_17_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_10_LC_17_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42772),
            .lcout(M_this_scroll_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42002),
            .ce(N__26326),
            .sr(N__43104));
    defparam M_this_scroll_q_esr_11_LC_17_18_1.C_ON=1'b0;
    defparam M_this_scroll_q_esr_11_LC_17_18_1.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_11_LC_17_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_11_LC_17_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41474),
            .lcout(M_this_scroll_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42002),
            .ce(N__26326),
            .sr(N__43104));
    defparam M_this_scroll_q_esr_12_LC_17_18_2.C_ON=1'b0;
    defparam M_this_scroll_q_esr_12_LC_17_18_2.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_12_LC_17_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_12_LC_17_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40786),
            .lcout(M_this_scroll_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42002),
            .ce(N__26326),
            .sr(N__43104));
    defparam M_this_scroll_q_esr_13_LC_17_18_3.C_ON=1'b0;
    defparam M_this_scroll_q_esr_13_LC_17_18_3.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_13_LC_17_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_13_LC_17_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40039),
            .lcout(M_this_scroll_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42002),
            .ce(N__26326),
            .sr(N__43104));
    defparam M_this_scroll_q_esr_14_LC_17_18_4.C_ON=1'b0;
    defparam M_this_scroll_q_esr_14_LC_17_18_4.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_14_LC_17_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_14_LC_17_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40420),
            .lcout(M_this_scroll_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42002),
            .ce(N__26326),
            .sr(N__43104));
    defparam M_this_scroll_q_esr_15_LC_17_18_5.C_ON=1'b0;
    defparam M_this_scroll_q_esr_15_LC_17_18_5.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_15_LC_17_18_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_15_LC_17_18_5 (
            .in0(N__39906),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42002),
            .ce(N__26326),
            .sr(N__43104));
    defparam M_this_scroll_q_esr_8_LC_17_18_6.C_ON=1'b0;
    defparam M_this_scroll_q_esr_8_LC_17_18_6.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_8_LC_17_18_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_8_LC_17_18_6 (
            .in0(N__42449),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42002),
            .ce(N__26326),
            .sr(N__43104));
    defparam M_this_scroll_q_esr_9_LC_17_18_7.C_ON=1'b0;
    defparam M_this_scroll_q_esr_9_LC_17_18_7.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_9_LC_17_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_9_LC_17_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39782),
            .lcout(M_this_scroll_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42002),
            .ce(N__26326),
            .sr(N__43104));
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_17_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_17_19_0 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_14_LC_17_19_0  (
            .in0(N__29320),
            .in1(N__28524),
            .in2(N__27163),
            .in3(N__27151),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_17_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_17_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_LC_17_19_1  (
            .in0(N__25981),
            .in1(N__28664),
            .in2(N__25993),
            .in3(N__27817),
            .lcout(\this_vga_signals.N_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_LC_17_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_LC_17_19_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_x2_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(N__28930),
            .in2(_gnd_net_),
            .in3(N__27433),
            .lcout(\this_vga_signals.g0_0_x2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m1_0_x2_1_LC_17_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m1_0_x2_1_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m1_0_x2_1_LC_17_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m1_0_x2_1_LC_17_19_5  (
            .in0(N__28931),
            .in1(N__27828),
            .in2(_gnd_net_),
            .in3(N__27004),
            .lcout(\this_vga_signals.if_m1_0_x2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_4_LC_17_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_4_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_4_LC_17_19_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_4_LC_17_19_7  (
            .in0(N__34973),
            .in1(N__35321),
            .in2(N__26228),
            .in3(N__30581),
            .lcout(\this_vga_signals.N_836_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_33_LC_17_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_33_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_33_LC_17_20_0 .LUT_INIT=16'b1001110000111001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_33_LC_17_20_0  (
            .in0(N__28904),
            .in1(N__28957),
            .in2(N__35491),
            .in3(N__27124),
            .lcout(\this_vga_signals.r_N_2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_17_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_17_20_1 .LUT_INIT=16'b0101100001011010;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_1_LC_17_20_1  (
            .in0(N__27116),
            .in1(N__25961),
            .in2(N__25885),
            .in3(N__30453),
            .lcout(),
            .ltout(\this_vga_signals.N_1043_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_1_LC_17_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_1_LC_17_20_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_1_LC_17_20_2 .LUT_INIT=16'b1110010011000100;
    LogicCell40 \this_vga_signals.M_lcounter_q_1_LC_17_20_2  (
            .in0(N__27333),
            .in1(N__25879),
            .in2(N__25942),
            .in3(N__25939),
            .lcout(this_vga_signals_M_lcounter_q_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42019),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_LC_17_20_3 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_LC_17_20_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.line_clk.M_last_q_LC_17_20_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.line_clk.M_last_q_LC_17_20_3  (
            .in0(N__25938),
            .in1(N__25918),
            .in2(N__25886),
            .in3(N__30454),
            .lcout(\this_ppu.M_last_q_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42019),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_17_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_17_20_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_17_20_4  (
            .in0(N__28903),
            .in1(N__27425),
            .in2(N__35490),
            .in3(N__27026),
            .lcout(N_771_0),
            .ltout(N_771_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_3_LC_17_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_3_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_3_LC_17_20_5 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_o2_3_LC_17_20_5  (
            .in0(N__35301),
            .in1(_gnd_net_),
            .in2(N__26203),
            .in3(N__34993),
            .lcout(\this_ppu.N_774_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_17_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_17_20_6 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_17_20_6  (
            .in0(N__34994),
            .in1(N__35302),
            .in2(_gnd_net_),
            .in3(N__34750),
            .lcout(\this_vga_signals.g1_0_0 ),
            .ltout(\this_vga_signals.g1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_17_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_17_20_7 .LUT_INIT=16'b0111000100010111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_36_LC_17_20_7  (
            .in0(N__34995),
            .in1(N__27956),
            .in2(N__26173),
            .in3(N__35153),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_17_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_17_21_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_22_LC_17_21_1  (
            .in0(N__27431),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27027),
            .lcout(\this_vga_signals.if_N_6_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIP1DV3_7_LC_17_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIP1DV3_7_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIP1DV3_7_LC_17_21_4 .LUT_INIT=16'b1101001000101101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIP1DV3_7_LC_17_21_4  (
            .in0(N__27991),
            .in1(N__30328),
            .in2(N__26164),
            .in3(N__35150),
            .lcout(),
            .ltout(\this_vga_signals.N_27_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_17_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_17_21_5 .LUT_INIT=16'b1100000001001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_35_LC_17_21_5  (
            .in0(N__35000),
            .in1(N__28423),
            .in2(N__26155),
            .in3(N__26152),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_33_N_4L6_LC_17_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_33_N_4L6_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_33_N_4L6_LC_17_21_6 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_33_N_4L6_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26146),
            .in3(N__28525),
            .lcout(\this_vga_signals.g0_33_N_4L6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_12_LC_17_21_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_12_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_12_LC_17_21_7 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_1_12_LC_17_21_7  (
            .in0(N__35783),
            .in1(N__36534),
            .in2(N__26143),
            .in3(N__27145),
            .lcout(\this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNI9A3Q6_6_LC_17_22_0 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNI9A3Q6_6_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNI9A3Q6_6_LC_17_22_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNI9A3Q6_6_LC_17_22_0  (
            .in0(N__26367),
            .in1(N__37696),
            .in2(N__36571),
            .in3(N__28039),
            .lcout(\this_ppu.N_753_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIO37G1_7_LC_17_22_2.C_ON=1'b0;
    defparam M_this_state_q_RNIO37G1_7_LC_17_22_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIO37G1_7_LC_17_22_2.LUT_INIT=16'b1111010011110000;
    LogicCell40 M_this_state_q_RNIO37G1_7_LC_17_22_2 (
            .in0(N__29053),
            .in1(N__30936),
            .in2(N__43251),
            .in3(N__43415),
            .lcout(N_1725_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIKQ691_7_LC_17_22_7.C_ON=1'b0;
    defparam M_this_state_q_RNIKQ691_7_LC_17_22_7.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIKQ691_7_LC_17_22_7.LUT_INIT=16'b1110111011001100;
    LogicCell40 M_this_state_q_RNIKQ691_7_LC_17_22_7 (
            .in0(N__43416),
            .in1(N__43232),
            .in2(_gnd_net_),
            .in3(N__29052),
            .lcout(N_1717_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_0_13_LC_17_23_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_0_13_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_0_13_LC_17_23_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_o2_0_13_LC_17_23_1  (
            .in0(_gnd_net_),
            .in1(N__35763),
            .in2(_gnd_net_),
            .in3(N__29190),
            .lcout(\this_ppu.N_1002_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_12_LC_17_23_2.C_ON=1'b0;
    defparam M_this_state_q_12_LC_17_23_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_12_LC_17_23_2.LUT_INIT=16'b1100110011001000;
    LogicCell40 M_this_state_q_12_LC_17_23_2 (
            .in0(N__36535),
            .in1(N__26314),
            .in2(N__33171),
            .in3(N__27384),
            .lcout(M_this_state_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42044),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_17_23_3 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_17_23_3 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_17_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_17_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26305),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42044),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNIR3631_1_LC_17_24_0.C_ON=1'b0;
    defparam M_this_oam_address_q_RNIR3631_1_LC_17_24_0.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNIR3631_1_LC_17_24_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_oam_address_q_RNIR3631_1_LC_17_24_0 (
            .in0(N__28168),
            .in1(N__26843),
            .in2(N__26890),
            .in3(N__43371),
            .lcout(un1_M_this_oam_address_q_c2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_0_o2_0_LC_17_24_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_0_o2_0_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_0_o2_0_LC_17_24_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_0_o2_0_LC_17_24_1  (
            .in0(N__26290),
            .in1(N__37427),
            .in2(N__26272),
            .in3(N__26254),
            .lcout(\this_ppu.N_767_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_17_24_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_17_24_3 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_17_24_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_17_24_3  (
            .in0(N__27588),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27675),
            .lcout(this_start_data_delay_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42056),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_data_tmp_d_1_sqmuxa_i_0_o3_LC_17_24_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_data_tmp_d_1_sqmuxa_i_0_o3_LC_17_24_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_data_tmp_d_1_sqmuxa_i_0_o3_LC_17_24_5 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \this_ppu.M_this_data_tmp_d_1_sqmuxa_i_0_o3_LC_17_24_5  (
            .in0(N__27587),
            .in1(N__27615),
            .in2(N__27681),
            .in3(N__28167),
            .lcout(N_778_0),
            .ltout(N_778_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI13IA1_0_1_LC_17_24_6.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI13IA1_0_1_LC_17_24_6.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI13IA1_0_1_LC_17_24_6.LUT_INIT=16'b1111111101000000;
    LogicCell40 M_this_oam_address_q_RNI13IA1_0_1_LC_17_24_6 (
            .in0(N__26887),
            .in1(N__26844),
            .in2(N__26566),
            .in3(N__43228),
            .lcout(N_1701_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_0_LC_17_25_3.C_ON=1'b0;
    defparam M_this_oam_address_q_0_LC_17_25_3.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_0_LC_17_25_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_oam_address_q_0_LC_17_25_3 (
            .in0(N__27464),
            .in1(N__26841),
            .in2(_gnd_net_),
            .in3(N__26789),
            .lcout(M_this_oam_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42067),
            .ce(),
            .sr(N__41641));
    defparam M_this_oam_address_q_5_LC_17_25_4.C_ON=1'b0;
    defparam M_this_oam_address_q_5_LC_17_25_4.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_5_LC_17_25_4.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_5_LC_17_25_4 (
            .in0(N__26497),
            .in1(N__27463),
            .in2(_gnd_net_),
            .in3(N__26527),
            .lcout(M_this_oam_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42067),
            .ce(),
            .sr(N__41641));
    defparam M_this_oam_address_q_RNIRA651_4_LC_17_25_5.C_ON=1'b0;
    defparam M_this_oam_address_q_RNIRA651_4_LC_17_25_5.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNIRA651_4_LC_17_25_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_oam_address_q_RNIRA651_4_LC_17_25_5 (
            .in0(N__26970),
            .in1(N__26426),
            .in2(N__26924),
            .in3(N__26397),
            .lcout(un1_M_this_oam_address_q_c5),
            .ltout(un1_M_this_oam_address_q_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_6_LC_17_25_6.C_ON=1'b0;
    defparam M_this_oam_address_q_6_LC_17_25_6.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_6_LC_17_25_6.LUT_INIT=16'b0000000001101100;
    LogicCell40 M_this_oam_address_q_6_LC_17_25_6 (
            .in0(N__26498),
            .in1(N__26447),
            .in2(N__26473),
            .in3(N__27466),
            .lcout(M_this_oam_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42067),
            .ce(),
            .sr(N__41641));
    defparam M_this_oam_address_q_3_LC_17_25_7.C_ON=1'b0;
    defparam M_this_oam_address_q_3_LC_17_25_7.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_3_LC_17_25_7.LUT_INIT=16'b0001010001010000;
    LogicCell40 M_this_oam_address_q_3_LC_17_25_7 (
            .in0(N__27465),
            .in1(N__26427),
            .in2(N__26981),
            .in3(N__26398),
            .lcout(M_this_oam_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42067),
            .ce(),
            .sr(N__41641));
    defparam M_this_oam_address_q_1_LC_17_26_0.C_ON=1'b0;
    defparam M_this_oam_address_q_1_LC_17_26_0.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_1_LC_17_26_0.LUT_INIT=16'b0001001000110000;
    LogicCell40 M_this_oam_address_q_1_LC_17_26_0 (
            .in0(N__26842),
            .in1(N__27482),
            .in2(N__26889),
            .in3(N__26796),
            .lcout(M_this_oam_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42078),
            .ce(),
            .sr(N__41639));
    defparam M_this_oam_address_q_2_LC_17_26_4.C_ON=1'b0;
    defparam M_this_oam_address_q_2_LC_17_26_4.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_2_LC_17_26_4.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_2_LC_17_26_4 (
            .in0(N__26399),
            .in1(N__27480),
            .in2(_gnd_net_),
            .in3(N__26431),
            .lcout(M_this_oam_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42078),
            .ce(),
            .sr(N__41639));
    defparam M_this_oam_address_q_4_LC_17_26_5.C_ON=1'b0;
    defparam M_this_oam_address_q_4_LC_17_26_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_4_LC_17_26_5.LUT_INIT=16'b0001010001010000;
    LogicCell40 M_this_oam_address_q_4_LC_17_26_5 (
            .in0(N__27481),
            .in1(N__26977),
            .in2(N__26925),
            .in3(N__26944),
            .lcout(M_this_oam_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42078),
            .ce(),
            .sr(N__41639));
    defparam \this_ppu.M_this_oam_ram_write_data_0_sqmuxa_0_a3_0_a2_LC_17_27_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_sqmuxa_0_a3_0_a2_LC_17_27_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_sqmuxa_0_a3_0_a2_LC_17_27_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_sqmuxa_0_a3_0_a2_LC_17_27_4  (
            .in0(N__26875),
            .in1(N__26845),
            .in2(_gnd_net_),
            .in3(N__26790),
            .lcout(M_this_oam_ram_write_data_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_18_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_18_17_0 .LUT_INIT=16'b0110011011011101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_18_17_0  (
            .in0(N__29929),
            .in1(N__29876),
            .in2(_gnd_net_),
            .in3(N__29842),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_c_0_1 ),
            .ltout(\this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_LC_18_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_LC_18_17_1 .LUT_INIT=16'b0011001000110001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_LC_18_17_1  (
            .in0(N__30535),
            .in1(N__27763),
            .in2(N__26572),
            .in3(N__29626),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_0_1 ),
            .ltout(\this_vga_signals.mult1_un47_sum_ac0_3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_18_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_18_17_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_18_17_2  (
            .in0(N__28702),
            .in1(_gnd_net_),
            .in2(N__26569),
            .in3(N__34990),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_18_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_18_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_18_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28293),
            .lcout(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42003),
            .ce(N__34246),
            .sr(N__34214));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_18_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_18_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_18_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30762),
            .lcout(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42003),
            .ce(N__34246),
            .sr(N__34214));
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_18_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_18_17_5 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_LC_18_17_5  (
            .in0(N__34991),
            .in1(N__28703),
            .in2(N__27187),
            .in3(N__28748),
            .lcout(\this_vga_signals.g0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_18_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_18_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_18_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30725),
            .lcout(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42003),
            .ce(N__34246),
            .sr(N__34214));
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_18_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_18_17_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_LC_18_17_7  (
            .in0(N__34992),
            .in1(N__28704),
            .in2(_gnd_net_),
            .in3(N__28749),
            .lcout(\this_vga_signals.mult1_un54_sum_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_18_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_18_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_18_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27708),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42009),
            .ce(N__34248),
            .sr(N__34215));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_18_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_18_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_18_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34277),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42009),
            .ce(N__34248),
            .sr(N__34215));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_18_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_18_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_18_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28292),
            .lcout(this_vga_signals_M_vcounter_q_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42009),
            .ce(N__34248),
            .sr(N__34215));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_18_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_18_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_18_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28325),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42009),
            .ce(N__34248),
            .sr(N__34215));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_18_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_18_19_1 .LUT_INIT=16'b0001001001111011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_18_19_1  (
            .in0(N__35408),
            .in1(N__35515),
            .in2(N__28986),
            .in3(N__35248),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_18_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_18_19_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_18_19_2  (
            .in0(N__28584),
            .in1(N__28977),
            .in2(_gnd_net_),
            .in3(N__35409),
            .lcout(\this_vga_signals.mult1_un61_sum_axb2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_0_LC_18_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_0_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_0_LC_18_19_3 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_0_LC_18_19_3  (
            .in0(N__29764),
            .in1(N__29714),
            .in2(_gnd_net_),
            .in3(N__29620),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI0FP_LC_18_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI0FP_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI0FP_LC_18_19_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI0FP_LC_18_19_4  (
            .in0(N__29715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28196),
            .lcout(\this_vga_signals.vaddress_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_LC_18_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_LC_18_19_6 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_LC_18_19_6  (
            .in0(N__27949),
            .in1(N__34881),
            .in2(_gnd_net_),
            .in3(N__27910),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_33_N_3L4_LC_18_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_33_N_3L4_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_33_N_3L4_LC_18_19_7 .LUT_INIT=16'b1010010100001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_33_N_3L4_LC_18_19_7  (
            .in0(N__28705),
            .in1(_gnd_net_),
            .in2(N__34943),
            .in3(N__28768),
            .lcout(\this_vga_signals.g0_33_N_3L4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_18_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_18_20_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_24_LC_18_20_0  (
            .in0(N__34967),
            .in1(N__28711),
            .in2(_gnd_net_),
            .in3(N__28766),
            .lcout(\this_vga_signals.mult1_un54_sum_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_18_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_18_20_1 .LUT_INIT=16'b1000100000101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_19_LC_18_20_1  (
            .in0(N__28424),
            .in1(N__27838),
            .in2(N__34999),
            .in3(N__28383),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_18_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_18_20_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_17_LC_18_20_2  (
            .in0(N__34966),
            .in1(N__28712),
            .in2(_gnd_net_),
            .in3(N__28767),
            .lcout(\this_vga_signals.mult1_un54_sum_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_18_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_18_20_3 .LUT_INIT=16'b0011100111000110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_LC_18_20_3  (
            .in0(N__29536),
            .in1(N__30112),
            .in2(N__29497),
            .in3(N__29572),
            .lcout(\this_vga_signals.mult1_un47_sum_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a3_1_12_LC_18_20_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a3_1_12_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a3_1_12_LC_18_20_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_a3_1_12_LC_18_20_4  (
            .in0(N__29201),
            .in1(N__36533),
            .in2(_gnd_net_),
            .in3(N__29289),
            .lcout(\this_ppu.N_1115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_33_N_5L8_LC_18_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_33_N_5L8_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_33_N_5L8_LC_18_20_5 .LUT_INIT=16'b0011011011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_33_N_5L8_LC_18_20_5  (
            .in0(N__29803),
            .in1(N__28666),
            .in2(N__27139),
            .in3(N__27130),
            .lcout(\this_vga_signals.g0_33_N_5L8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_18_21_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_18_21_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_18_21_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_18_21_0  (
            .in0(N__27326),
            .in1(N__27028),
            .in2(N__27118),
            .in3(N__27117),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_21_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__42037),
            .ce(),
            .sr(N__34219));
    defparam \this_vga_signals.M_vcounter_q_1_LC_18_21_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_18_21_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_18_21_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_18_21_1  (
            .in0(N__27328),
            .in1(N__27432),
            .in2(_gnd_net_),
            .in3(N__27010),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__42037),
            .ce(),
            .sr(N__34219));
    defparam \this_vga_signals.M_vcounter_q_2_LC_18_21_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_18_21_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_18_21_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_18_21_2  (
            .in0(N__27327),
            .in1(N__28928),
            .in2(_gnd_net_),
            .in3(N__27007),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__42037),
            .ce(),
            .sr(N__34219));
    defparam \this_vga_signals.M_vcounter_q_3_LC_18_21_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_18_21_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_18_21_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_18_21_3  (
            .in0(N__27329),
            .in1(N__35464),
            .in2(_gnd_net_),
            .in3(N__27208),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__42037),
            .ce(),
            .sr(N__34219));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_18_21_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_18_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_18_21_4  (
            .in0(_gnd_net_),
            .in1(N__35318),
            .in2(_gnd_net_),
            .in3(N__27205),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_18_21_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_18_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_18_21_5  (
            .in0(_gnd_net_),
            .in1(N__34947),
            .in2(_gnd_net_),
            .in3(N__27202),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_18_21_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_18_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_18_21_6  (
            .in0(_gnd_net_),
            .in1(N__34758),
            .in2(_gnd_net_),
            .in3(N__27199),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_18_21_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_18_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_18_21_7  (
            .in0(_gnd_net_),
            .in1(N__35151),
            .in2(_gnd_net_),
            .in3(N__27196),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_18_22_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_18_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_18_22_0  (
            .in0(_gnd_net_),
            .in1(N__30692),
            .in2(_gnd_net_),
            .in3(N__27193),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_18_22_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_18_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_18_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_18_22_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(N__30452),
            .in2(_gnd_net_),
            .in3(N__27190),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_18_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_18_22_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(N__27426),
            .in2(_gnd_net_),
            .in3(N__28905),
            .lcout(\this_vga_signals.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_o2_2_1_LC_18_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_o2_2_1_LC_18_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_o2_2_1_LC_18_22_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.IO_port_data_write_0_a2_i_o2_2_1_LC_18_22_3  (
            .in0(N__27874),
            .in1(N__30895),
            .in2(N__29155),
            .in3(N__36430),
            .lcout(\this_vga_signals.IO_port_data_write_0_a2_i_o2_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_18_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_18_22_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_18_22_5  (
            .in0(N__27427),
            .in1(N__35465),
            .in2(N__28929),
            .in3(N__35319),
            .lcout(\this_vga_signals.vsync_1_0_a3_0_a3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_13_LC_18_22_7.C_ON=1'b0;
    defparam M_this_state_q_13_LC_18_22_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_13_LC_18_22_7.LUT_INIT=16'b1111100000000000;
    LogicCell40 M_this_state_q_13_LC_18_22_7 (
            .in0(N__29082),
            .in1(N__27385),
            .in2(N__36442),
            .in3(N__31059),
            .lcout(M_this_state_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42045),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_data_count_qlde_i_0_o2_LC_18_23_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_data_count_qlde_i_0_o2_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_data_count_qlde_i_0_o2_LC_18_23_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.M_this_data_count_qlde_i_0_o2_LC_18_23_0  (
            .in0(N__27871),
            .in1(N__29144),
            .in2(_gnd_net_),
            .in3(N__27382),
            .lcout(N_816_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_1_18_LC_18_23_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_1_18_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_1_18_LC_18_23_1 .LUT_INIT=16'b0010001000100011;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_1_18_LC_18_23_1  (
            .in0(N__27616),
            .in1(N__43221),
            .in2(N__27682),
            .in3(N__27592),
            .lcout(\this_ppu.N_430_1_0 ),
            .ltout(\this_ppu.N_430_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_fast_13_LC_18_23_2.C_ON=1'b0;
    defparam M_this_state_q_fast_13_LC_18_23_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_fast_13_LC_18_23_2.LUT_INIT=16'b1111000010000000;
    LogicCell40 M_this_state_q_fast_13_LC_18_23_2 (
            .in0(N__29081),
            .in1(N__27383),
            .in2(N__27364),
            .in3(N__27361),
            .lcout(M_this_state_q_fastZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42057),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_18_LC_18_23_3.C_ON=1'b0;
    defparam M_this_state_q_18_LC_18_23_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_18_LC_18_23_3.LUT_INIT=16'b1110000010100000;
    LogicCell40 M_this_state_q_18_LC_18_23_3 (
            .in0(N__28163),
            .in1(N__29080),
            .in2(N__31075),
            .in3(N__27872),
            .lcout(M_this_state_qZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42057),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_38_i_0_a2_3_0_LC_18_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.N_38_i_0_a2_3_0_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_38_i_0_a2_3_0_LC_18_23_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.N_38_i_0_a2_3_0_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(N__27360),
            .in2(_gnd_net_),
            .in3(N__28162),
            .lcout(),
            .ltout(\this_vga_signals.N_38_i_0_a2_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_38_i_0_a2_3_x1_LC_18_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.N_38_i_0_a2_3_x1_LC_18_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_38_i_0_a2_3_x1_LC_18_23_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vga_signals.N_38_i_0_a2_3_x1_LC_18_23_5  (
            .in0(N__38588),
            .in1(N__29041),
            .in2(N__27352),
            .in3(N__37394),
            .lcout(),
            .ltout(\this_vga_signals.N_38_i_0_a2_3_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_38_i_0_a2_3_ns_LC_18_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.N_38_i_0_a2_3_ns_LC_18_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_38_i_0_a2_3_ns_LC_18_23_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vga_signals.N_38_i_0_a2_3_ns_LC_18_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27349),
            .in3(N__30805),
            .lcout(),
            .ltout(\this_vga_signals.N_38_i_0_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_38_i_0_o3_LC_18_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.N_38_i_0_o3_LC_18_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_38_i_0_o3_LC_18_23_7 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \this_vga_signals.N_38_i_0_o3_LC_18_23_7  (
            .in0(N__37426),
            .in1(N__27688),
            .in2(N__27691),
            .in3(N__36518),
            .lcout(N_38_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_38_i_0_a2_0_4_LC_18_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.N_38_i_0_a2_0_4_LC_18_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_38_i_0_a2_0_4_LC_18_24_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vga_signals.N_38_i_0_a2_0_4_LC_18_24_0  (
            .in0(N__30918),
            .in1(N__27883),
            .in2(N__36443),
            .in3(N__41060),
            .lcout(\this_vga_signals.N_38_i_0_a2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_0_15_LC_18_24_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_0_15_LC_18_24_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_0_15_LC_18_24_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_o2_0_15_LC_18_24_3  (
            .in0(N__27586),
            .in1(N__27679),
            .in2(_gnd_net_),
            .in3(N__27614),
            .lcout(\this_ppu.N_787_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_15_LC_18_24_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_15_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_15_LC_18_24_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_o2_15_LC_18_24_4  (
            .in0(N__27680),
            .in1(N__27613),
            .in2(_gnd_net_),
            .in3(N__27585),
            .lcout(N_765_0),
            .ltout(N_765_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_this_data_count_q4_i_0_366_i_0_1_LC_18_24_5 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_data_count_q4_i_0_366_i_0_1_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_data_count_q4_i_0_366_i_0_1_LC_18_24_5 .LUT_INIT=16'b0000000010101111;
    LogicCell40 \this_ppu.un1_M_this_data_count_q4_i_0_366_i_0_1_LC_18_24_5  (
            .in0(N__41061),
            .in1(_gnd_net_),
            .in2(N__27565),
            .in3(N__43219),
            .lcout(\this_ppu.N_229_1_0 ),
            .ltout(\this_ppu.N_229_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_this_data_count_q4_i_0_366_i_0_i_LC_18_24_6 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_data_count_q4_i_0_366_i_0_i_LC_18_24_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_data_count_q4_i_0_366_i_0_i_LC_18_24_6 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \this_ppu.un1_M_this_data_count_q4_i_0_366_i_0_i_LC_18_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27553),
            .in3(N__29194),
            .lcout(N_229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_data_count_d_5_sqmuxa_0_a3_i_o3_i_a2_LC_18_25_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_data_count_d_5_sqmuxa_0_a3_i_o3_i_a2_LC_18_25_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_data_count_d_5_sqmuxa_0_a3_i_o3_i_a2_LC_18_25_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_data_count_d_5_sqmuxa_0_a3_i_o3_i_a2_LC_18_25_2  (
            .in0(_gnd_net_),
            .in1(N__43372),
            .in2(_gnd_net_),
            .in3(N__29240),
            .lcout(N_1423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI99C6_5_LC_19_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI99C6_5_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI99C6_5_LC_19_17_1 .LUT_INIT=16'b0000011100000111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNI99C6_5_LC_19_17_1  (
            .in0(N__29705),
            .in1(N__29755),
            .in2(N__29644),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.SUM_2_i_i_1_0_3 ),
            .ltout(\this_vga_signals.SUM_2_i_i_1_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3GK81_8_LC_19_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3GK81_8_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3GK81_8_LC_19_17_2 .LUT_INIT=16'b1011110100100011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI3GK81_8_LC_19_17_2  (
            .in0(N__35137),
            .in1(N__30420),
            .in2(N__27436),
            .in3(N__30685),
            .lcout(\this_vga_signals.N_39_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_x1_LC_19_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_x1_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_x1_LC_19_17_3 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_x1_LC_19_17_3  (
            .in0(N__29703),
            .in1(N__29753),
            .in2(N__29643),
            .in3(N__27733),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_1_LC_19_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_1_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_1_LC_19_17_4 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_1_LC_19_17_4  (
            .in0(_gnd_net_),
            .in1(N__28229),
            .in2(N__28216),
            .in3(N__28253),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1 ),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_x0_LC_19_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_x0_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_x0_LC_19_17_5 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_x0_LC_19_17_5  (
            .in0(N__29704),
            .in1(_gnd_net_),
            .in2(N__27727),
            .in3(N__29754),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_1_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_ns_LC_19_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_ns_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_ns_LC_19_17_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_ns_LC_19_17_6  (
            .in0(_gnd_net_),
            .in1(N__29658),
            .in2(N__27724),
            .in3(N__27721),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_19_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_19_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_19_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_19_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28332),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42010),
            .ce(N__34247),
            .sr(N__34216));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_19_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_19_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_19_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_19_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27715),
            .lcout(this_vga_signals_M_vcounter_q_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42020),
            .ce(N__34250),
            .sr(N__34217));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIFI5N_LC_19_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIFI5N_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIFI5N_LC_19_18_2 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIFI5N_LC_19_18_2  (
            .in0(N__28195),
            .in1(N__35219),
            .in2(_gnd_net_),
            .in3(N__34705),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_18_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34284),
            .lcout(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42020),
            .ce(N__34250),
            .sr(N__34217));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_1_LC_19_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_1_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_1_LC_19_18_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_1_LC_19_18_4  (
            .in0(N__28194),
            .in1(N__29716),
            .in2(_gnd_net_),
            .in3(N__28237),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_0_ns_1_LC_19_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_0_ns_1_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_0_ns_1_LC_19_18_5 .LUT_INIT=16'b0100001000101000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_0_ns_1_LC_19_18_5  (
            .in0(N__29872),
            .in1(N__29831),
            .in2(N__29930),
            .in3(N__29621),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_ac0_3_0_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_0_ns_LC_19_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_0_ns_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_0_ns_LC_19_18_6 .LUT_INIT=16'b0110111110101111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_0_ns_LC_19_18_6  (
            .in0(N__29622),
            .in1(N__29765),
            .in2(N__27781),
            .in3(N__29717),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_0_0 ),
            .ltout(\this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_19_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_19_18_7 .LUT_INIT=16'b0000000010110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_19_18_7  (
            .in0(N__27778),
            .in1(N__27772),
            .in2(N__27766),
            .in3(N__27762),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m5_s_LC_19_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m5_s_LC_19_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m5_s_LC_19_19_0 .LUT_INIT=16'b0000011001100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m5_s_LC_19_19_0  (
            .in0(N__28937),
            .in1(N__35518),
            .in2(N__29008),
            .in3(N__28981),
            .lcout(),
            .ltout(\this_vga_signals.if_m5_s_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m5_LC_19_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m5_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m5_LC_19_19_1 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m5_LC_19_19_1  (
            .in0(N__28856),
            .in1(N__28650),
            .in2(N__27751),
            .in3(N__27742),
            .lcout(\this_vga_signals.mult1_un68_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_19_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_19_19_2 .LUT_INIT=16'b1111100110010000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_21_LC_19_19_2  (
            .in0(N__34735),
            .in1(N__34162),
            .in2(N__29988),
            .in3(N__34141),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_19_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_19_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_19_19_3 .LUT_INIT=16'b0000011001100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_0_LC_19_19_3  (
            .in0(N__35516),
            .in1(N__28935),
            .in2(N__27748),
            .in3(N__29002),
            .lcout(\this_vga_signals.N_2840_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_ns_LC_19_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_ns_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_ns_LC_19_19_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_ns_LC_19_19_4  (
            .in0(_gnd_net_),
            .in1(N__35553),
            .in2(N__28435),
            .in3(N__28597),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m5_d_LC_19_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m5_d_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m5_d_LC_19_19_5 .LUT_INIT=16'b0101110011000101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m5_d_LC_19_19_5  (
            .in0(N__35517),
            .in1(N__28936),
            .in2(N__27745),
            .in3(N__29003),
            .lcout(\this_vga_signals.if_m5_d ),
            .ltout(\this_vga_signals.if_m5_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_19_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_19_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_19_19_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_18_LC_19_19_6  (
            .in0(N__28651),
            .in1(N__28855),
            .in2(N__27736),
            .in3(N__27844),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_1_LC_19_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_1_LC_19_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_1_LC_19_19_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_1_LC_19_19_7  (
            .in0(N__27909),
            .in1(N__35684),
            .in2(_gnd_net_),
            .in3(N__27945),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIS9T25_0_9_LC_19_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIS9T25_0_9_LC_19_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIS9T25_0_9_LC_19_20_0 .LUT_INIT=16'b1001001101101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIS9T25_0_9_LC_19_20_0  (
            .in0(N__28030),
            .in1(N__27914),
            .in2(N__27990),
            .in3(N__28785),
            .lcout(\this_vga_signals.N_27_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_LC_19_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_LC_19_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_LC_19_20_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_LC_19_20_1  (
            .in0(N__27787),
            .in1(N__28425),
            .in2(_gnd_net_),
            .in3(N__28516),
            .lcout(\this_vga_signals.g0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNICUI21_LC_19_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNICUI21_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNICUI21_LC_19_20_2 .LUT_INIT=16'b1100100110011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNICUI21_LC_19_20_2  (
            .in0(N__34716),
            .in1(N__35146),
            .in2(N__35300),
            .in3(N__28201),
            .lcout(\this_vga_signals.vaddress_7 ),
            .ltout(\this_vga_signals.vaddress_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIS9T25_9_LC_19_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIS9T25_9_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIS9T25_9_LC_19_20_3 .LUT_INIT=16'b1001011001001011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIS9T25_9_LC_19_20_3  (
            .in0(N__28784),
            .in1(N__27982),
            .in2(N__27832),
            .in3(N__28029),
            .lcout(\this_vga_signals.N_27_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_N_3_i_LC_19_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_N_3_i_LC_19_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_N_3_i_LC_19_20_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_N_3_i_LC_19_20_4  (
            .in0(N__28456),
            .in1(N__27829),
            .in2(N__27816),
            .in3(N__28858),
            .lcout(),
            .ltout(\this_vga_signals.g1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_19_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_19_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_19_20_5 .LUT_INIT=16'b1101011100101000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_9_LC_19_20_5  (
            .in0(N__28603),
            .in1(N__28792),
            .in2(N__27799),
            .in3(N__28828),
            .lcout(\this_vga_signals.if_m6_i_x2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA65T2_9_LC_19_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA65T2_9_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA65T2_9_LC_19_21_1 .LUT_INIT=16'b0000000100000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIA65T2_9_LC_19_21_1  (
            .in0(N__30429),
            .in1(N__28359),
            .in2(N__28031),
            .in3(_gnd_net_),
            .lcout(N_842_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_19_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_19_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_19_21_3 .LUT_INIT=16'b1001111010100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_3_LC_19_21_3  (
            .in0(N__27964),
            .in1(N__27915),
            .in2(N__35013),
            .in3(N__27958),
            .lcout(\this_vga_signals.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_19_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_19_21_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_32_LC_19_21_4  (
            .in0(_gnd_net_),
            .in1(N__35460),
            .in2(_gnd_net_),
            .in3(N__28909),
            .lcout(\this_vga_signals.g0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_6_LC_19_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_6_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_6_LC_19_21_5 .LUT_INIT=16'b1100110011001001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI65531_6_LC_19_21_5  (
            .in0(N__30540),
            .in1(N__30670),
            .in2(N__35155),
            .in3(N__34745),
            .lcout(\this_vga_signals.vaddress_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_1_9_LC_19_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_1_9_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_1_9_LC_19_21_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_1_9_LC_19_21_6  (
            .in0(N__30571),
            .in1(N__30428),
            .in2(_gnd_net_),
            .in3(N__30539),
            .lcout(this_vga_signals_CO0_0_i_i),
            .ltout(this_vga_signals_CO0_0_i_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGBA04_9_LC_19_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGBA04_9_LC_19_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGBA04_9_LC_19_21_7 .LUT_INIT=16'b0011110011001111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGBA04_9_LC_19_21_7  (
            .in0(_gnd_net_),
            .in1(N__28786),
            .in2(N__27994),
            .in3(N__27989),
            .lcout(\this_vga_signals.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_3_LC_19_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_3_LC_19_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_3_LC_19_22_6 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_3_LC_19_22_6  (
            .in0(N__35286),
            .in1(N__27957),
            .in2(N__27919),
            .in3(N__34746),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_38_i_0_a2_0_4_1_LC_19_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.N_38_i_0_a2_0_4_1_LC_19_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_38_i_0_a2_0_4_1_LC_19_23_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.N_38_i_0_a2_0_4_1_LC_19_23_0  (
            .in0(_gnd_net_),
            .in1(N__30833),
            .in2(_gnd_net_),
            .in3(N__28164),
            .lcout(\this_vga_signals.N_38_i_0_a2_0_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_17_LC_19_23_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_17_LC_19_23_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_17_LC_19_23_1 .LUT_INIT=16'b0101000101110011;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_1_17_LC_19_23_1  (
            .in0(N__29222),
            .in1(N__27873),
            .in2(N__29206),
            .in3(N__43355),
            .lcout(),
            .ltout(\this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_17_LC_19_23_2.C_ON=1'b0;
    defparam M_this_state_q_17_LC_19_23_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_17_LC_19_23_2.LUT_INIT=16'b1000100000001100;
    LogicCell40 M_this_state_q_17_LC_19_23_2 (
            .in0(N__43356),
            .in1(N__29062),
            .in2(N__27877),
            .in3(N__28166),
            .lcout(M_this_state_qZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42068),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQ6821_8_LC_19_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQ6821_8_LC_19_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQ6821_8_LC_19_23_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIQ6821_8_LC_19_23_3  (
            .in0(N__30693),
            .in1(N__30457),
            .in2(_gnd_net_),
            .in3(N__35152),
            .lcout(\this_vga_signals.vsync_1_0_a3_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam led_1_7_5__m12_0_a3_0_a3_0_o2_LC_19_23_5.C_ON=1'b0;
    defparam led_1_7_5__m12_0_a3_0_a3_0_o2_LC_19_23_5.SEQ_MODE=4'b0000;
    defparam led_1_7_5__m12_0_a3_0_a3_0_o2_LC_19_23_5.LUT_INIT=16'b0000000000010001;
    LogicCell40 led_1_7_5__m12_0_a3_0_a3_0_o2_LC_19_23_5 (
            .in0(N__29221),
            .in1(N__36099),
            .in2(_gnd_net_),
            .in3(N__29271),
            .lcout(N_773_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_4_LC_19_23_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_4_LC_19_23_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_4_LC_19_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a3_4_LC_19_23_6  (
            .in0(_gnd_net_),
            .in1(N__31034),
            .in2(_gnd_net_),
            .in3(N__38587),
            .lcout(\this_ppu.N_1162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_this_state_q_8_0_i_0_0_i_LC_19_23_7 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_state_q_8_0_i_0_0_i_LC_19_23_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_state_q_8_0_i_0_0_i_LC_19_23_7 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \this_ppu.un1_M_this_state_q_8_0_i_0_0_i_LC_19_23_7  (
            .in0(N__28165),
            .in1(N__43354),
            .in2(N__36532),
            .in3(N__30836),
            .lcout(N_247),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_19_24_0.C_ON=1'b0;
    defparam M_this_state_q_7_LC_19_24_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_19_24_0.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_7_LC_19_24_0 (
            .in0(N__30296),
            .in1(N__31054),
            .in2(N__29116),
            .in3(N__29046),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42079),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_8_LC_19_24_2.C_ON=1'b0;
    defparam M_this_state_q_8_LC_19_24_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_8_LC_19_24_2.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_8_LC_19_24_2 (
            .in0(N__30297),
            .in1(N__31055),
            .in2(N__29101),
            .in3(N__30928),
            .lcout(M_this_state_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42079),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_q_0_i_0_o2_1_LC_19_24_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_o2_1_LC_19_24_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_o2_1_LC_19_24_7 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_o2_1_LC_19_24_7  (
            .in0(N__43365),
            .in1(N__36354),
            .in2(_gnd_net_),
            .in3(N__38586),
            .lcout(N_794_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0_LC_19_25_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0_LC_19_25_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0_LC_19_25_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_ppu.M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0_LC_19_25_5  (
            .in0(_gnd_net_),
            .in1(N__43234),
            .in2(_gnd_net_),
            .in3(N__36113),
            .lcout(this_ppu_M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_a2_3_LC_19_26_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_a2_3_LC_19_26_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_a2_3_LC_19_26_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_1_0_a2_3_LC_19_26_2  (
            .in0(N__36513),
            .in1(N__43401),
            .in2(_gnd_net_),
            .in3(N__36444),
            .lcout(\this_ppu.N_1322 ),
            .ltout(\this_ppu.N_1322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_0_LC_19_26_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_0_LC_19_26_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_0_LC_19_26_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_1_0_i_0_LC_19_26_3  (
            .in0(N__42444),
            .in1(N__40751),
            .in2(N__28129),
            .in3(N__36514),
            .lcout(M_this_spr_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_0_6_LC_20_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_0_6_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_0_6_LC_20_17_0 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI65531_0_6_LC_20_17_0  (
            .in0(N__30684),
            .in1(N__34704),
            .in2(N__35154),
            .in3(N__30502),
            .lcout(\this_vga_signals.N_1247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_0_LC_20_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_0_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_0_LC_20_17_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_0_LC_20_17_1  (
            .in0(N__28270),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28231),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_2_LC_20_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_2_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_2_LC_20_17_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_2_LC_20_17_2  (
            .in0(N__30683),
            .in1(N__34703),
            .in2(N__28336),
            .in3(N__30501),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_20_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_20_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_20_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_20_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28333),
            .lcout(this_vga_signals_M_vcounter_q_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42021),
            .ce(N__34249),
            .sr(N__34218));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_20_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_20_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_20_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_9_LC_20_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28300),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42021),
            .ce(N__34249),
            .sr(N__34218));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_1_1_LC_20_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_1_1_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_1_1_LC_20_17_5 .LUT_INIT=16'b0001100010000111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_1_1_LC_20_17_5  (
            .in0(N__28269),
            .in1(N__28230),
            .in2(N__28260),
            .in3(N__28215),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_0_1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_20_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_20_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_20_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_20_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30766),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42021),
            .ce(N__34249),
            .sr(N__34218));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_20_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_20_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_20_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_20_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30730),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42021),
            .ce(N__34249),
            .sr(N__34218));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_20_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_20_18_0 .LUT_INIT=16'b0111100010000111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_20_18_0  (
            .in0(N__28693),
            .in1(N__28769),
            .in2(N__35293),
            .in3(N__28200),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_20_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_20_18_1 .LUT_INIT=16'b0100011011001111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_20_18_1  (
            .in0(N__34971),
            .in1(N__35240),
            .in2(N__28171),
            .in3(N__34123),
            .lcout(\this_vga_signals.mult1_un54_sum_c2_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_20_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_20_18_2 .LUT_INIT=16'b0010101111010100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_LC_20_18_2  (
            .in0(N__34039),
            .in1(N__28444),
            .in2(N__28459),
            .in3(N__30037),
            .lcout(\this_vga_signals.g0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_20_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_20_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_20_18_3  (
            .in0(_gnd_net_),
            .in1(N__35602),
            .in2(_gnd_net_),
            .in3(N__34070),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_20_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_20_18_4 .LUT_INIT=16'b0110100101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_29_LC_20_18_4  (
            .in0(N__30073),
            .in1(N__29488),
            .in2(N__28447),
            .in3(N__29531),
            .lcout(\this_vga_signals.mult1_un47_sum_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_20_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_20_18_5 .LUT_INIT=16'b0110100110100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_20_18_5  (
            .in0(N__35663),
            .in1(N__35603),
            .in2(N__35705),
            .in3(N__34071),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc1 ),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x1_LC_20_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x1_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x1_LC_20_18_6 .LUT_INIT=16'b0010111100001010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x1_LC_20_18_6  (
            .in0(N__35241),
            .in1(N__34972),
            .in2(N__28438),
            .in3(N__34131),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_20_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_20_18_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_1_LC_20_18_7  (
            .in0(N__34132),
            .in1(N__30028),
            .in2(_gnd_net_),
            .in3(N__29987),
            .lcout(\this_vga_signals.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_20_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_20_19_0 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_20_19_0  (
            .in0(N__30017),
            .in1(N__29982),
            .in2(N__34137),
            .in3(N__35384),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_20_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_20_19_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_20_19_1  (
            .in0(N__35317),
            .in1(_gnd_net_),
            .in2(N__35405),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_LC_20_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_LC_20_19_2 .LUT_INIT=16'b1000101000100010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_LC_20_19_2  (
            .in0(N__28426),
            .in1(N__28387),
            .in2(N__34946),
            .in3(N__28369),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x0_LC_20_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x0_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x0_LC_20_19_3 .LUT_INIT=16'b0111101100110011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x0_LC_20_19_3  (
            .in0(N__35315),
            .in1(N__30016),
            .in2(N__34944),
            .in3(N__34125),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_3_1_LC_20_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_3_1_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_3_1_LC_20_19_4 .LUT_INIT=16'b0111100000011110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_3_1_LC_20_19_4  (
            .in0(N__34130),
            .in1(N__29983),
            .in2(N__28947),
            .in3(N__35566),
            .lcout(\this_vga_signals.g0_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m3_i_m2_LC_20_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m3_i_m2_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m3_i_m2_LC_20_19_5 .LUT_INIT=16'b0010111000111100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m3_i_m2_LC_20_19_5  (
            .in0(N__35316),
            .in1(N__34152),
            .in2(N__34945),
            .in3(N__34126),
            .lcout(),
            .ltout(\this_vga_signals.if_N_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m3_LC_20_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m3_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m3_LC_20_19_6 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m3_LC_20_19_6  (
            .in0(N__35514),
            .in1(N__35552),
            .in2(N__28591),
            .in3(N__35380),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_d ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_20_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_20_19_7 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_20_19_7  (
            .in0(N__28588),
            .in1(N__28539),
            .in2(N__28564),
            .in3(N__30079),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_20_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_20_20_0 .LUT_INIT=16'b1100011001100011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_15_LC_20_20_0  (
            .in0(N__30031),
            .in1(N__35400),
            .in2(N__28561),
            .in3(N__29989),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_20_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_20_20_1 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_LC_20_20_1  (
            .in0(N__28549),
            .in1(N__28540),
            .in2(N__28528),
            .in3(N__28517),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_20_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_20_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_LC_20_20_2  (
            .in0(N__30196),
            .in1(N__29014),
            .in2(N__28492),
            .in3(N__28489),
            .lcout(\this_vga_signals.N_3_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_20_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_20_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_LC_20_20_3  (
            .in0(N__35399),
            .in1(N__28648),
            .in2(N__28474),
            .in3(N__28982),
            .lcout(\this_vga_signals.g0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_20_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_20_20_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_0_LC_20_20_4  (
            .in0(N__29007),
            .in1(_gnd_net_),
            .in2(N__28987),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_c2_LC_20_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_c2_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_c2_LC_20_20_5 .LUT_INIT=16'b1101010001110001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_c2_LC_20_20_5  (
            .in0(N__28948),
            .in1(N__28649),
            .in2(N__35521),
            .in3(N__28857),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_3_LC_20_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_3_LC_20_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_3_LC_20_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_3_LC_20_20_6  (
            .in0(N__35323),
            .in1(N__35401),
            .in2(N__28837),
            .in3(N__28834),
            .lcout(\this_vga_signals.g0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_20_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_20_21_0 .LUT_INIT=16'b1001111100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_LC_20_21_0  (
            .in0(N__35410),
            .in1(N__28822),
            .in2(N__28813),
            .in3(N__28798),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_20_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_20_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_LC_20_21_1  (
            .in0(_gnd_net_),
            .in1(N__28713),
            .in2(_gnd_net_),
            .in3(N__28770),
            .lcout(\this_vga_signals.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_9_LC_20_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_9_LC_20_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_9_LC_20_21_3 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_9_LC_20_21_3  (
            .in0(N__30455),
            .in1(N__30567),
            .in2(_gnd_net_),
            .in3(N__30533),
            .lcout(\this_vga_signals.vaddress_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_1_LC_20_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_1_LC_20_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_1_LC_20_21_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_x2_1_LC_20_21_4  (
            .in0(N__28771),
            .in1(_gnd_net_),
            .in2(N__28717),
            .in3(N__34986),
            .lcout(\this_vga_signals.N_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_LC_20_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_LC_20_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_LC_20_21_5 .LUT_INIT=16'b1001111101101111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_LC_20_21_5  (
            .in0(N__35489),
            .in1(N__28665),
            .in2(N__28618),
            .in3(N__30211),
            .lcout(\this_vga_signals.if_m5_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_1_LC_20_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_1_LC_20_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_1_LC_20_22_1 .LUT_INIT=16'b0011001110010011;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_1_LC_20_22_1  (
            .in0(N__35322),
            .in1(N__35099),
            .in2(N__35005),
            .in3(N__34747),
            .lcout(\this_vga_signals.g1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1_0_LC_20_22_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1_0_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1_0_LC_20_22_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1_0_LC_20_22_3  (
            .in0(N__30929),
            .in1(N__30887),
            .in2(_gnd_net_),
            .in3(N__43224),
            .lcout(\this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_16_LC_20_22_5.C_ON=1'b0;
    defparam M_this_state_q_16_LC_20_22_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_16_LC_20_22_5.LUT_INIT=16'b1111000010000000;
    LogicCell40 M_this_state_q_16_LC_20_22_5 (
            .in0(N__29143),
            .in1(N__29089),
            .in2(N__31090),
            .in3(N__30838),
            .lcout(M_this_state_qZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42069),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_2_15_LC_20_22_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_2_15_LC_20_22_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_2_15_LC_20_22_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_2_15_LC_20_22_6  (
            .in0(N__43225),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35784),
            .lcout(\this_ppu.N_235_2_0 ),
            .ltout(\this_ppu.N_235_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_0_15_LC_20_22_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_0_15_LC_20_22_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_0_15_LC_20_22_7 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_0_15_LC_20_22_7  (
            .in0(N__29142),
            .in1(N__43471),
            .in2(N__29056),
            .in3(N__30837),
            .lcout(\this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_1_LC_20_23_0.C_ON=1'b0;
    defparam M_this_state_q_1_LC_20_23_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_20_23_0.LUT_INIT=16'b1111100010001000;
    LogicCell40 M_this_state_q_1_LC_20_23_0 (
            .in0(N__40862),
            .in1(N__31067),
            .in2(N__29449),
            .in3(N__30969),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42080),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_10_LC_20_23_2.C_ON=1'b0;
    defparam M_this_state_q_10_LC_20_23_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_10_LC_20_23_2.LUT_INIT=16'b1110101011000000;
    LogicCell40 M_this_state_q_10_LC_20_23_2 (
            .in0(N__31137),
            .in1(N__31065),
            .in2(N__36114),
            .in3(N__33015),
            .lcout(M_this_state_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42080),
            .ce(),
            .sr(_gnd_net_));
    defparam led_1_7_5__m17_0_a3_0_a3_0_o2_LC_20_23_3.C_ON=1'b0;
    defparam led_1_7_5__m17_0_a3_0_a3_0_o2_LC_20_23_3.SEQ_MODE=4'b0000;
    defparam led_1_7_5__m17_0_a3_0_a3_0_o2_LC_20_23_3.LUT_INIT=16'b0000000000010001;
    LogicCell40 led_1_7_5__m17_0_a3_0_a3_0_o2_LC_20_23_3 (
            .in0(N__40861),
            .in1(N__29042),
            .in2(_gnd_net_),
            .in3(N__37386),
            .lcout(N_815_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_20_23_4.C_ON=1'b0;
    defparam M_this_state_q_4_LC_20_23_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_20_23_4.LUT_INIT=16'b1110101010101010;
    LogicCell40 M_this_state_q_4_LC_20_23_4 (
            .in0(N__29020),
            .in1(N__36160),
            .in2(N__32866),
            .in3(N__30793),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42080),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_9_LC_20_23_5.C_ON=1'b0;
    defparam M_this_state_q_9_LC_20_23_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_9_LC_20_23_5.LUT_INIT=16'b1010111000001100;
    LogicCell40 M_this_state_q_9_LC_20_23_5 (
            .in0(N__31068),
            .in1(N__31138),
            .in2(N__33022),
            .in3(N__29281),
            .lcout(M_this_state_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42080),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_11_LC_20_23_6.C_ON=1'b0;
    defparam M_this_state_q_11_LC_20_23_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_11_LC_20_23_6.LUT_INIT=16'b1111100010001000;
    LogicCell40 M_this_state_q_11_LC_20_23_6 (
            .in0(N__29107),
            .in1(N__30792),
            .in2(N__29244),
            .in3(N__31066),
            .lcout(M_this_state_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42080),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_15_LC_20_23_7.C_ON=1'b0;
    defparam M_this_state_q_15_LC_20_23_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_15_LC_20_23_7.LUT_INIT=16'b0100000011001100;
    LogicCell40 M_this_state_q_15_LC_20_23_7 (
            .in0(N__29205),
            .in1(N__29161),
            .in2(N__29151),
            .in3(N__37455),
            .lcout(M_this_state_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42080),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_7_LC_20_24_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_7_LC_20_24_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_7_LC_20_24_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_7_LC_20_24_0  (
            .in0(N__36154),
            .in1(N__36298),
            .in2(_gnd_net_),
            .in3(N__35846),
            .lcout(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_0_0_LC_20_24_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_0_0_LC_20_24_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_0_0_LC_20_24_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_0_a2_0_0_LC_20_24_2  (
            .in0(N__42616),
            .in1(N__35777),
            .in2(N__29445),
            .in3(N__43235),
            .lcout(\this_ppu.N_1425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_11_LC_20_24_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_11_LC_20_24_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_11_LC_20_24_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_11_LC_20_24_3  (
            .in0(N__32927),
            .in1(N__33013),
            .in2(_gnd_net_),
            .in3(N__33088),
            .lcout(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_8_LC_20_24_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_8_LC_20_24_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_8_LC_20_24_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_8_LC_20_24_4  (
            .in0(N__36155),
            .in1(N__36299),
            .in2(_gnd_net_),
            .in3(N__35847),
            .lcout(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_o2_6_LC_20_24_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_o2_6_LC_20_24_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_o2_6_LC_20_24_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_o2_6_LC_20_24_6  (
            .in0(N__33089),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32928),
            .lcout(\this_ppu.N_807_0 ),
            .ltout(\this_ppu.N_807_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_this_state_q_11_0_0_m3_LC_20_24_7 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_state_q_11_0_0_m3_LC_20_24_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_state_q_11_0_0_m3_LC_20_24_7 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \this_ppu.un1_M_this_state_q_11_0_0_m3_LC_20_24_7  (
            .in0(N__36300),
            .in1(N__33014),
            .in2(N__29092),
            .in3(N__36242),
            .lcout(\this_ppu.N_969 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_2_LC_20_25_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_2_LC_20_25_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_2_LC_20_25_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_2_LC_20_25_2  (
            .in0(N__32981),
            .in1(N__33091),
            .in2(_gnd_net_),
            .in3(N__32935),
            .lcout(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a2_0_1_LC_20_25_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a2_0_1_LC_20_25_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a2_0_1_LC_20_25_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a2_0_1_LC_20_25_3  (
            .in0(N__32934),
            .in1(N__32980),
            .in2(N__36210),
            .in3(N__33090),
            .lcout(\this_ppu.N_1341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_2_LC_20_26_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_2_LC_20_26_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_2_LC_20_26_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_1_0_i_2_LC_20_26_2  (
            .in0(N__42773),
            .in1(N__35976),
            .in2(N__40436),
            .in3(N__36531),
            .lcout(M_this_spr_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_5_LC_21_15_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_5_LC_21_15_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_5_LC_21_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_5_LC_21_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29341),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42011),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_21_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_21_17_0 .LUT_INIT=16'b1101010000101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_20_LC_21_17_0  (
            .in0(N__30030),
            .in1(N__29980),
            .in2(N__29299),
            .in3(N__35407),
            .lcout(\this_vga_signals.mult1_un54_sum_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_a3_0_LC_21_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_a3_0_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_a3_0_LC_21_17_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_a3_0_LC_21_17_1  (
            .in0(_gnd_net_),
            .in1(N__35320),
            .in2(_gnd_net_),
            .in3(N__35548),
            .lcout(\this_vga_signals.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_21_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_21_17_2 .LUT_INIT=16'b0101100110100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_11_LC_21_17_2  (
            .in0(N__30108),
            .in1(N__29527),
            .in2(N__29490),
            .in3(N__29571),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_21_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_21_17_3 .LUT_INIT=16'b1011001100110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_8_LC_21_17_3  (
            .in0(N__34186),
            .in1(N__34174),
            .in2(N__29308),
            .in3(N__29305),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_21_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_21_17_4 .LUT_INIT=16'b0100101110110100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_23_LC_21_17_4  (
            .in0(N__29480),
            .in1(N__29523),
            .in2(N__29776),
            .in3(N__29569),
            .lcout(\this_vga_signals.mult1_un47_sum_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_21_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_21_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_21_17_5 .LUT_INIT=16'b0110010110011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_28_LC_21_17_5  (
            .in0(N__29570),
            .in1(N__29481),
            .in2(N__29532),
            .in3(N__30107),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_21_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_21_17_6 .LUT_INIT=16'b1101010000101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_38_LC_21_17_6  (
            .in0(N__30029),
            .in1(N__29981),
            .in2(N__29806),
            .in3(N__35406),
            .lcout(\this_vga_signals.mult1_un54_sum_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_3_0_LC_21_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_3_0_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_3_0_LC_21_17_7 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_3_0_LC_21_17_7  (
            .in0(N__29880),
            .in1(N__29843),
            .in2(N__29937),
            .in3(N__29642),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_0_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_0_LC_21_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_0_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_o2_0_LC_21_18_0 .LUT_INIT=16'b1010000010100001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_o2_0_LC_21_18_0  (
            .in0(N__30688),
            .in1(N__34706),
            .in2(N__35136),
            .in3(N__30520),
            .lcout(\this_ppu.m18_i_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_21_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_21_18_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_25_LC_21_18_1  (
            .in0(N__34069),
            .in1(_gnd_net_),
            .in2(N__35616),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_5_LC_21_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_5_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_5_LC_21_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_5_LC_21_18_2  (
            .in0(_gnd_net_),
            .in1(N__29767),
            .in2(_gnd_net_),
            .in3(N__29719),
            .lcout(N_814_0),
            .ltout(N_814_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_1_LC_21_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_1_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_1_LC_21_18_3 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_1_LC_21_18_3  (
            .in0(N__29665),
            .in1(N__29659),
            .in2(N__29647),
            .in3(N__29635),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc3_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_2_LC_21_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_2_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_2_LC_21_18_4 .LUT_INIT=16'b1110000001110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_2_LC_21_18_4  (
            .in0(N__35100),
            .in1(N__30421),
            .in2(N__29578),
            .in3(N__30669),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_2_2 ),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc3_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_21_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_21_18_5 .LUT_INIT=16'b1100111100110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_21_18_5  (
            .in0(_gnd_net_),
            .in1(N__29476),
            .in2(N__29575),
            .in3(N__29557),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_21_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_21_18_6 .LUT_INIT=16'b0101100110100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_21_18_6  (
            .in0(N__29558),
            .in1(N__29522),
            .in2(N__29489),
            .in3(N__34068),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc3_x1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_21_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_21_18_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_21_18_7  (
            .in0(N__35604),
            .in1(_gnd_net_),
            .in2(N__30133),
            .in3(N__30130),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_21_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_21_19_0 .LUT_INIT=16'b0111000111110101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_21_19_0  (
            .in0(N__35656),
            .in1(N__35609),
            .in2(N__35713),
            .in3(N__34072),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_21_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_21_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_21_19_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_21_19_1  (
            .in0(N__30124),
            .in1(N__30103),
            .in2(N__30085),
            .in3(N__34118),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_21_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_21_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_21_19_2 .LUT_INIT=16'b1011010000101101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_21_19_2  (
            .in0(N__34119),
            .in1(N__30018),
            .in2(N__30082),
            .in3(N__29978),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_1_LC_21_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_1_LC_21_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_1_LC_21_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_1_LC_21_19_3  (
            .in0(N__30072),
            .in1(N__34880),
            .in2(N__30052),
            .in3(N__35386),
            .lcout(\this_vga_signals.g0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_2_LC_21_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_2_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_2_LC_21_19_4 .LUT_INIT=16'b0101100110011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_x2_2_LC_21_19_4  (
            .in0(N__35385),
            .in1(N__30019),
            .in2(N__34136),
            .in3(N__29979),
            .lcout(\this_vga_signals.N_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_LC_21_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_LC_21_19_5 .LUT_INIT=16'b1110110001110011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_LC_21_19_5  (
            .in0(N__29851),
            .in1(N__29938),
            .in2(N__29902),
            .in3(N__29887),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_3_LC_21_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_3_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_3_LC_21_19_6 .LUT_INIT=16'b1101111100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_3_LC_21_19_6  (
            .in0(N__29886),
            .in1(N__29850),
            .in2(N__30186),
            .in3(N__30156),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_3 ),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb1_LC_21_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb1_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb1_LC_21_19_7 .LUT_INIT=16'b1010000001011111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb1_LC_21_19_7  (
            .in0(N__35608),
            .in1(_gnd_net_),
            .in2(N__30280),
            .in3(N__35709),
            .lcout(\this_vga_signals.mult1_un47_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIPMQM_6_LC_21_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIPMQM_6_LC_21_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIPMQM_6_LC_21_20_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIPMQM_6_LC_21_20_0  (
            .in0(N__35089),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34748),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_8_LC_21_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_8_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_8_LC_21_20_1 .LUT_INIT=16'b0010001101010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_8_LC_21_20_1  (
            .in0(N__30534),
            .in1(N__30459),
            .in2(N__30277),
            .in3(N__30651),
            .lcout(\this_vga_signals.N_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3GK81_0_8_LC_21_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3GK81_0_8_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3GK81_0_8_LC_21_20_2 .LUT_INIT=16'b1010001011011011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI3GK81_0_8_LC_21_20_2  (
            .in0(N__30652),
            .in1(N__30274),
            .in2(N__35133),
            .in3(N__30458),
            .lcout(\this_vga_signals.N_39_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_21_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_21_20_3 .LUT_INIT=16'b0011100011100111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_26_LC_21_20_3  (
            .in0(N__30240),
            .in1(N__34879),
            .in2(N__34633),
            .in3(N__30259),
            .lcout(),
            .ltout(\this_vga_signals.g1_3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_LC_21_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_LC_21_20_4 .LUT_INIT=16'b0110111111111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_LC_21_20_4  (
            .in0(N__30250),
            .in1(N__30241),
            .in2(N__30229),
            .in3(N__35304),
            .lcout(),
            .ltout(\this_vga_signals.g3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_21_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_21_20_5 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_13_LC_21_20_5  (
            .in0(N__30226),
            .in1(N__35329),
            .in2(N__30220),
            .in3(N__30217),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_21_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_21_20_6 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_21_20_6  (
            .in0(N__35305),
            .in1(N__35398),
            .in2(N__35520),
            .in3(N__30205),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_1_0_LC_21_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_1_0_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_1_0_LC_21_21_0 .LUT_INIT=16'b0000100011111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_1_0_LC_21_21_0  (
            .in0(N__30638),
            .in1(N__30187),
            .in2(N__35135),
            .in3(N__30157),
            .lcout(\this_vga_signals.g2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_21_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_21_21_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_21_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_21_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30755),
            .lcout(this_vga_signals_M_vcounter_q_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42070),
            .ce(N__34252),
            .sr(N__34221));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_21_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_21_21_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_21_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_21_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30726),
            .lcout(this_vga_signals_M_vcounter_q_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42070),
            .ce(N__34252),
            .sr(N__34221));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIN3821_6_LC_21_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIN3821_6_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIN3821_6_LC_21_21_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIN3821_6_LC_21_21_3  (
            .in0(N__35075),
            .in1(N__30637),
            .in2(_gnd_net_),
            .in3(N__34744),
            .lcout(N_1001_0),
            .ltout(N_1001_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_0_9_LC_21_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_0_9_LC_21_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_0_9_LC_21_21_4 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_0_9_LC_21_21_4  (
            .in0(_gnd_net_),
            .in1(N__30532),
            .in2(N__30475),
            .in3(N__30456),
            .lcout(\this_vga_signals.g4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_3_15_LC_21_22_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_3_15_LC_21_22_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_3_15_LC_21_22_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_o2_3_15_LC_21_22_1  (
            .in0(_gnd_net_),
            .in1(N__30835),
            .in2(_gnd_net_),
            .in3(N__36100),
            .lcout(\this_ppu.N_856_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a2_3_LC_21_22_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a2_3_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a2_3_LC_21_22_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a2_3_LC_21_22_2  (
            .in0(N__36000),
            .in1(N__36307),
            .in2(N__36250),
            .in3(N__35840),
            .lcout(\this_ppu.N_1278 ),
            .ltout(\this_ppu.N_1278_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_3_LC_21_22_3.C_ON=1'b0;
    defparam M_this_state_q_3_LC_21_22_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_21_22_3.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_3_LC_21_22_3 (
            .in0(N__31129),
            .in1(N__31089),
            .in2(N__30319),
            .in3(N__36343),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42081),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_0_a3_0_LC_21_22_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a3_0_LC_21_22_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a3_0_LC_21_22_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_0_a3_0_LC_21_22_4  (
            .in0(N__36001),
            .in1(N__36306),
            .in2(N__31123),
            .in3(N__30315),
            .lcout(),
            .ltout(\this_ppu.N_1149_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_0_LC_21_22_5.C_ON=1'b0;
    defparam M_this_state_q_0_LC_21_22_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_0_LC_21_22_5.LUT_INIT=16'b0000101100001010;
    LogicCell40 M_this_state_q_0_LC_21_22_5 (
            .in0(N__30316),
            .in1(N__30301),
            .in2(N__30283),
            .in3(N__30943),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42081),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_0_0_tz_0_LC_21_22_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_0_0_tz_0_LC_21_22_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_0_0_tz_0_LC_21_22_6 .LUT_INIT=16'b0011111100010101;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_0_0_tz_0_LC_21_22_6  (
            .in0(N__31088),
            .in1(N__35793),
            .in2(N__30955),
            .in3(N__35841),
            .lcout(\this_ppu.M_this_state_q_srsts_0_0_0_tz_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam led_1_7_5__m17_0_a3_0_a3_0_a3_LC_21_22_7.C_ON=1'b0;
    defparam led_1_7_5__m17_0_a3_0_a3_0_a3_LC_21_22_7.SEQ_MODE=4'b0000;
    defparam led_1_7_5__m17_0_a3_0_a3_0_a3_LC_21_22_7.LUT_INIT=16'b0100000001000000;
    LogicCell40 led_1_7_5__m17_0_a3_0_a3_0_a3_LC_21_22_7 (
            .in0(N__30937),
            .in1(N__30888),
            .in2(N__35797),
            .in3(_gnd_net_),
            .lcout(led_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_6_LC_21_23_0.C_ON=1'b0;
    defparam M_this_state_q_6_LC_21_23_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_21_23_0.LUT_INIT=16'b1111111110000000;
    LogicCell40 M_this_state_q_6_LC_21_23_0 (
            .in0(N__30791),
            .in1(N__33020),
            .in2(N__30847),
            .in3(N__30775),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42091),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_0_sqmuxa_i_i_o3_0_a2_LC_21_23_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_0_sqmuxa_i_i_o3_0_a2_LC_21_23_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_0_sqmuxa_i_i_o3_0_a2_LC_21_23_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_0_sqmuxa_i_i_o3_0_a2_LC_21_23_1  (
            .in0(_gnd_net_),
            .in1(N__30834),
            .in2(_gnd_net_),
            .in3(N__38275),
            .lcout(N_1415),
            .ltout(N_1415_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_0_sqmuxa_i_i_o3_0_o3_LC_21_23_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_0_sqmuxa_i_i_o3_0_o3_LC_21_23_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_0_sqmuxa_i_i_o3_0_o3_LC_21_23_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_0_sqmuxa_i_i_o3_0_o3_LC_21_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30796),
            .in3(N__43460),
            .lcout(N_296_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_5_LC_21_23_3.C_ON=1'b0;
    defparam M_this_state_q_5_LC_21_23_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_21_23_3.LUT_INIT=16'b1110101011000000;
    LogicCell40 M_this_state_q_5_LC_21_23_3 (
            .in0(N__31064),
            .in1(N__30790),
            .in2(N__30994),
            .in3(N__37387),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42091),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_6_LC_21_23_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_6_LC_21_23_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_6_LC_21_23_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a3_6_LC_21_23_4  (
            .in0(N__38276),
            .in1(N__31063),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.N_1166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a2_1_LC_21_23_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a2_1_LC_21_23_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a2_1_LC_21_23_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a2_1_LC_21_23_5  (
            .in0(N__34486),
            .in1(N__43756),
            .in2(N__36287),
            .in3(N__35839),
            .lcout(\this_ppu.N_1263 ),
            .ltout(\this_ppu.N_1263_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_1_10_LC_21_23_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_1_10_LC_21_23_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_1_10_LC_21_23_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a3_0_1_10_LC_21_23_6  (
            .in0(N__33052),
            .in1(N__36243),
            .in2(N__30769),
            .in3(N__32932),
            .lcout(\this_ppu.N_1176_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_3_LC_21_23_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_3_LC_21_23_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_3_LC_21_23_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_3_LC_21_23_7  (
            .in0(N__33021),
            .in1(N__33051),
            .in2(N__32942),
            .in3(N__36153),
            .lcout(\this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_0_m2_0_LC_21_24_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_0_m2_0_LC_21_24_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_0_m2_0_LC_21_24_0 .LUT_INIT=16'b1111010110000010;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_0_m2_0_LC_21_24_0  (
            .in0(N__33019),
            .in1(N__36226),
            .in2(N__33087),
            .in3(N__32933),
            .lcout(\this_ppu.N_893 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_this_state_q_11_0_0_LC_21_24_5 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_state_q_11_0_0_LC_21_24_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_state_q_11_0_0_LC_21_24_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_ppu.un1_M_this_state_q_11_0_0_LC_21_24_5  (
            .in0(N__42615),
            .in1(N__31096),
            .in2(N__31111),
            .in3(N__35773),
            .lcout(),
            .ltout(un1_M_this_state_q_11_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_LC_21_24_6.C_ON=1'b0;
    defparam M_this_substate_q_LC_21_24_6.SEQ_MODE=4'b1000;
    defparam M_this_substate_q_LC_21_24_6.LUT_INIT=16'b1010110000001100;
    LogicCell40 M_this_substate_q_LC_21_24_6 (
            .in0(N__32856),
            .in1(N__36156),
            .in2(N__31102),
            .in3(N__36124),
            .lcout(M_this_substate_qZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42100),
            .ce(),
            .sr(N__43106));
    defparam \this_ppu.un1_M_this_state_q_11_0_0_0_LC_21_25_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_state_q_11_0_0_0_LC_21_25_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_state_q_11_0_0_0_LC_21_25_0 .LUT_INIT=16'b0010111100000000;
    LogicCell40 \this_ppu.un1_M_this_state_q_11_0_0_0_LC_21_25_0  (
            .in0(N__32988),
            .in1(N__33074),
            .in2(N__32947),
            .in3(N__35845),
            .lcout(),
            .ltout(\this_ppu.un1_M_this_state_q_11_0_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_this_state_q_11_0_0_1_LC_21_25_1 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_state_q_11_0_0_1_LC_21_25_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_state_q_11_0_0_1_LC_21_25_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \this_ppu.un1_M_this_state_q_11_0_0_1_LC_21_25_1  (
            .in0(N__33075),
            .in1(N__32989),
            .in2(N__31099),
            .in3(N__36196),
            .lcout(\this_ppu.un1_M_this_state_q_11_0_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_2_LC_21_25_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_2_LC_21_25_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_a3_2_LC_21_25_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_a3_2_LC_21_25_3  (
            .in0(_gnd_net_),
            .in1(N__37781),
            .in2(_gnd_net_),
            .in3(N__31079),
            .lcout(),
            .ltout(\this_ppu.N_1158_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_2_LC_21_25_4.C_ON=1'b0;
    defparam M_this_state_q_2_LC_21_25_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_21_25_4.LUT_INIT=16'b1111010011110000;
    LogicCell40 M_this_state_q_2_LC_21_25_4 (
            .in0(N__36195),
            .in1(N__30990),
            .in2(N__30973),
            .in3(N__30970),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42108),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_substate_d_0_sqmuxa_3_0_a3_0_a2_LC_21_25_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_substate_d_0_sqmuxa_3_0_a3_0_a2_LC_21_25_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_substate_d_0_sqmuxa_3_0_a3_0_a2_LC_21_25_7 .LUT_INIT=16'b0000000100000001;
    LogicCell40 \this_ppu.M_this_substate_d_0_sqmuxa_3_0_a3_0_a2_LC_21_25_7  (
            .in0(N__33073),
            .in1(N__32987),
            .in2(N__32943),
            .in3(_gnd_net_),
            .lcout(N_1422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_spr_address_q_0_LC_22_14_0.C_ON=1'b1;
    defparam M_this_spr_address_q_0_LC_22_14_0.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_0_LC_22_14_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_0_LC_22_14_0 (
            .in0(N__33210),
            .in1(N__32661),
            .in2(N__36379),
            .in3(N__36378),
            .lcout(M_this_spr_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_22_14_0_),
            .carryout(un1_M_this_spr_address_q_cry_0),
            .clk(N__42012),
            .ce(),
            .sr(N__41653));
    defparam M_this_spr_address_q_1_LC_22_14_1.C_ON=1'b1;
    defparam M_this_spr_address_q_1_LC_22_14_1.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_1_LC_22_14_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_1_LC_22_14_1 (
            .in0(N__33214),
            .in1(N__32441),
            .in2(_gnd_net_),
            .in3(N__32398),
            .lcout(M_this_spr_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_0),
            .carryout(un1_M_this_spr_address_q_cry_1),
            .clk(N__42012),
            .ce(),
            .sr(N__41653));
    defparam M_this_spr_address_q_2_LC_22_14_2.C_ON=1'b1;
    defparam M_this_spr_address_q_2_LC_22_14_2.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_2_LC_22_14_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_2_LC_22_14_2 (
            .in0(N__33211),
            .in1(N__32211),
            .in2(_gnd_net_),
            .in3(N__32191),
            .lcout(M_this_spr_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_1),
            .carryout(un1_M_this_spr_address_q_cry_2),
            .clk(N__42012),
            .ce(),
            .sr(N__41653));
    defparam M_this_spr_address_q_3_LC_22_14_3.C_ON=1'b1;
    defparam M_this_spr_address_q_3_LC_22_14_3.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_3_LC_22_14_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_3_LC_22_14_3 (
            .in0(N__33215),
            .in1(N__31998),
            .in2(_gnd_net_),
            .in3(N__31975),
            .lcout(M_this_spr_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_2),
            .carryout(un1_M_this_spr_address_q_cry_3),
            .clk(N__42012),
            .ce(),
            .sr(N__41653));
    defparam M_this_spr_address_q_4_LC_22_14_4.C_ON=1'b1;
    defparam M_this_spr_address_q_4_LC_22_14_4.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_4_LC_22_14_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_4_LC_22_14_4 (
            .in0(N__33212),
            .in1(N__31779),
            .in2(_gnd_net_),
            .in3(N__31759),
            .lcout(M_this_spr_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_3),
            .carryout(un1_M_this_spr_address_q_cry_4),
            .clk(N__42012),
            .ce(),
            .sr(N__41653));
    defparam M_this_spr_address_q_5_LC_22_14_5.C_ON=1'b1;
    defparam M_this_spr_address_q_5_LC_22_14_5.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_5_LC_22_14_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_5_LC_22_14_5 (
            .in0(N__33216),
            .in1(N__31581),
            .in2(_gnd_net_),
            .in3(N__31549),
            .lcout(M_this_spr_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_4),
            .carryout(un1_M_this_spr_address_q_cry_5),
            .clk(N__42012),
            .ce(),
            .sr(N__41653));
    defparam M_this_spr_address_q_6_LC_22_14_6.C_ON=1'b1;
    defparam M_this_spr_address_q_6_LC_22_14_6.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_6_LC_22_14_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_6_LC_22_14_6 (
            .in0(N__33213),
            .in1(N__31371),
            .in2(_gnd_net_),
            .in3(N__31351),
            .lcout(M_this_spr_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_5),
            .carryout(un1_M_this_spr_address_q_cry_6),
            .clk(N__42012),
            .ce(),
            .sr(N__41653));
    defparam M_this_spr_address_q_7_LC_22_14_7.C_ON=1'b1;
    defparam M_this_spr_address_q_7_LC_22_14_7.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_7_LC_22_14_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_7_LC_22_14_7 (
            .in0(N__33217),
            .in1(N__31159),
            .in2(_gnd_net_),
            .in3(N__31141),
            .lcout(M_this_spr_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_6),
            .carryout(un1_M_this_spr_address_q_cry_7),
            .clk(N__42012),
            .ce(),
            .sr(N__41653));
    defparam M_this_spr_address_q_8_LC_22_15_0.C_ON=1'b1;
    defparam M_this_spr_address_q_8_LC_22_15_0.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_8_LC_22_15_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_8_LC_22_15_0 (
            .in0(N__33206),
            .in1(N__33700),
            .in2(_gnd_net_),
            .in3(N__33682),
            .lcout(M_this_spr_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_22_15_0_),
            .carryout(un1_M_this_spr_address_q_cry_8),
            .clk(N__42022),
            .ce(),
            .sr(N__41652));
    defparam M_this_spr_address_q_9_LC_22_15_1.C_ON=1'b1;
    defparam M_this_spr_address_q_9_LC_22_15_1.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_9_LC_22_15_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_9_LC_22_15_1 (
            .in0(N__33209),
            .in1(N__33482),
            .in2(_gnd_net_),
            .in3(N__33457),
            .lcout(M_this_spr_address_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_8),
            .carryout(un1_M_this_spr_address_q_cry_9),
            .clk(N__42022),
            .ce(),
            .sr(N__41652));
    defparam M_this_spr_address_q_10_LC_22_15_2.C_ON=1'b1;
    defparam M_this_spr_address_q_10_LC_22_15_2.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_10_LC_22_15_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_10_LC_22_15_2 (
            .in0(N__33204),
            .in1(N__33264),
            .in2(_gnd_net_),
            .in3(N__33226),
            .lcout(M_this_spr_address_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_9),
            .carryout(un1_M_this_spr_address_q_cry_10),
            .clk(N__42022),
            .ce(),
            .sr(N__41652));
    defparam M_this_spr_address_q_11_LC_22_15_3.C_ON=1'b1;
    defparam M_this_spr_address_q_11_LC_22_15_3.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_11_LC_22_15_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_11_LC_22_15_3 (
            .in0(N__33208),
            .in1(N__38846),
            .in2(_gnd_net_),
            .in3(N__33223),
            .lcout(M_this_spr_address_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_10),
            .carryout(un1_M_this_spr_address_q_cry_11),
            .clk(N__42022),
            .ce(),
            .sr(N__41652));
    defparam M_this_spr_address_q_12_LC_22_15_4.C_ON=1'b1;
    defparam M_this_spr_address_q_12_LC_22_15_4.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_12_LC_22_15_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_12_LC_22_15_4 (
            .in0(N__33205),
            .in1(N__38902),
            .in2(_gnd_net_),
            .in3(N__33220),
            .lcout(M_this_spr_address_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_11),
            .carryout(un1_M_this_spr_address_q_cry_12),
            .clk(N__42022),
            .ce(),
            .sr(N__41652));
    defparam M_this_spr_address_q_13_LC_22_15_5.C_ON=1'b0;
    defparam M_this_spr_address_q_13_LC_22_15_5.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_13_LC_22_15_5.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_spr_address_q_13_LC_22_15_5 (
            .in0(N__38755),
            .in1(N__33207),
            .in2(_gnd_net_),
            .in3(N__33118),
            .lcout(M_this_spr_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42022),
            .ce(),
            .sr(N__41652));
    defparam \this_spr_ram.mem_radreg_11_LC_22_16_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_11_LC_22_16_0 .SEQ_MODE=4'b1000;
    defparam \this_spr_ram.mem_radreg_11_LC_22_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_spr_ram.mem_radreg_11_LC_22_16_0  (
            .in0(N__33115),
            .in1(N__43935),
            .in2(_gnd_net_),
            .in3(N__38205),
            .lcout(\this_spr_ram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42028),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_12_LC_22_16_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_12_LC_22_16_4 .SEQ_MODE=4'b1000;
    defparam \this_spr_ram.mem_radreg_12_LC_22_16_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_spr_ram.mem_radreg_12_LC_22_16_4  (
            .in0(N__34027),
            .in1(N__41602),
            .in2(_gnd_net_),
            .in3(N__38206),
            .lcout(\this_spr_ram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42028),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_6_LC_22_17_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_6_LC_22_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_6_LC_22_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_6_LC_22_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33109),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42038),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_22_17_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_22_17_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_22_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_22_17_2  (
            .in0(N__39107),
            .in1(N__34021),
            .in2(_gnd_net_),
            .in3(N__34006),
            .lcout(),
            .ltout(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_22_17_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_22_17_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_22_17_3 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_22_17_3  (
            .in0(N__37027),
            .in1(N__36978),
            .in2(N__33988),
            .in3(N__36628),
            .lcout(),
            .ltout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_22_17_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_22_17_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_22_17_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_22_17_4  (
            .in0(N__36979),
            .in1(N__37861),
            .in2(N__33985),
            .in3(N__36754),
            .lcout(M_this_spr_ram_read_data_2),
            .ltout(M_this_spr_ram_read_data_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNITTE65_5_LC_22_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNITTE65_5_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNITTE65_5_LC_22_17_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNITTE65_5_LC_22_17_5  (
            .in0(N__34476),
            .in1(N__37122),
            .in2(N__33982),
            .in3(N__34437),
            .lcout(M_this_ppu_vram_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_22_17_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_22_17_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_22_17_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_22_17_6  (
            .in0(N__39106),
            .in1(N__33964),
            .in2(_gnd_net_),
            .in3(N__33949),
            .lcout(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_22_18_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_22_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_22_18_0  (
            .in0(N__39121),
            .in1(N__33931),
            .in2(_gnd_net_),
            .in3(N__33919),
            .lcout(),
            .ltout(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_22_18_1 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_22_18_1 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_22_18_1 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_22_18_1  (
            .in0(N__39019),
            .in1(N__36995),
            .in2(N__33898),
            .in3(N__37038),
            .lcout(),
            .ltout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_22_18_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_22_18_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_22_18_2  (
            .in0(N__36999),
            .in1(N__36790),
            .in2(N__33895),
            .in3(N__36013),
            .lcout(M_this_spr_ram_read_data_1),
            .ltout(M_this_spr_ram_read_data_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.vram_en_iv_i_0_o2_LC_22_18_3 .C_ON=1'b0;
    defparam \this_ppu.vram_en_iv_i_0_o2_LC_22_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.vram_en_iv_i_0_o2_LC_22_18_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.vram_en_iv_i_0_o2_LC_22_18_3  (
            .in0(N__36945),
            .in1(N__34384),
            .in2(N__34378),
            .in3(N__34296),
            .lcout(\this_ppu.N_1000_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_RNIB2R65_4_LC_22_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_RNIB2R65_4_LC_22_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_RNIB2R65_4_LC_22_18_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_ppu.M_screen_y_q_RNIB2R65_4_LC_22_18_5  (
            .in0(N__34477),
            .in1(N__34430),
            .in2(N__37345),
            .in3(N__34336),
            .lcout(M_this_ppu_vram_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_22_18_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_22_18_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_22_18_6 .LUT_INIT=16'b1110001100100011;
    LogicCell40 \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_22_18_6  (
            .in0(N__36826),
            .in1(N__36712),
            .in2(N__37003),
            .in3(N__34312),
            .lcout(M_this_spr_ram_read_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_22_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_22_19_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_22_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_22_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34285),
            .lcout(this_vga_signals_M_vcounter_q_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42058),
            .ce(N__34251),
            .sr(N__34220));
    defparam \this_vga_signals.un5_vaddress_g0_3_2_LC_22_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_2_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_2_LC_22_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_2_LC_22_19_1  (
            .in0(_gnd_net_),
            .in1(N__34842),
            .in2(_gnd_net_),
            .in3(N__35306),
            .lcout(\this_vga_signals.N_5_i_0 ),
            .ltout(\this_vga_signals.N_5_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_22_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_22_19_2 .LUT_INIT=16'b0111100010000111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_12_LC_22_19_2  (
            .in0(N__34074),
            .in1(N__35610),
            .in2(N__34177),
            .in3(N__35710),
            .lcout(\this_vga_signals.mult1_un47_sum_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_21_1_LC_22_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_21_1_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_21_1_LC_22_19_3 .LUT_INIT=16'b0011011011111010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_21_1_LC_22_19_3  (
            .in0(N__35314),
            .in1(N__35611),
            .in2(N__34938),
            .in3(N__34073),
            .lcout(\this_vga_signals.g0_21_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_40_LC_22_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_40_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_40_LC_22_19_4 .LUT_INIT=16'b0010111000111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_40_LC_22_19_4  (
            .in0(N__35307),
            .in1(N__34153),
            .in2(N__34897),
            .in3(N__34124),
            .lcout(\this_vga_signals.if_N_7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_22_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_22_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_22_19_6 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_30_LC_22_19_6  (
            .in0(N__34075),
            .in1(N__35712),
            .in2(N__35617),
            .in3(N__35665),
            .lcout(\this_vga_signals.mult1_un47_sum_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_43_LC_22_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_43_LC_22_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_43_LC_22_19_7 .LUT_INIT=16'b1001011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_43_LC_22_19_7  (
            .in0(N__35711),
            .in1(N__35664),
            .in2(N__35629),
            .in3(N__35615),
            .lcout(\this_vga_signals.mult1_un47_sum_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_45_LC_22_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_45_LC_22_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_45_LC_22_20_2 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_45_LC_22_20_2  (
            .in0(N__35557),
            .in1(N__35527),
            .in2(N__35519),
            .in3(N__35392),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_d_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_6_LC_22_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_6_LC_22_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_6_LC_22_20_3 .LUT_INIT=16'b1100110010010011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_6_LC_22_20_3  (
            .in0(N__35303),
            .in1(N__35134),
            .in2(N__34942),
            .in3(N__34749),
            .lcout(\this_vga_signals.vaddress_0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNILD7F7_6_LC_22_21_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNILD7F7_6_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNILD7F7_6_LC_22_21_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNILD7F7_6_LC_22_21_1  (
            .in0(N__36560),
            .in1(N__39460),
            .in2(N__34624),
            .in3(N__37736),
            .lcout(\this_ppu.M_screen_y_q_esr_RNILD7F7Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_3_LC_22_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_3_LC_22_21_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_3_LC_22_21_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_1_0_i_3_LC_22_21_4  (
            .in0(N__35992),
            .in1(N__41510),
            .in2(N__39898),
            .in3(N__36484),
            .lcout(M_this_spr_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_1_x_0_LC_22_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_1_x_0_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_1_x_0_LC_22_21_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_0_a2_1_x_0_LC_22_21_5  (
            .in0(N__42649),
            .in1(N__35782),
            .in2(_gnd_net_),
            .in3(N__43222),
            .lcout(\this_ppu.M_this_state_q_srsts_0_0_a2_1_xZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIUUE65_6_LC_22_21_6 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIUUE65_6_LC_22_21_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIUUE65_6_LC_22_21_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIUUE65_6_LC_22_21_6  (
            .in0(N__34469),
            .in1(N__34438),
            .in2(N__36567),
            .in3(N__36949),
            .lcout(M_this_ppu_vram_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_en_0_i_0_0_0_LC_22_22_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_en_0_i_0_0_0_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_en_0_i_0_0_0_LC_22_22_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \this_ppu.M_this_spr_ram_write_en_0_i_0_0_0_LC_22_22_0  (
            .in0(N__36477),
            .in1(N__36437),
            .in2(_gnd_net_),
            .in3(N__43431),
            .lcout(M_this_spr_ram_write_en_0_i_1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_1_0_LC_22_22_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_1_0_LC_22_22_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_1_0_LC_22_22_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_0_a2_1_0_LC_22_22_1  (
            .in0(N__43799),
            .in1(N__42648),
            .in2(_gnd_net_),
            .in3(N__35719),
            .lcout(\this_ppu.N_1257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_1_LC_22_22_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_1_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_1_LC_22_22_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_1_0_i_1_LC_22_22_2  (
            .in0(N__36478),
            .in1(N__39783),
            .in2(N__40052),
            .in3(N__35988),
            .lcout(M_this_spr_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_14_LC_22_22_7.C_ON=1'b0;
    defparam M_this_state_q_14_LC_22_22_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_14_LC_22_22_7.LUT_INIT=16'b0000000010001000;
    LogicCell40 M_this_state_q_14_LC_22_22_7 (
            .in0(N__43432),
            .in1(N__36438),
            .in2(_gnd_net_),
            .in3(N__43241),
            .lcout(M_this_state_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42092),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a2_1_1_LC_22_23_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a2_1_1_LC_22_23_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a2_1_1_LC_22_23_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a2_1_1_LC_22_23_0  (
            .in0(_gnd_net_),
            .in1(N__36335),
            .in2(_gnd_net_),
            .in3(N__38595),
            .lcout(N_1258),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam led_1_7_5__m17_0_a3_0_a3_0_a2_LC_22_23_2.C_ON=1'b0;
    defparam led_1_7_5__m17_0_a3_0_a3_0_a2_LC_22_23_2.SEQ_MODE=4'b0000;
    defparam led_1_7_5__m17_0_a3_0_a3_0_a2_LC_22_23_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 led_1_7_5__m17_0_a3_0_a3_0_a2_LC_22_23_2 (
            .in0(_gnd_net_),
            .in1(N__35830),
            .in2(_gnd_net_),
            .in3(N__37785),
            .lcout(N_1416),
            .ltout(N_1416_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam led_1_7_5__m17_0_a3_0_a3_0_a3_2_LC_22_23_3.C_ON=1'b0;
    defparam led_1_7_5__m17_0_a3_0_a3_0_a3_2_LC_22_23_3.SEQ_MODE=4'b0000;
    defparam led_1_7_5__m17_0_a3_0_a3_0_a3_2_LC_22_23_3.LUT_INIT=16'b0000000011000000;
    LogicCell40 led_1_7_5__m17_0_a3_0_a3_0_a3_2_LC_22_23_3 (
            .in0(_gnd_net_),
            .in1(N__42240),
            .in2(N__35800),
            .in3(N__38287),
            .lcout(N_1151_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_4_LC_22_23_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_4_LC_22_23_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_4_LC_22_23_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a3_1_4_LC_22_23_4  (
            .in0(N__43489),
            .in1(N__40747),
            .in2(_gnd_net_),
            .in3(N__38597),
            .lcout(N_1066),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_1_sx_0_LC_22_23_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_1_sx_0_LC_22_23_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_0_a2_1_sx_0_LC_22_23_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_0_a2_1_sx_0_LC_22_23_5  (
            .in0(N__43855),
            .in1(N__35781),
            .in2(N__43894),
            .in3(N__43220),
            .lcout(\this_ppu.M_this_state_q_srsts_0_0_a2_1_sxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a2_0_5_LC_22_23_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a2_0_5_LC_22_23_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a2_0_5_LC_22_23_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a2_0_5_LC_22_23_6  (
            .in0(N__43488),
            .in1(N__36336),
            .in2(_gnd_net_),
            .in3(N__38596),
            .lcout(N_1276),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_en_0_i_0_0_i_0_LC_22_23_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_en_0_i_0_0_i_0_LC_22_23_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_en_0_i_0_0_i_0_LC_22_23_7 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \this_ppu.M_this_spr_ram_write_en_0_i_0_0_i_0_LC_22_23_7  (
            .in0(N__36476),
            .in1(N__36445),
            .in2(_gnd_net_),
            .in3(N__43487),
            .lcout(M_this_spr_ram_write_en_0_i_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_q_0_i_0_o2_5_LC_22_24_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_o2_5_LC_22_24_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_o2_5_LC_22_24_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_o2_5_LC_22_24_3  (
            .in0(N__36350),
            .in1(N__43502),
            .in2(_gnd_net_),
            .in3(N__38605),
            .lcout(N_801_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1_LC_22_24_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1_LC_22_24_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1_LC_22_24_4 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \this_ppu.M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1_LC_22_24_4  (
            .in0(N__42614),
            .in1(N__36272),
            .in2(N__36235),
            .in3(N__36152),
            .lcout(this_ppu_M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_1_1_LC_22_25_2.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_1_1_LC_22_25_2.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_1_1_LC_22_25_2.LUT_INIT=16'b0011001100100010;
    LogicCell40 M_this_map_address_q_RNO_1_1_LC_22_25_2 (
            .in0(N__39381),
            .in1(N__42499),
            .in2(_gnd_net_),
            .in3(N__38534),
            .lcout(),
            .ltout(M_this_map_address_qc_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_0_1_LC_22_25_3.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_0_1_LC_22_25_3.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_0_1_LC_22_25_3.LUT_INIT=16'b1011000011110000;
    LogicCell40 M_this_map_address_q_RNO_0_1_LC_22_25_3 (
            .in0(N__39781),
            .in1(N__43503),
            .in2(N__36118),
            .in3(N__38606),
            .lcout(M_this_map_address_qc_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a2_1_LC_22_26_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a2_1_LC_22_26_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a2_1_LC_22_26_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a2_1_LC_22_26_3  (
            .in0(N__42262),
            .in1(N__43501),
            .in2(_gnd_net_),
            .in3(N__36115),
            .lcout(N_1242),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_i_0_0_LC_22_29_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_0_LC_22_29_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_0_LC_22_29_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_i_0_0_LC_22_29_3  (
            .in0(_gnd_net_),
            .in1(N__42443),
            .in2(_gnd_net_),
            .in3(N__40122),
            .lcout(N_169_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam led_1_7_5__N_1048_i_LC_23_8_4.C_ON=1'b0;
    defparam led_1_7_5__N_1048_i_LC_23_8_4.SEQ_MODE=4'b0000;
    defparam led_1_7_5__N_1048_i_LC_23_8_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 led_1_7_5__N_1048_i_LC_23_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38482),
            .lcout(N_1048_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_23_15_1 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_23_15_1 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_23_15_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_23_15_1  (
            .in0(N__36043),
            .in1(N__36028),
            .in2(_gnd_net_),
            .in3(N__39117),
            .lcout(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_23_16_7 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_23_16_7 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_23_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_23_16_7  (
            .in0(N__36784),
            .in1(N__36769),
            .in2(_gnd_net_),
            .in3(N__39105),
            .lcout(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_23_17_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_23_17_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_23_17_0  (
            .in0(N__39100),
            .in1(N__36748),
            .in2(_gnd_net_),
            .in3(N__36730),
            .lcout(),
            .ltout(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_23_17_1 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_23_17_1 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_23_17_1 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_23_17_1  (
            .in0(N__37037),
            .in1(N__37002),
            .in2(N__36715),
            .in3(N__39139),
            .lcout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_7_0_wclke_3_LC_23_17_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_7_0_wclke_3_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_7_0_wclke_3_LC_23_17_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_spr_ram.mem_mem_7_0_wclke_3_LC_23_17_3  (
            .in0(N__38923),
            .in1(N__38847),
            .in2(N__38795),
            .in3(N__38709),
            .lcout(\this_spr_ram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_13_LC_23_17_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_13_LC_23_17_4 .SEQ_MODE=4'b1000;
    defparam \this_spr_ram.mem_radreg_13_LC_23_17_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_spr_ram.mem_radreg_13_LC_23_17_4  (
            .in0(N__36676),
            .in1(N__39006),
            .in2(_gnd_net_),
            .in3(N__38204),
            .lcout(\this_spr_ram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42046),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_23_17_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_23_17_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_23_17_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_23_17_6  (
            .in0(N__39099),
            .in1(N__36661),
            .in2(_gnd_net_),
            .in3(N__36640),
            .lcout(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_23_17_7 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_23_17_7 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_23_17_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_23_17_7  (
            .in0(N__39098),
            .in1(N__36622),
            .in2(_gnd_net_),
            .in3(N__36610),
            .lcout(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_6_LC_23_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_6_LC_23_18_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_6_LC_23_18_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_6_LC_23_18_1  (
            .in0(N__37344),
            .in1(N__37290),
            .in2(N__37134),
            .in3(N__36595),
            .lcout(\this_ppu.M_screen_y_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42059),
            .ce(N__37177),
            .sr(N__43098));
    defparam \this_ppu.M_screen_y_q_esr_5_LC_23_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_5_LC_23_18_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_5_LC_23_18_2 .LUT_INIT=16'b0111100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_5_LC_23_18_2  (
            .in0(N__37343),
            .in1(N__37291),
            .in2(N__37133),
            .in3(N__37264),
            .lcout(\this_ppu.M_screen_y_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42059),
            .ce(N__37177),
            .sr(N__43098));
    defparam \this_ppu.M_screen_y_q_esr_RNIJB7F7_5_LC_23_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIJB7F7_5_LC_23_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIJB7F7_5_LC_23_18_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIJB7F7_5_LC_23_18_4  (
            .in0(N__37123),
            .in1(N__39492),
            .in2(N__37093),
            .in3(N__37734),
            .lcout(\this_ppu.M_screen_y_q_esr_RNIJB7F7Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNITCNI1_12_LC_23_18_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_12_LC_23_18_5 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_12_LC_23_18_5 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_spr_ram.mem_radreg_RNITCNI1_12_LC_23_18_5  (
            .in0(N__37000),
            .in1(N__36865),
            .in2(N__37042),
            .in3(N__37009),
            .lcout(),
            .ltout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNINL8S2_11_LC_23_18_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_11_LC_23_18_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_11_LC_23_18_6 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \this_spr_ram.mem_radreg_RNINL8S2_11_LC_23_18_6  (
            .in0(N__36901),
            .in1(N__37001),
            .in2(N__36952),
            .in3(N__37819),
            .lcout(M_this_spr_ram_read_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_23_19_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_23_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_23_19_2  (
            .in0(N__36934),
            .in1(N__36919),
            .in2(_gnd_net_),
            .in3(N__39110),
            .lcout(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_23_19_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_23_19_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_23_19_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_23_19_3  (
            .in0(N__39109),
            .in1(N__36895),
            .in2(_gnd_net_),
            .in3(N__36880),
            .lcout(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_23_19_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_23_19_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_23_19_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_23_19_4  (
            .in0(N__36859),
            .in1(N__36838),
            .in2(_gnd_net_),
            .in3(N__39112),
            .lcout(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_23_19_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_23_19_5 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_23_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_23_19_5  (
            .in0(N__39113),
            .in1(N__36820),
            .in2(_gnd_net_),
            .in3(N__36802),
            .lcout(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_LC_23_19_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_LC_23_19_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_LC_23_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_3_1_RNISI5G_LC_23_19_6  (
            .in0(N__37891),
            .in1(N__37873),
            .in2(_gnd_net_),
            .in3(N__39108),
            .lcout(\this_spr_ram.mem_mem_3_1_RNISI5GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_23_19_7 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_23_19_7 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_23_19_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_23_19_7  (
            .in0(N__39111),
            .in1(_gnd_net_),
            .in2(N__37849),
            .in3(N__37831),
            .lcout(\this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_ext_address_q_9_LC_23_20_0.C_ON=1'b0;
    defparam M_this_ext_address_q_9_LC_23_20_0.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_9_LC_23_20_0.LUT_INIT=16'b1010111010100010;
    LogicCell40 M_this_ext_address_q_9_LC_23_20_0 (
            .in0(N__40606),
            .in1(N__43543),
            .in2(N__41153),
            .in3(N__39784),
            .lcout(M_this_ext_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42082),
            .ce(),
            .sr(N__43100));
    defparam M_this_ctrl_flags_q_7_LC_23_21_2.C_ON=1'b0;
    defparam M_this_ctrl_flags_q_7_LC_23_21_2.SEQ_MODE=4'b1000;
    defparam M_this_ctrl_flags_q_7_LC_23_21_2.LUT_INIT=16'b1110001010101010;
    LogicCell40 M_this_ctrl_flags_q_7_LC_23_21_2 (
            .in0(N__37800),
            .in1(N__40880),
            .in2(N__39897),
            .in3(N__43544),
            .lcout(M_this_ctrl_flags_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42093),
            .ce(),
            .sr(N__43103));
    defparam led_1_7_5__m5_i_a2_i_o3_i_a3_LC_23_22_3.C_ON=1'b0;
    defparam led_1_7_5__m5_i_a2_i_o3_i_a3_LC_23_22_3.SEQ_MODE=4'b0000;
    defparam led_1_7_5__m5_i_a2_i_o3_i_a3_LC_23_22_3.LUT_INIT=16'b0000000001010101;
    LogicCell40 led_1_7_5__m5_i_a2_i_o3_i_a3_LC_23_22_3 (
            .in0(N__37399),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37789),
            .lcout(m5_i_a2_i_o3_i_a3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam N_38_i_0_sbtinv_LC_23_22_7.C_ON=1'b0;
    defparam N_38_i_0_sbtinv_LC_23_22_7.SEQ_MODE=4'b0000;
    defparam N_38_i_0_sbtinv_LC_23_22_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 N_38_i_0_sbtinv_LC_23_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37748),
            .lcout(N_38_i_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_this_state_q_7_i_0_0_0_LC_23_23_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_state_q_7_i_0_0_0_LC_23_23_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_state_q_7_i_0_0_0_LC_23_23_0 .LUT_INIT=16'b1100111001001110;
    LogicCell40 \this_ppu.un1_M_this_state_q_7_i_0_0_0_LC_23_23_0  (
            .in0(N__37459),
            .in1(N__43485),
            .in2(N__42261),
            .in3(N__38285),
            .lcout(this_ppu_un1_M_this_state_q_7_i_0_0_0),
            .ltout(this_ppu_un1_M_this_state_q_7_i_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_0_c_RNO_LC_23_23_1.C_ON=1'b0;
    defparam un1_M_this_map_address_q_cry_0_c_RNO_LC_23_23_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_0_c_RNO_LC_23_23_1.LUT_INIT=16'b0000000011110000;
    LogicCell40 un1_M_this_map_address_q_cry_0_c_RNO_LC_23_23_1 (
            .in0(_gnd_net_),
            .in1(N__39563),
            .in2(N__37441),
            .in3(N__39198),
            .lcout(un1_M_this_map_address_q_cry_0_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam led_1_7_5__m12_0_a3_0_a3_0_a3_LC_23_23_2.C_ON=1'b0;
    defparam led_1_7_5__m12_0_a3_0_a3_0_a3_LC_23_23_2.SEQ_MODE=4'b0000;
    defparam led_1_7_5__m12_0_a3_0_a3_0_a3_LC_23_23_2.LUT_INIT=16'b0000000010000000;
    LogicCell40 led_1_7_5__m12_0_a3_0_a3_0_a3_LC_23_23_2 (
            .in0(N__37437),
            .in1(N__37405),
            .in2(N__41130),
            .in3(N__37395),
            .lcout(led_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_2_LC_23_23_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_2_LC_23_23_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_2_LC_23_23_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a3_1_2_LC_23_23_3  (
            .in0(N__43486),
            .in1(N__42774),
            .in2(_gnd_net_),
            .in3(N__38598),
            .lcout(N_1058),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_this_state_q_7_i_0_a3_0_0_LC_23_23_4 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_state_q_7_i_0_a3_0_0_LC_23_23_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_state_q_7_i_0_a3_0_0_LC_23_23_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.un1_M_this_state_q_7_i_0_a3_0_0_LC_23_23_4  (
            .in0(N__40840),
            .in1(N__43484),
            .in2(_gnd_net_),
            .in3(N__38286),
            .lcout(un1_M_this_state_q_7_i_0_a3_0_0),
            .ltout(un1_M_this_state_q_7_i_0_a3_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_1_0_LC_23_23_5.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_1_0_LC_23_23_5.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_1_0_LC_23_23_5.LUT_INIT=16'b1111010100001010;
    LogicCell40 M_this_map_address_q_RNO_1_0_LC_23_23_5 (
            .in0(N__38260),
            .in1(_gnd_net_),
            .in2(N__38254),
            .in3(N__39562),
            .lcout(un1_M_this_map_address_q_axb_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_23_23_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_23_23_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_23_23_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_23_23_6  (
            .in0(N__38251),
            .in1(N__38226),
            .in2(_gnd_net_),
            .in3(N__38198),
            .lcout(read_data_RNI4PFJ1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_2_LC_23_24_0.C_ON=1'b0;
    defparam M_this_map_address_q_2_LC_23_24_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_2_LC_23_24_0.LUT_INIT=16'b0000100000001010;
    LogicCell40 M_this_map_address_q_2_LC_23_24_0 (
            .in0(N__38503),
            .in1(N__39298),
            .in2(N__37912),
            .in3(N__42259),
            .lcout(M_this_map_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42115),
            .ce(),
            .sr(N__41643));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_3_LC_23_24_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_3_LC_23_24_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_3_LC_23_24_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a3_1_3_LC_23_24_3  (
            .in0(N__41509),
            .in1(N__43499),
            .in2(_gnd_net_),
            .in3(N__38608),
            .lcout(),
            .ltout(N_1062_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_3_LC_23_24_4.C_ON=1'b0;
    defparam M_this_map_address_q_3_LC_23_24_4.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_3_LC_23_24_4.LUT_INIT=16'b0000100000001010;
    LogicCell40 M_this_map_address_q_3_LC_23_24_4 (
            .in0(N__37897),
            .in1(N__39253),
            .in2(N__37900),
            .in3(N__42260),
            .lcout(M_this_map_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42115),
            .ce(),
            .sr(N__41643));
    defparam M_this_map_address_q_RNO_0_3_LC_23_24_5.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_0_3_LC_23_24_5.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_0_3_LC_23_24_5.LUT_INIT=16'b0011001100100010;
    LogicCell40 M_this_map_address_q_RNO_0_3_LC_23_24_5 (
            .in0(N__39273),
            .in1(N__42529),
            .in2(_gnd_net_),
            .in3(N__38532),
            .lcout(M_this_map_address_qc_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_0_4_LC_23_24_6.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_0_4_LC_23_24_6.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_0_4_LC_23_24_6.LUT_INIT=16'b0000111100001010;
    LogicCell40 M_this_map_address_q_RNO_0_4_LC_23_24_6 (
            .in0(N__38533),
            .in1(_gnd_net_),
            .in2(N__42542),
            .in3(N__39228),
            .lcout(),
            .ltout(M_this_map_address_qc_6_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_4_LC_23_24_7.C_ON=1'b0;
    defparam M_this_map_address_q_4_LC_23_24_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_4_LC_23_24_7.LUT_INIT=16'b0011000000010000;
    LogicCell40 M_this_map_address_q_4_LC_23_24_7 (
            .in0(N__42258),
            .in1(N__38617),
            .in2(N__38611),
            .in3(N__39208),
            .lcout(M_this_map_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42115),
            .ce(),
            .sr(N__41643));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_0_LC_23_25_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_0_LC_23_25_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_1_0_LC_23_25_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a3_1_0_LC_23_25_0  (
            .in0(N__42445),
            .in1(N__43500),
            .in2(_gnd_net_),
            .in3(N__38607),
            .lcout(N_1097),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_0_0_LC_23_25_3.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_0_0_LC_23_25_3.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_0_0_LC_23_25_3.LUT_INIT=16'b0011001100100010;
    LogicCell40 M_this_map_address_q_RNO_0_0_LC_23_25_3 (
            .in0(N__39547),
            .in1(N__42507),
            .in2(_gnd_net_),
            .in3(N__38535),
            .lcout(M_this_map_address_qc_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_0_2_LC_23_25_6.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_0_2_LC_23_25_6.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_0_2_LC_23_25_6.LUT_INIT=16'b0000000011101110;
    LogicCell40 M_this_map_address_q_RNO_0_2_LC_23_25_6 (
            .in0(N__38536),
            .in1(N__39318),
            .in2(_gnd_net_),
            .in3(N__42508),
            .lcout(M_this_map_address_qc_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_i_0_1_LC_23_29_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_1_LC_23_29_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_1_LC_23_29_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_i_0_1_LC_23_29_1  (
            .in0(_gnd_net_),
            .in1(N__39761),
            .in2(_gnd_net_),
            .in3(N__40150),
            .lcout(N_918_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam N_1048_sbtinv_LC_23_30_0.C_ON=1'b0;
    defparam N_1048_sbtinv_LC_23_30_0.SEQ_MODE=4'b0000;
    defparam N_1048_sbtinv_LC_23_30_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 N_1048_sbtinv_LC_23_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38478),
            .lcout(N_1048_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_0_wclke_3_LC_24_14_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_0_wclke_3_LC_24_14_0 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_0_wclke_3_LC_24_14_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_spr_ram.mem_mem_1_0_wclke_3_LC_24_14_0  (
            .in0(N__38921),
            .in1(N__38859),
            .in2(N__38793),
            .in3(N__38719),
            .lcout(\this_spr_ram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_0_wclke_3_LC_24_15_1 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_0_wclke_3_LC_24_15_1 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_0_wclke_3_LC_24_15_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_spr_ram.mem_mem_3_0_wclke_3_LC_24_15_1  (
            .in0(N__38717),
            .in1(N__38904),
            .in2(N__38858),
            .in3(N__38759),
            .lcout(\this_spr_ram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_0_wclke_3_LC_24_15_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_0_wclke_3_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_0_wclke_3_LC_24_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_spr_ram.mem_mem_0_0_wclke_3_LC_24_15_2  (
            .in0(N__38903),
            .in1(N__38839),
            .in2(N__38776),
            .in3(N__38716),
            .lcout(\this_spr_ram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_0_wclke_3_LC_24_16_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_0_wclke_3_LC_24_16_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_0_wclke_3_LC_24_16_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_spr_ram.mem_mem_2_0_wclke_3_LC_24_16_4  (
            .in0(N__38922),
            .in1(N__38865),
            .in2(N__38794),
            .in3(N__38718),
            .lcout(\this_spr_ram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_24_17_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_24_17_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_24_17_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_24_17_6  (
            .in0(N__39163),
            .in1(N__39097),
            .in2(_gnd_net_),
            .in3(N__39154),
            .lcout(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_24_18_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_24_18_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_24_18_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_24_18_2  (
            .in0(N__39133),
            .in1(N__39104),
            .in2(_gnd_net_),
            .in3(N__39034),
            .lcout(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.IO_port_data_write_i_m2_i_m2_7_LC_24_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.IO_port_data_write_i_m2_i_m2_7_LC_24_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.IO_port_data_write_i_m2_i_m2_7_LC_24_19_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vga_signals.IO_port_data_write_i_m2_i_m2_7_LC_24_19_4  (
            .in0(N__39415),
            .in1(N__43681),
            .in2(_gnd_net_),
            .in3(N__39010),
            .lcout(IO_port_data_write_i_m2_i_m2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_4_0_wclke_3_LC_24_19_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_4_0_wclke_3_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_4_0_wclke_3_LC_24_19_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_spr_ram.mem_mem_4_0_wclke_3_LC_24_19_5  (
            .in0(N__38924),
            .in1(N__38861),
            .in2(N__38796),
            .in3(N__38701),
            .lcout(\this_spr_ram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_5_0_wclke_3_LC_24_19_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_5_0_wclke_3_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_5_0_wclke_3_LC_24_19_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_spr_ram.mem_mem_5_0_wclke_3_LC_24_19_6  (
            .in0(N__38702),
            .in1(N__38789),
            .in2(N__38866),
            .in3(N__38925),
            .lcout(\this_spr_ram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_6_0_wclke_3_LC_24_19_7 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_6_0_wclke_3_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_6_0_wclke_3_LC_24_19_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_spr_ram.mem_mem_6_0_wclke_3_LC_24_19_7  (
            .in0(N__38926),
            .in1(N__38860),
            .in2(N__38797),
            .in3(N__38703),
            .lcout(\this_spr_ram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_ext_address_q_0_LC_24_21_0.C_ON=1'b0;
    defparam M_this_ext_address_q_0_LC_24_21_0.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_0_LC_24_21_0.LUT_INIT=16'b0101101000010010;
    LogicCell40 M_this_ext_address_q_0_LC_24_21_0 (
            .in0(N__40312),
            .in1(N__43528),
            .in2(N__40281),
            .in3(N__41145),
            .lcout(M_this_ext_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42101),
            .ce(),
            .sr(N__43101));
    defparam M_this_status_flags_q_7_LC_24_21_1.C_ON=1'b0;
    defparam M_this_status_flags_q_7_LC_24_21_1.SEQ_MODE=4'b1000;
    defparam M_this_status_flags_q_7_LC_24_21_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 M_this_status_flags_q_7_LC_24_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39461),
            .lcout(M_this_status_flags_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42101),
            .ce(),
            .sr(N__43101));
    defparam M_this_map_address_q_1_LC_24_22_7.C_ON=1'b0;
    defparam M_this_map_address_q_1_LC_24_22_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_1_LC_24_22_7.LUT_INIT=16'b0100110011000100;
    LogicCell40 M_this_map_address_q_1_LC_24_22_7 (
            .in0(N__42288),
            .in1(N__39406),
            .in2(N__39377),
            .in3(N__39340),
            .lcout(M_this_map_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42109),
            .ce(),
            .sr(N__41647));
    defparam un1_M_this_map_address_q_cry_0_c_LC_24_23_0.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_0_c_LC_24_23_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_0_c_LC_24_23_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_map_address_q_cry_0_c_LC_24_23_0 (
            .in0(_gnd_net_),
            .in1(N__39394),
            .in2(N__39564),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_24_23_0_),
            .carryout(un1_M_this_map_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_0_THRU_LUT4_0_LC_24_23_1.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_0_THRU_LUT4_0_LC_24_23_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_0_THRU_LUT4_0_LC_24_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_map_address_q_cry_0_THRU_LUT4_0_LC_24_23_1 (
            .in0(_gnd_net_),
            .in1(N__39364),
            .in2(_gnd_net_),
            .in3(N__39334),
            .lcout(un1_M_this_map_address_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_0),
            .carryout(un1_M_this_map_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_1_2_LC_24_23_2.C_ON=1'b1;
    defparam M_this_map_address_q_RNO_1_2_LC_24_23_2.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_1_2_LC_24_23_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_RNO_1_2_LC_24_23_2 (
            .in0(_gnd_net_),
            .in1(N__39317),
            .in2(_gnd_net_),
            .in3(N__39292),
            .lcout(M_this_map_address_q_RNO_1Z0Z_2),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_1),
            .carryout(un1_M_this_map_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_1_3_LC_24_23_3.C_ON=1'b1;
    defparam M_this_map_address_q_RNO_1_3_LC_24_23_3.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_1_3_LC_24_23_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_RNO_1_3_LC_24_23_3 (
            .in0(_gnd_net_),
            .in1(N__39272),
            .in2(_gnd_net_),
            .in3(N__39247),
            .lcout(M_this_map_address_q_RNO_1Z0Z_3),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_2),
            .carryout(un1_M_this_map_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_1_4_LC_24_23_4.C_ON=1'b1;
    defparam M_this_map_address_q_RNO_1_4_LC_24_23_4.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_1_4_LC_24_23_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_RNO_1_4_LC_24_23_4 (
            .in0(_gnd_net_),
            .in1(N__39227),
            .in2(_gnd_net_),
            .in3(N__39202),
            .lcout(M_this_map_address_q_RNO_1Z0Z_4),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_3),
            .carryout(un1_M_this_map_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_1_5_LC_24_23_5.C_ON=1'b1;
    defparam M_this_map_address_q_RNO_1_5_LC_24_23_5.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_1_5_LC_24_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_map_address_q_RNO_1_5_LC_24_23_5 (
            .in0(_gnd_net_),
            .in1(N__39199),
            .in2(N__42183),
            .in3(N__39187),
            .lcout(M_this_map_address_q_RNO_1Z0Z_5),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_4),
            .carryout(un1_M_this_map_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_5_THRU_LUT4_0_LC_24_23_6.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_5_THRU_LUT4_0_LC_24_23_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_5_THRU_LUT4_0_LC_24_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_map_address_q_cry_5_THRU_LUT4_0_LC_24_23_6 (
            .in0(_gnd_net_),
            .in1(N__39632),
            .in2(_gnd_net_),
            .in3(N__39805),
            .lcout(un1_M_this_map_address_q_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_5),
            .carryout(un1_M_this_map_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_6_THRU_LUT4_0_LC_24_23_7.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_6_THRU_LUT4_0_LC_24_23_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_6_THRU_LUT4_0_LC_24_23_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_map_address_q_cry_6_THRU_LUT4_0_LC_24_23_7 (
            .in0(_gnd_net_),
            .in1(N__42869),
            .in2(_gnd_net_),
            .in3(N__39802),
            .lcout(un1_M_this_map_address_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_6),
            .carryout(un1_M_this_map_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_map_address_q_cry_7_THRU_LUT4_0_LC_24_24_0.C_ON=1'b1;
    defparam un1_M_this_map_address_q_cry_7_THRU_LUT4_0_LC_24_24_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_map_address_q_cry_7_THRU_LUT4_0_LC_24_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_map_address_q_cry_7_THRU_LUT4_0_LC_24_24_0 (
            .in0(_gnd_net_),
            .in1(N__41542),
            .in2(_gnd_net_),
            .in3(N__39799),
            .lcout(un1_M_this_map_address_q_cry_7_THRU_CO),
            .ltout(),
            .carryin(bfn_24_24_0_),
            .carryout(un1_M_this_map_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_9_LC_24_24_1.C_ON=1'b0;
    defparam M_this_map_address_q_9_LC_24_24_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_9_LC_24_24_1.LUT_INIT=16'b0100110010001100;
    LogicCell40 M_this_map_address_q_9_LC_24_24_1 (
            .in0(N__40808),
            .in1(N__40651),
            .in2(N__42295),
            .in3(N__39796),
            .lcout(M_this_map_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42120),
            .ce(),
            .sr(N__41645));
    defparam M_this_map_address_q_RNO_0_6_LC_24_25_0.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_0_6_LC_24_25_0.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_0_6_LC_24_25_0.LUT_INIT=16'b1100010100001101;
    LogicCell40 M_this_map_address_q_RNO_0_6_LC_24_25_0 (
            .in0(N__42834),
            .in1(N__42283),
            .in2(N__39633),
            .in3(N__39793),
            .lcout(),
            .ltout(M_this_map_address_qc_8_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_6_LC_24_25_1.C_ON=1'b0;
    defparam M_this_map_address_q_6_LC_24_25_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_6_LC_24_25_1.LUT_INIT=16'b0000000000001011;
    LogicCell40 M_this_map_address_q_6_LC_24_25_1 (
            .in0(N__39777),
            .in1(N__42588),
            .in2(N__39649),
            .in3(N__42541),
            .lcout(M_this_map_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42124),
            .ce(),
            .sr(N__41644));
    defparam M_this_map_address_q_8_LC_24_25_5.C_ON=1'b0;
    defparam M_this_map_address_q_8_LC_24_25_5.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_8_LC_24_25_5.LUT_INIT=16'b0111110100000000;
    LogicCell40 M_this_map_address_q_8_LC_24_25_5 (
            .in0(N__42284),
            .in1(N__39604),
            .in2(N__41550),
            .in3(N__41383),
            .lcout(M_this_map_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42124),
            .ce(),
            .sr(N__41644));
    defparam M_this_map_address_q_0_LC_24_26_2.C_ON=1'b0;
    defparam M_this_map_address_q_0_LC_24_26_2.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_0_LC_24_26_2.LUT_INIT=16'b0000100000001100;
    LogicCell40 M_this_map_address_q_0_LC_24_26_2 (
            .in0(N__39598),
            .in1(N__39589),
            .in2(N__39583),
            .in3(N__42289),
            .lcout(M_this_map_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42129),
            .ce(),
            .sr(N__41642));
    defparam \this_ppu.M_this_map_ram_write_data_i_0_4_LC_24_27_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_4_LC_24_27_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_4_LC_24_27_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_i_0_4_LC_24_27_6  (
            .in0(N__40685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40129),
            .lcout(N_921_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_i_0_2_LC_24_28_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_2_LC_24_28_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_2_LC_24_28_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_i_0_2_LC_24_28_6  (
            .in0(N__42750),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40151),
            .lcout(N_919_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_i_0_6_LC_24_29_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_6_LC_24_29_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_6_LC_24_29_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_i_0_6_LC_24_29_0  (
            .in0(N__40153),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40397),
            .lcout(N_923_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_i_0_3_LC_24_29_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_3_LC_24_29_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_3_LC_24_29_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_i_0_3_LC_24_29_5  (
            .in0(N__41466),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40152),
            .lcout(N_920_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_i_0_5_LC_24_30_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_5_LC_24_30_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_5_LC_24_30_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_i_0_5_LC_24_30_5  (
            .in0(_gnd_net_),
            .in1(N__40154),
            .in2(_gnd_net_),
            .in3(N__40061),
            .lcout(N_922_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_i_0_7_LC_24_30_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_7_LC_24_30_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_i_0_7_LC_24_30_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_i_0_7_LC_24_30_7  (
            .in0(_gnd_net_),
            .in1(N__40155),
            .in2(_gnd_net_),
            .in3(N__39905),
            .lcout(N_924_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_ext_address_q_13_LC_26_18_0.C_ON=1'b0;
    defparam M_this_ext_address_q_13_LC_26_18_0.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_13_LC_26_18_0.LUT_INIT=16'b1010111010100010;
    LogicCell40 M_this_ext_address_q_13_LC_26_18_0 (
            .in0(N__40555),
            .in1(N__43566),
            .in2(N__41160),
            .in3(N__40012),
            .lcout(M_this_ext_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42096),
            .ce(),
            .sr(N__43097));
    defparam M_this_ctrl_flags_q_5_LC_26_18_1.C_ON=1'b0;
    defparam M_this_ctrl_flags_q_5_LC_26_18_1.SEQ_MODE=4'b1000;
    defparam M_this_ctrl_flags_q_5_LC_26_18_1.LUT_INIT=16'b1110010011001100;
    LogicCell40 M_this_ctrl_flags_q_5_LC_26_18_1 (
            .in0(N__43564),
            .in1(N__39945),
            .in2(N__40032),
            .in3(N__40890),
            .lcout(M_this_ctrl_flags_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42096),
            .ce(),
            .sr(N__43097));
    defparam M_this_ext_address_q_2_LC_26_18_2.C_ON=1'b0;
    defparam M_this_ext_address_q_2_LC_26_18_2.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_2_LC_26_18_2.LUT_INIT=16'b0101101000010010;
    LogicCell40 M_this_ext_address_q_2_LC_26_18_2 (
            .in0(N__40210),
            .in1(N__43568),
            .in2(N__40236),
            .in3(N__41152),
            .lcout(M_this_ext_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42096),
            .ce(),
            .sr(N__43097));
    defparam M_this_ext_address_q_15_LC_26_18_3.C_ON=1'b0;
    defparam M_this_ext_address_q_15_LC_26_18_3.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_15_LC_26_18_3.LUT_INIT=16'b1110111101000000;
    LogicCell40 M_this_ext_address_q_15_LC_26_18_3 (
            .in0(N__41151),
            .in1(N__39838),
            .in2(N__43576),
            .in3(N__41035),
            .lcout(M_this_ext_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42096),
            .ce(),
            .sr(N__43097));
    defparam M_this_ctrl_flags_q_6_LC_26_18_5.C_ON=1'b0;
    defparam M_this_ctrl_flags_q_6_LC_26_18_5.SEQ_MODE=4'b1000;
    defparam M_this_ctrl_flags_q_6_LC_26_18_5.LUT_INIT=16'b1110010011001100;
    LogicCell40 M_this_ctrl_flags_q_6_LC_26_18_5 (
            .in0(N__43565),
            .in1(N__40458),
            .in2(N__40419),
            .in3(N__40891),
            .lcout(M_this_ctrl_flags_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42096),
            .ce(),
            .sr(N__43097));
    defparam M_this_ext_address_q_14_LC_26_18_6.C_ON=1'b0;
    defparam M_this_ext_address_q_14_LC_26_18_6.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_14_LC_26_18_6.LUT_INIT=16'b1010111010100010;
    LogicCell40 M_this_ext_address_q_14_LC_26_18_6 (
            .in0(N__40519),
            .in1(N__43567),
            .in2(N__41161),
            .in3(N__40404),
            .lcout(M_this_ext_address_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42096),
            .ce(),
            .sr(N__43097));
    defparam un1_M_this_ext_address_q_cry_0_c_LC_26_21_0.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_0_c_LC_26_21_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_0_c_LC_26_21_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_ext_address_q_cry_0_c_LC_26_21_0 (
            .in0(_gnd_net_),
            .in1(N__40311),
            .in2(N__40280),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_26_21_0_),
            .carryout(un1_M_this_ext_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_0_THRU_LUT4_0_LC_26_21_1.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_0_THRU_LUT4_0_LC_26_21_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_0_THRU_LUT4_0_LC_26_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_0_THRU_LUT4_0_LC_26_21_1 (
            .in0(_gnd_net_),
            .in1(N__41288),
            .in2(_gnd_net_),
            .in3(N__40249),
            .lcout(un1_M_this_ext_address_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_0),
            .carryout(un1_M_this_ext_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_1_THRU_LUT4_0_LC_26_21_2.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_1_THRU_LUT4_0_LC_26_21_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_1_THRU_LUT4_0_LC_26_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_1_THRU_LUT4_0_LC_26_21_2 (
            .in0(_gnd_net_),
            .in1(N__40232),
            .in2(_gnd_net_),
            .in3(N__40201),
            .lcout(un1_M_this_ext_address_q_cry_1_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_1),
            .carryout(un1_M_this_ext_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_2_THRU_LUT4_0_LC_26_21_3.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_2_THRU_LUT4_0_LC_26_21_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_2_THRU_LUT4_0_LC_26_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_2_THRU_LUT4_0_LC_26_21_3 (
            .in0(_gnd_net_),
            .in1(N__41249),
            .in2(_gnd_net_),
            .in3(N__40198),
            .lcout(un1_M_this_ext_address_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_2),
            .carryout(un1_M_this_ext_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_3_THRU_LUT4_0_LC_26_21_4.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_3_THRU_LUT4_0_LC_26_21_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_3_THRU_LUT4_0_LC_26_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_3_THRU_LUT4_0_LC_26_21_4 (
            .in0(_gnd_net_),
            .in1(N__41213),
            .in2(_gnd_net_),
            .in3(N__40195),
            .lcout(un1_M_this_ext_address_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_3),
            .carryout(un1_M_this_ext_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_4_THRU_LUT4_0_LC_26_21_5.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_4_THRU_LUT4_0_LC_26_21_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_4_THRU_LUT4_0_LC_26_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_4_THRU_LUT4_0_LC_26_21_5 (
            .in0(_gnd_net_),
            .in1(N__41177),
            .in2(_gnd_net_),
            .in3(N__40192),
            .lcout(un1_M_this_ext_address_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_4),
            .carryout(un1_M_this_ext_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_5_THRU_LUT4_0_LC_26_21_6.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_5_THRU_LUT4_0_LC_26_21_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_5_THRU_LUT4_0_LC_26_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_5_THRU_LUT4_0_LC_26_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43275),
            .in3(N__40189),
            .lcout(un1_M_this_ext_address_q_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_5),
            .carryout(un1_M_this_ext_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_6_THRU_LUT4_0_LC_26_21_7.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_6_THRU_LUT4_0_LC_26_21_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_6_THRU_LUT4_0_LC_26_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_6_THRU_LUT4_0_LC_26_21_7 (
            .in0(_gnd_net_),
            .in1(N__40971),
            .in2(_gnd_net_),
            .in3(N__40642),
            .lcout(un1_M_this_ext_address_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_6),
            .carryout(un1_M_this_ext_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_7_c_RNIQ14F_LC_26_22_0.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_7_c_RNIQ14F_LC_26_22_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_7_c_RNIQ14F_LC_26_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_7_c_RNIQ14F_LC_26_22_0 (
            .in0(_gnd_net_),
            .in1(N__41322),
            .in2(_gnd_net_),
            .in3(N__40639),
            .lcout(un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0),
            .ltout(),
            .carryin(bfn_26_22_0_),
            .carryout(un1_M_this_ext_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_8_c_RNIS45F_LC_26_22_1.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_8_c_RNIS45F_LC_26_22_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_8_c_RNIS45F_LC_26_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_8_c_RNIS45F_LC_26_22_1 (
            .in0(_gnd_net_),
            .in1(N__40626),
            .in2(_gnd_net_),
            .in3(N__40594),
            .lcout(un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_8),
            .carryout(un1_M_this_ext_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_9_c_RNI55NH_LC_26_22_2.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_9_c_RNI55NH_LC_26_22_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_9_c_RNI55NH_LC_26_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_9_c_RNI55NH_LC_26_22_2 (
            .in0(_gnd_net_),
            .in1(N__41004),
            .in2(_gnd_net_),
            .in3(N__40591),
            .lcout(un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_9),
            .carryout(un1_M_this_ext_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_10_c_RNIEGOA_LC_26_22_3.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_10_c_RNIEGOA_LC_26_22_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_10_c_RNIEGOA_LC_26_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_10_c_RNIEGOA_LC_26_22_3 (
            .in0(_gnd_net_),
            .in1(N__40929),
            .in2(_gnd_net_),
            .in3(N__40588),
            .lcout(un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_10),
            .carryout(un1_M_this_ext_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_11_c_RNIGJPA_LC_26_22_4.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_11_c_RNIGJPA_LC_26_22_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_11_c_RNIGJPA_LC_26_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_11_c_RNIGJPA_LC_26_22_4 (
            .in0(_gnd_net_),
            .in1(N__40902),
            .in2(_gnd_net_),
            .in3(N__40585),
            .lcout(un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_11),
            .carryout(un1_M_this_ext_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_12_c_RNIIMQA_LC_26_22_5.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_12_c_RNIIMQA_LC_26_22_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_12_c_RNIIMQA_LC_26_22_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_12_c_RNIIMQA_LC_26_22_5 (
            .in0(_gnd_net_),
            .in1(N__40572),
            .in2(_gnd_net_),
            .in3(N__40546),
            .lcout(un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_12),
            .carryout(un1_M_this_ext_address_q_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_13_c_RNIKPRA_LC_26_22_6.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_13_c_RNIKPRA_LC_26_22_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_13_c_RNIKPRA_LC_26_22_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_13_c_RNIKPRA_LC_26_22_6 (
            .in0(_gnd_net_),
            .in1(N__40536),
            .in2(_gnd_net_),
            .in3(N__40510),
            .lcout(un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_13),
            .carryout(un1_M_this_ext_address_q_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_14_c_RNIMSSA_LC_26_22_7.C_ON=1'b0;
    defparam un1_M_this_ext_address_q_cry_14_c_RNIMSSA_LC_26_22_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_14_c_RNIMSSA_LC_26_22_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_M_this_ext_address_q_cry_14_c_RNIMSSA_LC_26_22_7 (
            .in0(_gnd_net_),
            .in1(N__40503),
            .in2(_gnd_net_),
            .in3(N__41038),
            .lcout(un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_ext_address_q_10_LC_26_23_0.C_ON=1'b0;
    defparam M_this_ext_address_q_10_LC_26_23_0.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_10_LC_26_23_0.LUT_INIT=16'b1011100010101010;
    LogicCell40 M_this_ext_address_q_10_LC_26_23_0 (
            .in0(N__41026),
            .in1(N__41097),
            .in2(N__42757),
            .in3(N__43561),
            .lcout(M_this_ext_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42125),
            .ce(),
            .sr(N__43102));
    defparam M_this_ext_address_q_7_LC_26_23_1.C_ON=1'b0;
    defparam M_this_ext_address_q_7_LC_26_23_1.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_7_LC_26_23_1.LUT_INIT=16'b0010001110001100;
    LogicCell40 M_this_ext_address_q_7_LC_26_23_1 (
            .in0(N__41096),
            .in1(N__40967),
            .in2(N__43575),
            .in3(N__40993),
            .lcout(M_this_ext_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42125),
            .ce(),
            .sr(N__43102));
    defparam M_this_ext_address_q_11_LC_26_23_2.C_ON=1'b0;
    defparam M_this_ext_address_q_11_LC_26_23_2.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_11_LC_26_23_2.LUT_INIT=16'b1010110010101010;
    LogicCell40 M_this_ext_address_q_11_LC_26_23_2 (
            .in0(N__40948),
            .in1(N__41454),
            .in2(N__41129),
            .in3(N__43562),
            .lcout(M_this_ext_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42125),
            .ce(),
            .sr(N__43102));
    defparam M_this_ext_address_q_12_LC_26_23_3.C_ON=1'b0;
    defparam M_this_ext_address_q_12_LC_26_23_3.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_12_LC_26_23_3.LUT_INIT=16'b1110111101000000;
    LogicCell40 M_this_ext_address_q_12_LC_26_23_3 (
            .in0(N__41095),
            .in1(N__40709),
            .in2(N__43574),
            .in3(N__40918),
            .lcout(M_this_ext_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42125),
            .ce(),
            .sr(N__43102));
    defparam M_this_ctrl_flags_q_4_LC_26_23_4.C_ON=1'b0;
    defparam M_this_ctrl_flags_q_4_LC_26_23_4.SEQ_MODE=4'b1000;
    defparam M_this_ctrl_flags_q_4_LC_26_23_4.LUT_INIT=16'b1110010011001100;
    LogicCell40 M_this_ctrl_flags_q_4_LC_26_23_4 (
            .in0(N__40881),
            .in1(N__40839),
            .in2(N__40726),
            .in3(N__43563),
            .lcout(M_this_ctrl_flags_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42125),
            .ce(),
            .sr(N__43102));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_9_LC_26_24_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_9_LC_26_24_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_9_LC_26_24_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a3_9_LC_26_24_5  (
            .in0(_gnd_net_),
            .in1(N__40812),
            .in2(_gnd_net_),
            .in3(N__42828),
            .lcout(),
            .ltout(N_1081_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_0_9_LC_26_24_6.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_0_9_LC_26_24_6.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_0_9_LC_26_24_6.LUT_INIT=16'b0000000000001011;
    LogicCell40 M_this_map_address_q_RNO_0_9_LC_26_24_6 (
            .in0(N__40705),
            .in1(N__42593),
            .in2(N__40654),
            .in3(N__42543),
            .lcout(M_this_map_address_qc_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_5_LC_26_25_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_5_LC_26_25_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_5_LC_26_25_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a3_5_LC_26_25_4  (
            .in0(_gnd_net_),
            .in1(N__42167),
            .in2(_gnd_net_),
            .in3(N__42829),
            .lcout(N_1068),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_8_LC_26_25_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_8_LC_26_25_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_8_LC_26_25_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a3_8_LC_26_25_5  (
            .in0(N__42830),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41549),
            .lcout(),
            .ltout(N_1078_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_0_8_LC_26_25_6.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_0_8_LC_26_25_6.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_0_8_LC_26_25_6.LUT_INIT=16'b0000001000000011;
    LogicCell40 M_this_map_address_q_RNO_0_8_LC_26_25_6 (
            .in0(N__41470),
            .in1(N__42540),
            .in2(N__41386),
            .in3(N__42594),
            .lcout(M_this_map_address_qc_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_2_LC_26_30_6 .C_ON=1'b0;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_2_LC_26_30_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_2_LC_26_30_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.IO_port_data_write_0_a2_i_2_LC_26_30_6  (
            .in0(N__43703),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41364),
            .lcout(N_726_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_ext_address_q_8_LC_27_22_0.C_ON=1'b0;
    defparam M_this_ext_address_q_8_LC_27_22_0.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_8_LC_27_22_0.LUT_INIT=16'b1011100010101010;
    LogicCell40 M_this_ext_address_q_8_LC_27_22_0 (
            .in0(N__41341),
            .in1(N__41133),
            .in2(N__42463),
            .in3(N__43545),
            .lcout(M_this_ext_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42126),
            .ce(),
            .sr(N__43099));
    defparam M_this_ext_address_q_1_LC_27_22_2.C_ON=1'b0;
    defparam M_this_ext_address_q_1_LC_27_22_2.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_1_LC_27_22_2.LUT_INIT=16'b0100100001011010;
    LogicCell40 M_this_ext_address_q_1_LC_27_22_2 (
            .in0(N__41311),
            .in1(N__41134),
            .in2(N__41295),
            .in3(N__43546),
            .lcout(M_this_ext_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42126),
            .ce(),
            .sr(N__43099));
    defparam M_this_ext_address_q_3_LC_27_22_4.C_ON=1'b0;
    defparam M_this_ext_address_q_3_LC_27_22_4.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_3_LC_27_22_4.LUT_INIT=16'b0100100001011010;
    LogicCell40 M_this_ext_address_q_3_LC_27_22_4 (
            .in0(N__41272),
            .in1(N__41135),
            .in2(N__41256),
            .in3(N__43547),
            .lcout(M_this_ext_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42126),
            .ce(),
            .sr(N__43099));
    defparam M_this_ext_address_q_4_LC_27_22_5.C_ON=1'b0;
    defparam M_this_ext_address_q_4_LC_27_22_5.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_4_LC_27_22_5.LUT_INIT=16'b0010001110001100;
    LogicCell40 M_this_ext_address_q_4_LC_27_22_5 (
            .in0(N__41131),
            .in1(N__41214),
            .in2(N__43572),
            .in3(N__41233),
            .lcout(M_this_ext_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42126),
            .ce(),
            .sr(N__43099));
    defparam M_this_ext_address_q_5_LC_27_22_6.C_ON=1'b0;
    defparam M_this_ext_address_q_5_LC_27_22_6.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_5_LC_27_22_6.LUT_INIT=16'b0100100001011010;
    LogicCell40 M_this_ext_address_q_5_LC_27_22_6 (
            .in0(N__41197),
            .in1(N__41136),
            .in2(N__41184),
            .in3(N__43548),
            .lcout(M_this_ext_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42126),
            .ce(),
            .sr(N__43099));
    defparam M_this_ext_address_q_6_LC_27_22_7.C_ON=1'b0;
    defparam M_this_ext_address_q_6_LC_27_22_7.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_6_LC_27_22_7.LUT_INIT=16'b0010001110001100;
    LogicCell40 M_this_ext_address_q_6_LC_27_22_7 (
            .in0(N__41132),
            .in1(N__43271),
            .in2(N__43573),
            .in3(N__43285),
            .lcout(M_this_ext_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42126),
            .ce(),
            .sr(N__43099));
    defparam M_this_map_address_q_7_LC_27_23_3.C_ON=1'b0;
    defparam M_this_map_address_q_7_LC_27_23_3.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_7_LC_27_23_3.LUT_INIT=16'b0010100010101010;
    LogicCell40 M_this_map_address_q_7_LC_27_23_3 (
            .in0(N__42655),
            .in1(N__42895),
            .in2(N__42870),
            .in3(N__42293),
            .lcout(M_this_map_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42132),
            .ce(),
            .sr(N__41650));
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_7_LC_27_24_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_7_LC_27_24_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_0_a3_7_LC_27_24_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_0_a3_7_LC_27_24_0  (
            .in0(_gnd_net_),
            .in1(N__42859),
            .in2(_gnd_net_),
            .in3(N__42835),
            .lcout(),
            .ltout(N_1075_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_0_7_LC_27_24_1.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_0_7_LC_27_24_1.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_0_7_LC_27_24_1.LUT_INIT=16'b0000000000001011;
    LogicCell40 M_this_map_address_q_RNO_0_7_LC_27_24_1 (
            .in0(N__42710),
            .in1(N__42595),
            .in2(N__42658),
            .in3(N__42544),
            .lcout(M_this_map_address_qc_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_substate_d_0_sqmuxa_3_0_o2_LC_27_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_substate_d_0_sqmuxa_3_0_o2_LC_27_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_substate_d_0_sqmuxa_3_0_o2_LC_27_24_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_substate_d_0_sqmuxa_3_0_o2_LC_27_24_3  (
            .in0(N__43854),
            .in1(N__42636),
            .in2(N__43887),
            .in3(N__43813),
            .lcout(N_459_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_RNO_0_5_LC_27_25_5.C_ON=1'b0;
    defparam M_this_map_address_q_RNO_0_5_LC_27_25_5.SEQ_MODE=4'b0000;
    defparam M_this_map_address_q_RNO_0_5_LC_27_25_5.LUT_INIT=16'b0000000000110001;
    LogicCell40 M_this_map_address_q_RNO_0_5_LC_27_25_5 (
            .in0(N__42592),
            .in1(N__42539),
            .in2(N__42459),
            .in3(N__42319),
            .lcout(M_this_map_address_qc_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_5_LC_27_26_2.C_ON=1'b0;
    defparam M_this_map_address_q_5_LC_27_26_2.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_5_LC_27_26_2.LUT_INIT=16'b1000100010101010;
    LogicCell40 M_this_map_address_q_5_LC_27_26_2 (
            .in0(N__42313),
            .in1(N__42307),
            .in2(_gnd_net_),
            .in3(N__42294),
            .lcout(M_this_map_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42137),
            .ce(),
            .sr(N__41646));
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_6_LC_28_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_6_LC_28_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_6_LC_28_19_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.IO_port_data_write_0_a2_i_6_LC_28_19_5  (
            .in0(N__43696),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41601),
            .lcout(N_734_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_5_LC_28_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_5_LC_28_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_5_LC_28_19_6 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \this_vga_signals.IO_port_data_write_0_a2_i_5_LC_28_19_6  (
            .in0(N__43936),
            .in1(N__43695),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_996_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_substate_d_0_sqmuxa_3_0_o2_x_LC_28_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_substate_d_0_sqmuxa_3_0_o2_x_LC_28_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_substate_d_0_sqmuxa_3_0_o2_x_LC_28_23_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_this_substate_d_0_sqmuxa_3_0_o2_x_LC_28_23_7  (
            .in0(N__43874),
            .in1(N__43847),
            .in2(_gnd_net_),
            .in3(N__43806),
            .lcout(M_this_substate_d_0_sqmuxa_3_0_o2_x),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_4_LC_28_27_5 .C_ON=1'b0;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_4_LC_28_27_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_4_LC_28_27_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.IO_port_data_write_0_a2_i_4_LC_28_27_5  (
            .in0(N__43704),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43746),
            .lcout(N_730_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_3_LC_28_29_1 .C_ON=1'b0;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_3_LC_28_29_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.IO_port_data_write_0_a2_i_3_LC_28_29_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.IO_port_data_write_0_a2_i_3_LC_28_29_1  (
            .in0(N__43705),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43608),
            .lcout(N_728_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
