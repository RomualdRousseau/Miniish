-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 10 2022 20:23:05

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \VCCG0\ : std_logic;
signal \N_377_i\ : std_logic;
signal port_nmib_0_i : std_logic;
signal port_clk_c : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal rgb_c_0 : std_logic;
signal i7_mux_0 : std_logic;
signal rgb_c_1 : std_logic;
signal \N_28_0\ : std_logic;
signal rgb_c_5 : std_logic;
signal \this_vga_signals.new_pixel_1_1_cascade_\ : std_logic;
signal \debug_c_0_cascade_\ : std_logic;
signal rgb_c_3 : std_logic;
signal \N_37\ : std_logic;
signal rgb_c_4 : std_logic;
signal \this_vga_signals.new_pixel_1_3_1_cascade_\ : std_logic;
signal \this_vga_signals.new_pixel_sx_0\ : std_logic;
signal this_vga_signals_vvisibility_i : std_logic;
signal \N_60\ : std_logic;
signal i7_mux : std_logic;
signal \N_50_cascade_\ : std_logic;
signal debug_c_0 : std_logic;
signal rgb_c_2 : std_logic;
signal \M_hcounter_q_esr_RNIH8GJ4_9\ : std_logic;
signal \bfn_6_21_0_\ : std_logic;
signal \this_vga_signals.new_pixel_1Z0Z_1\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_0\ : std_logic;
signal \this_vga_signals.new_pixel_1_2\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_1\ : std_logic;
signal \this_vga_signals.new_pixel_1_3\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_2\ : std_logic;
signal \this_vga_signals.new_pixel_1_4\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_3\ : std_logic;
signal \this_vga_signals.new_pixel_1_5\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_4\ : std_logic;
signal \this_vga_signals.new_pixel_1_6\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_5\ : std_logic;
signal \this_vga_signals.M_hcounter_q_i_7\ : std_logic;
signal \this_vga_signals.new_pixel_1_7\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_6\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_7\ : std_logic;
signal \this_vga_signals.new_pixel_1_8\ : std_logic;
signal \bfn_6_22_0_\ : std_logic;
signal \this_vga_signals.new_pixel_1_9\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_8\ : std_logic;
signal \this_vga_signals.new_pixel_1_10\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_9\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_10\ : std_logic;
signal \this_vga_signals.new_pixel_1_11\ : std_logic;
signal \this_vga_signals.un4_hsynclt8_0\ : std_logic;
signal this_vga_signals_hsync_1_i : std_logic;
signal debug_c_i_1 : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNIG53K_1Z0Z_9\ : std_logic;
signal \this_vga_signals.un3_hsynclt8_0\ : std_logic;
signal \this_vga_signals.new_pixel_1_i_0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNIUA42NDZ0Z_1\ : std_logic;
signal \this_vga_signals.new_pixel_1_cry_0_c_RNOZ0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNIG53KZ0Z_9\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_\ : std_logic;
signal \this_vga_signals.g0_13_N_3L3_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_2_0_0\ : std_logic;
signal \this_vga_signals.g0_13_N_3L3_x1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_cascade_\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \this_vga_signals.M_hcounter_d6lt9_cascade_\ : std_logic;
signal \this_pixel_clock_M_counter_q_i_1\ : std_logic;
signal \this_pixel_clock_M_counter_q_0\ : std_logic;
signal \this_vga_signals.M_hcounter_d6_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNIUKG82Z0Z_9\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_1_sx_cascade_\ : std_logic;
signal \this_vga_signals.if_m2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_i_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_1\ : std_logic;
signal \this_vga_signals.N_4_i_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_ac0_1_cascade_\ : std_logic;
signal \this_vga_signals.N_4_i\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9_cascade_\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TAZ0Z7\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_i_0_3\ : std_logic;
signal \this_vga_signals.un1_haddress_0_axb_2_l_ofxZ0\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44VZ0Z02\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_1\ : std_logic;
signal \this_vga_signals.un1_haddress_0_axb_3_l_fxZ0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_i_3\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9DZ0\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_2\ : std_logic;
signal \this_vga_signals.un1_haddress_0_axb_4_l_fxZ0\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4TZ0Z72\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_3\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJLZ0\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_4\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_5_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_5\ : std_logic;
signal \this_vga_signals.un1_haddress_0_axb_7\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQUZ0\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_6\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_7_i\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_7\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBSZ0Z7\ : std_logic;
signal \this_vga_signals.m8_0_1_tz_cascade_\ : std_logic;
signal \this_vga_signals.g1_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_0_cascade_\ : std_logic;
signal \this_vga_signals.N_75_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_m_1_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_m_1_1_cascade_\ : std_logic;
signal \this_vga_signals.N_75\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_m_x0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_m_x1_1\ : std_logic;
signal \this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOMZ0Z71_cascade_\ : std_logic;
signal \this_vga_signals.m8_0_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_i_0_3_cascade_\ : std_logic;
signal \this_vga_signals.g1_6_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3\ : std_logic;
signal \this_vga_signals.g0_13_N_3L3_ns\ : std_logic;
signal \this_vga_signals.g0_13_N_2L1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_0_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5\ : std_logic;
signal \this_vga_signals.if_m2_0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5_cascade_\ : std_logic;
signal \this_vga_signals.g0_10_3_0_a2_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_1\ : std_logic;
signal \this_vga_signals.g1_0\ : std_logic;
signal \this_vga_signals.g0_10_3_0_a2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_x0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_x1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_i_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_3_0_1_x1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_3_0_1_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_3_0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_i\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc2\ : std_logic;
signal \this_vga_signals.N_510_i\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1_i_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_ac0_3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.new_pixel_1_axb_1_N_4L5_xZ0Z1_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNIPIQRNRZ0Z_2\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNI5HOBQCZ0Z_1\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNI8TTVN32Z0Z_2_cascade_\ : std_logic;
signal \this_vga_signals.new_pixel_1_axb_1\ : std_logic;
signal \this_vga_signals.N_510_cascade_\ : std_logic;
signal \this_vga_signals.un1_haddress_0_axb_6\ : std_logic;
signal \this_vga_signals.un1_haddress_0\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_\ : std_logic;
signal \this_vga_signals.un1_haddress_0_cry_1_c_RNOZ0\ : std_logic;
signal \this_vga_signals.m8_0_1_tz\ : std_logic;
signal \this_vga_signals.ANC2_4_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_q_7_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_hcounter_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fastZ0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.M_hcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_hcounter_q_9_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fast_esr_RNIHH441Z0Z_5_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fast_esr_RNIN6RRZ0Z_7\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.N_550_1\ : std_logic;
signal \this_vga_signals.m8_0_2\ : std_logic;
signal \this_vga_signals.g1_0_1\ : std_logic;
signal \this_vga_signals.g4_1_1_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fast_esr_RNI52HLZ0Z_9\ : std_logic;
signal \this_vga_signals.m8_0_1_0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_8_repZ0Z1\ : std_logic;
signal \this_vga_signals.m8_0_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3\ : std_logic;
signal \this_vga_signals.g1_1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_2_0\ : std_logic;
signal \this_vga_signals.g1_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_6_0\ : std_logic;
signal \this_vga_signals.g4_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_1_1\ : std_logic;
signal \this_vga_signals.g0_13_N_4L5\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_1_3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_i_1_0_0\ : std_logic;
signal \this_vga_signals.g4\ : std_logic;
signal \this_vga_signals.g0_0_2_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_1_0_0\ : std_logic;
signal \this_vga_signals.N_4_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_0_3_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_a2_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3\ : std_logic;
signal \this_vga_signals.N_19\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_3_0_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_i_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_1_0\ : std_logic;
signal \this_vga_signals.g0_i_x2_0_0_a2_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.if_i4_mux_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_a2\ : std_logic;
signal \this_vga_signals.g0_i_x2_0_0_a2_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0\ : std_logic;
signal \this_vga_signals.g1_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_0_3\ : std_logic;
signal \this_vga_signals.g0_0_a2_4\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axb2_i\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_ac0_3_0_0\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1_i\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_i_0_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_m_ns_1\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \this_vga_signals.new_pixel_1\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.N_583_g\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRDZ0\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.g0_4_0\ : std_logic;
signal debug_c_1 : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.g0_0_a2_1\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_1_2\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_1_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c2\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_4\ : std_logic;
signal \this_vga_signals.un2_vsynclt8\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \M_this_vga_signals_address_6\ : std_logic;
signal \this_vga_signals.if_N_9\ : std_logic;
signal \this_vga_signals.if_N_10_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_i\ : std_logic;
signal \this_vga_signals.SUM_2\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c2\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axb2_0_3\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c2_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axb2_3_tz\ : std_logic;
signal \this_vga_signals.vaddress_7\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt8_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt9_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lto8_1\ : std_logic;
signal \this_vga_signals.un6_vvisibilitylt9_0_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_c5_i\ : std_logic;
signal \this_vga_signals.vvisibility\ : std_logic;
signal \this_vga_signals.vsync_1_0_cascade_\ : std_logic;
signal \this_vga_signals.vsync_1_4\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_ns_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_cascade_\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_i_1_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3\ : std_logic;
signal \M_this_vga_signals_address_10\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_bm\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2\ : std_logic;
signal \this_vga_signals.if_N_10\ : std_logic;
signal \M_this_vga_signals_address_9\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc2_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc2\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0_0\ : std_logic;
signal \M_this_vga_signals_address_8\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_ns_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axb2_0_3_1_1\ : std_logic;
signal \this_vga_signals.M_hcounter_d6_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \this_vga_signals.GZ0Z_296\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_0_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_1_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_2_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_3_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_4_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_5_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c2\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_i_3\ : std_logic;
signal \this_vga_signals.vaddress_8\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x1\ : std_logic;
signal port_dmab_c_i : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal \un1_M_this_data_count_q_cry_0\ : std_logic;
signal \un1_M_this_data_count_q_cry_1\ : std_logic;
signal \un1_M_this_data_count_q_cry_2\ : std_logic;
signal \un1_M_this_data_count_q_cry_3\ : std_logic;
signal \un1_M_this_data_count_q_cry_4\ : std_logic;
signal \un1_M_this_data_count_q_cry_5\ : std_logic;
signal \un1_M_this_data_count_q_cry_6\ : std_logic;
signal \un1_M_this_data_count_q_cry_7\ : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal \un1_M_this_data_count_q_cry_8\ : std_logic;
signal \un1_M_this_data_count_q_cry_9\ : std_logic;
signal \un1_M_this_data_count_q_cry_10\ : std_logic;
signal \un1_M_this_data_count_q_cry_11\ : std_logic;
signal \un1_M_this_data_count_q_cry_12\ : std_logic;
signal \un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO\ : std_logic;
signal \GNDG0\ : std_logic;
signal \un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO\ : std_logic;
signal \un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO\ : std_logic;
signal \bfn_16_25_0_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_1_c2_1_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2Z0Z_9\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_1_c2_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.mult1_un54_sum1_i_1_3\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \this_vga_signals.vaddress_c2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_3\ : std_logic;
signal \this_vga_signals.N_550_2\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.N_550_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_i_1_2_cascade_\ : std_logic;
signal \this_start_data_delay.N_389_1\ : std_logic;
signal port_dmab_c : std_logic;
signal \port_dmab_c_cascade_\ : std_logic;
signal \this_start_data_delay.N_385_cascade_\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_i_a2_1_9Z0Z_1\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_i_a2_1_6Z0Z_1_cascade_\ : std_logic;
signal \this_start_data_delay.N_413\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_i_a2_1_8Z0Z_1\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_i_a2_1_7Z0Z_1\ : std_logic;
signal \M_this_state_q_RNI20CEZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \M_this_state_q_nss_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \this_start_data_delay.N_353_0\ : std_logic;
signal \M_this_start_data_delay_out_0_cascade_\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_11\ : std_logic;
signal port_rw_in : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_0_a2_1_4\ : std_logic;
signal \this_start_data_delay.N_352_0_cascade_\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_0_0_4\ : std_logic;
signal port_enb_c : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal \this_start_data_delay.M_last_qZ0\ : std_logic;
signal \this_start_data_delay.N_352_0\ : std_logic;
signal \this_start_data_delay.N_407_cascade_\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_1\ : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_4\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_9\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_2\ : std_logic;
signal \this_start_data_delay.N_407\ : std_logic;
signal \this_start_data_delay.N_398\ : std_logic;
signal \this_start_data_delay.M_this_state_dZ0Z29\ : std_logic;
signal \this_start_data_delay.N_396\ : std_logic;
signal \this_start_data_delay.M_this_state_dZ0Z27\ : std_logic;
signal port_address_in_0 : std_logic;
signal port_address_in_1 : std_logic;
signal \this_start_data_delay.M_this_state_dZ0Z28\ : std_logic;
signal \M_this_vga_signals_address_13\ : std_logic;
signal \M_this_vga_signals_address_12\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_5\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_3\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_7\ : std_logic;
signal \N_346_0\ : std_logic;
signal \M_this_internal_address_q_RNI6EA12Z0Z_0\ : std_logic;
signal \bfn_20_21_0_\ : std_logic;
signal \M_this_internal_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_internal_address_q_cry_0_c_RNI4MQIZ0\ : std_logic;
signal \un1_M_this_internal_address_q_cry_0\ : std_logic;
signal \M_this_internal_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_internal_address_q_cry_1_c_RNI6PRIZ0\ : std_logic;
signal \un1_M_this_internal_address_q_cry_1\ : std_logic;
signal \M_this_internal_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_internal_address_q_cry_2_c_RNI8SSIZ0\ : std_logic;
signal \un1_M_this_internal_address_q_cry_2\ : std_logic;
signal \M_this_internal_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_internal_address_q_cry_3_c_RNIAVTIZ0\ : std_logic;
signal \un1_M_this_internal_address_q_cry_3\ : std_logic;
signal \M_this_internal_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_internal_address_q_cry_4_c_RNIC2VIZ0\ : std_logic;
signal \un1_M_this_internal_address_q_cry_4\ : std_logic;
signal \un1_M_this_internal_address_q_cry_5\ : std_logic;
signal \M_this_internal_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_internal_address_q_cry_6_c_RNIG81JZ0\ : std_logic;
signal \un1_M_this_internal_address_q_cry_6\ : std_logic;
signal \un1_M_this_internal_address_q_cry_7\ : std_logic;
signal \bfn_20_22_0_\ : std_logic;
signal \M_this_internal_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_internal_address_q_cry_8_c_RNIKE3JZ0\ : std_logic;
signal \un1_M_this_internal_address_q_cry_8\ : std_logic;
signal \un1_M_this_internal_address_q_cry_9\ : std_logic;
signal \un1_M_this_internal_address_q_cry_10_c_RNI6I0DZ0\ : std_logic;
signal \un1_M_this_internal_address_q_cry_10\ : std_logic;
signal \un1_M_this_internal_address_q_cry_11\ : std_logic;
signal \un1_M_this_internal_address_q_cry_12\ : std_logic;
signal \M_this_internal_address_qZ0Z_0\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_0\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_10\ : std_logic;
signal \un1_M_this_internal_address_q_cry_9_c_RNITQCIZ0\ : std_logic;
signal \M_this_internal_address_qZ0Z_10\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_12\ : std_logic;
signal \un1_M_this_internal_address_q_cry_11_c_RNI8L1DZ0\ : std_logic;
signal \un1_M_this_internal_address_q_cry_5_c_RNIE50JZ0\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_13\ : std_logic;
signal \un1_M_this_internal_address_q_cry_12_c_RNIAO2DZ0\ : std_logic;
signal \un1_M_this_internal_address_q_cry_7_c_RNIIB2JZ0\ : std_logic;
signal \M_this_internal_address_q_3_sm0_0\ : std_logic;
signal \this_vram.mem_out_bus4_1\ : std_logic;
signal \this_vram.mem_out_bus0_1\ : std_logic;
signal \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_11\ : std_logic;
signal \this_vram.mem_DOUT_7_i_m2_ns_1_1\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \M_this_internal_address_qZ0Z_6\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_6\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal \M_this_internal_address_qZ0Z_8\ : std_logic;
signal \this_vram.M_this_internal_address_q_3_ns_1Z0Z_8\ : std_logic;
signal port_address_in_3 : std_logic;
signal port_address_in_2 : std_logic;
signal \this_start_data_delay.M_this_state_d27Z0Z_2\ : std_logic;
signal \this_vram.mem_WE_14\ : std_logic;
signal \this_vram.mem_out_bus6_1\ : std_logic;
signal \this_vram.mem_out_bus2_1\ : std_logic;
signal \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus7_1\ : std_logic;
signal \this_vram.mem_out_bus3_1\ : std_logic;
signal \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \this_vram.mem_DOUT_7_i_m2_ns_1_2_cascade_\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \this_vram.mem_radregZ0Z_11\ : std_logic;
signal \this_vram.mem_DOUT_7_i_m2_ns_1_0\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal port_data_c_1 : std_logic;
signal port_data_c_5 : std_logic;
signal \M_this_vram_write_data_0_i_1\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal port_data_c_0 : std_logic;
signal port_data_c_4 : std_logic;
signal \M_this_vram_write_data_0_sqmuxa_cascade_\ : std_logic;
signal \M_this_vram_write_data_0_i_0\ : std_logic;
signal \M_this_start_data_delay_out_0\ : std_logic;
signal \this_start_data_delay.N_351_0\ : std_logic;
signal \this_vram.mem_WE_8\ : std_logic;
signal \this_vram.mem_WE_12\ : std_logic;
signal \this_vram.mem_WE_10\ : std_logic;
signal \this_vram.mem_out_bus4_2\ : std_logic;
signal \this_vram.mem_out_bus0_2\ : std_logic;
signal \this_vram.mem_mem_0_1_RNISOIZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus5_3\ : std_logic;
signal \this_vram.mem_out_bus1_3\ : std_logic;
signal \this_vram.mem_out_bus3_3\ : std_logic;
signal \this_vram.mem_out_bus7_3\ : std_logic;
signal \this_vram.mem_DOUT_6_i_m2_ns_1_3_cascade_\ : std_logic;
signal \this_vram.mem_N_102\ : std_logic;
signal \this_vram.mem_out_bus4_3\ : std_logic;
signal \this_vram.mem_out_bus0_3\ : std_logic;
signal \this_vram.mem_out_bus6_3\ : std_logic;
signal \this_vram.mem_out_bus2_3\ : std_logic;
signal \this_vram.mem_DOUT_3_i_m2_ns_1_3_cascade_\ : std_logic;
signal \this_vram.mem_radregZ0Z_12\ : std_logic;
signal \this_vram.mem_N_105\ : std_logic;
signal \this_vram.mem_out_bus0_0\ : std_logic;
signal \this_vram.mem_out_bus4_0\ : std_logic;
signal \this_vram.mem_mem_0_0_RNIQOIZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus6_0\ : std_logic;
signal \this_vram.mem_out_bus2_0\ : std_logic;
signal \this_vram.mem_mem_2_0_RNIU0NZ0Z11\ : std_logic;
signal \this_vram.mem_WE_6\ : std_logic;
signal \this_vram.mem_out_bus1_1\ : std_logic;
signal \this_vram.mem_out_bus5_1\ : std_logic;
signal \this_vram.mem_mem_1_0_RNISSK11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus5_2\ : std_logic;
signal \this_vram.mem_out_bus1_2\ : std_logic;
signal \this_vram.mem_mem_1_1_RNIUSKZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus7_2\ : std_logic;
signal \this_vram.mem_out_bus3_2\ : std_logic;
signal \this_vram.mem_mem_3_1_RNI25PZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus7_0\ : std_logic;
signal \this_vram.mem_out_bus3_0\ : std_logic;
signal \this_vram.mem_mem_3_0_RNI05PZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus2_2\ : std_logic;
signal \this_vram.mem_out_bus6_2\ : std_logic;
signal \this_vram.mem_mem_2_1_RNI01NZ0Z11\ : std_logic;
signal \this_vram.mem_radregZ0Z_13\ : std_logic;
signal \this_vram.mem_out_bus5_0\ : std_logic;
signal \this_vram.mem_out_bus1_0\ : std_logic;
signal \this_vram.mem_mem_1_0_RNISSKZ0Z11\ : std_logic;
signal port_data_c_3 : std_logic;
signal port_data_c_7 : std_logic;
signal \M_this_vram_write_data_0_i_3\ : std_logic;
signal \this_vram.mem_WE_4\ : std_logic;
signal port_data_c_2 : std_logic;
signal port_data_c_6 : std_logic;
signal \M_this_vram_write_data_0_sqmuxa\ : std_logic;
signal \this_start_data_delay.un1_M_this_state_q_0\ : std_logic;
signal \M_this_vram_write_data_0_i_2\ : std_logic;
signal \this_vram.mem_WE_0\ : std_logic;
signal \M_this_internal_address_qZ0Z_12\ : std_logic;
signal \M_this_internal_address_qZ0Z_11\ : std_logic;
signal \M_this_internal_address_qZ0Z_13\ : std_logic;
signal \M_this_vram_write_en_0_0\ : std_logic;
signal \this_vram.mem_WE_2\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal \M_this_external_address_qZ0Z_0\ : std_logic;
signal \bfn_30_23_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_external_address_q_cry_0\ : std_logic;
signal \M_this_external_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_external_address_q_cry_1\ : std_logic;
signal \M_this_external_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_external_address_q_cry_2\ : std_logic;
signal \M_this_external_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_external_address_q_cry_3\ : std_logic;
signal \M_this_external_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_external_address_q_cry_4\ : std_logic;
signal \M_this_external_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_5\ : std_logic;
signal \M_this_external_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_external_address_q_cry_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_7\ : std_logic;
signal \M_this_external_address_qZ0Z_8\ : std_logic;
signal \bfn_30_24_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_external_address_q_cry_8\ : std_logic;
signal \M_this_external_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_external_address_q_cry_9\ : std_logic;
signal \M_this_external_address_qZ0Z_11\ : std_logic;
signal \un1_M_this_external_address_q_cry_10\ : std_logic;
signal \M_this_external_address_qZ0Z_12\ : std_logic;
signal \un1_M_this_external_address_q_cry_11\ : std_logic;
signal \M_this_external_address_qZ0Z_13\ : std_logic;
signal \un1_M_this_external_address_q_cry_12\ : std_logic;
signal \M_this_external_address_qZ0Z_14\ : std_logic;
signal \un1_M_this_external_address_q_cry_13\ : std_logic;
signal \M_this_state_qZ0Z_0\ : std_logic;
signal \un1_M_this_external_address_q_cry_14\ : std_logic;
signal \M_this_external_address_qZ0Z_15\ : std_logic;
signal clk_0_c_g : std_logic;
signal \M_this_state_q_nss_g_0\ : std_logic;
signal port_address_in_5 : std_logic;
signal port_address_in_6 : std_logic;
signal port_address_in_7 : std_logic;
signal port_address_in_4 : std_logic;
signal \this_start_data_delay.M_this_state_d27Z0Z_6\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \this_vram.mem_out_bus0_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= \N__12467\&\N__12311\&\N__12131\&\N__12647\&\N__11732\&\N__13955\&\N__9974\&\N__8198\&\N__10370\&\N__10562\&\N__10784\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= \N__17300\&\N__16601\&\N__17642\&\N__16733\&\N__17879\&\N__16868\&\N__17000\&\N__17132\&\N__16256\&\N__16400\&\N__17450\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18184\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18887\&'0'&'0'&'0';
    \this_vram.mem_out_bus0_3\ <= \this_vram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_2\ <= \this_vram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_1_physical_RADDR_wire\ <= \N__12461\&\N__12305\&\N__12125\&\N__12641\&\N__11726\&\N__13949\&\N__9968\&\N__8192\&\N__10364\&\N__10556\&\N__10778\;
    \this_vram.mem_mem_0_1_physical_WADDR_wire\ <= \N__17294\&\N__16595\&\N__17636\&\N__16727\&\N__17873\&\N__16862\&\N__16994\&\N__17126\&\N__16250\&\N__16394\&\N__17444\;
    \this_vram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19442\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20855\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_1\ <= \this_vram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_0\ <= \this_vram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_0_physical_RADDR_wire\ <= \N__12455\&\N__12299\&\N__12119\&\N__12635\&\N__11720\&\N__13943\&\N__9962\&\N__8186\&\N__10358\&\N__10550\&\N__10772\;
    \this_vram.mem_mem_1_0_physical_WADDR_wire\ <= \N__17288\&\N__16589\&\N__17630\&\N__16721\&\N__17867\&\N__16856\&\N__16988\&\N__17120\&\N__16244\&\N__16388\&\N__17438\;
    \this_vram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18180\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18883\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_3\ <= \this_vram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_2\ <= \this_vram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_1_physical_RADDR_wire\ <= \N__12449\&\N__12293\&\N__12113\&\N__12629\&\N__11714\&\N__13937\&\N__9956\&\N__8180\&\N__10352\&\N__10544\&\N__10766\;
    \this_vram.mem_mem_1_1_physical_WADDR_wire\ <= \N__17282\&\N__16583\&\N__17624\&\N__16715\&\N__17861\&\N__16850\&\N__16982\&\N__17114\&\N__16238\&\N__16382\&\N__17432\;
    \this_vram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19438\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20851\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_1\ <= \this_vram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_0\ <= \this_vram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_0_physical_RADDR_wire\ <= \N__12443\&\N__12287\&\N__12107\&\N__12623\&\N__11708\&\N__13931\&\N__9950\&\N__8174\&\N__10346\&\N__10538\&\N__10760\;
    \this_vram.mem_mem_2_0_physical_WADDR_wire\ <= \N__17276\&\N__16577\&\N__17618\&\N__16709\&\N__17855\&\N__16844\&\N__16976\&\N__17108\&\N__16232\&\N__16376\&\N__17426\;
    \this_vram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18164\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18876\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_3\ <= \this_vram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_2\ <= \this_vram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_1_physical_RADDR_wire\ <= \N__12437\&\N__12281\&\N__12101\&\N__12617\&\N__11702\&\N__13925\&\N__9944\&\N__8168\&\N__10340\&\N__10532\&\N__10754\;
    \this_vram.mem_mem_2_1_physical_WADDR_wire\ <= \N__17270\&\N__16571\&\N__17612\&\N__16703\&\N__17849\&\N__16838\&\N__16970\&\N__17102\&\N__16226\&\N__16370\&\N__17420\;
    \this_vram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19431\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20844\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_1\ <= \this_vram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_0\ <= \this_vram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_0_physical_RADDR_wire\ <= \N__12431\&\N__12275\&\N__12095\&\N__12611\&\N__11696\&\N__13919\&\N__9938\&\N__8162\&\N__10334\&\N__10526\&\N__10748\;
    \this_vram.mem_mem_3_0_physical_WADDR_wire\ <= \N__17264\&\N__16565\&\N__17606\&\N__16697\&\N__17843\&\N__16832\&\N__16964\&\N__17096\&\N__16220\&\N__16364\&\N__17414\;
    \this_vram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18185\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18866\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_3\ <= \this_vram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_2\ <= \this_vram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_1_physical_RADDR_wire\ <= \N__12425\&\N__12269\&\N__12089\&\N__12605\&\N__11690\&\N__13913\&\N__9932\&\N__8156\&\N__10328\&\N__10520\&\N__10742\;
    \this_vram.mem_mem_3_1_physical_WADDR_wire\ <= \N__17258\&\N__16559\&\N__17600\&\N__16691\&\N__17837\&\N__16826\&\N__16958\&\N__17090\&\N__16214\&\N__16358\&\N__17408\;
    \this_vram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19421\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20834\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_1\ <= \this_vram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_0\ <= \this_vram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_0_physical_RADDR_wire\ <= \N__12419\&\N__12263\&\N__12083\&\N__12599\&\N__11684\&\N__13907\&\N__9926\&\N__8150\&\N__10322\&\N__10514\&\N__10736\;
    \this_vram.mem_mem_4_0_physical_WADDR_wire\ <= \N__17252\&\N__16553\&\N__17594\&\N__16685\&\N__17831\&\N__16820\&\N__16952\&\N__17084\&\N__16208\&\N__16352\&\N__17402\;
    \this_vram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18171\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18853\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_3\ <= \this_vram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_2\ <= \this_vram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_1_physical_RADDR_wire\ <= \N__12413\&\N__12257\&\N__12077\&\N__12593\&\N__11678\&\N__13901\&\N__9920\&\N__8144\&\N__10316\&\N__10508\&\N__10730\;
    \this_vram.mem_mem_4_1_physical_WADDR_wire\ <= \N__17246\&\N__16547\&\N__17588\&\N__16679\&\N__17825\&\N__16814\&\N__16946\&\N__17078\&\N__16202\&\N__16346\&\N__17396\;
    \this_vram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19388\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20801\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_1\ <= \this_vram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_0\ <= \this_vram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_0_physical_RADDR_wire\ <= \N__12407\&\N__12251\&\N__12071\&\N__12587\&\N__11672\&\N__13895\&\N__9914\&\N__8138\&\N__10310\&\N__10502\&\N__10724\;
    \this_vram.mem_mem_5_0_physical_WADDR_wire\ <= \N__17240\&\N__16541\&\N__17582\&\N__16673\&\N__17819\&\N__16808\&\N__16940\&\N__17072\&\N__16196\&\N__16340\&\N__17390\;
    \this_vram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18131\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18831\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_3\ <= \this_vram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_2\ <= \this_vram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_1_physical_RADDR_wire\ <= \N__12401\&\N__12245\&\N__12065\&\N__12581\&\N__11666\&\N__13889\&\N__9908\&\N__8132\&\N__10304\&\N__10496\&\N__10718\;
    \this_vram.mem_mem_5_1_physical_WADDR_wire\ <= \N__17234\&\N__16535\&\N__17576\&\N__16667\&\N__17813\&\N__16802\&\N__16934\&\N__17066\&\N__16190\&\N__16334\&\N__17384\;
    \this_vram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19402\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20815\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_1\ <= \this_vram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_0\ <= \this_vram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_0_physical_RADDR_wire\ <= \N__12395\&\N__12239\&\N__12059\&\N__12575\&\N__11660\&\N__13883\&\N__9902\&\N__8126\&\N__10298\&\N__10490\&\N__10712\;
    \this_vram.mem_mem_6_0_physical_WADDR_wire\ <= \N__17228\&\N__16529\&\N__17570\&\N__16661\&\N__17807\&\N__16796\&\N__16928\&\N__17060\&\N__16184\&\N__16328\&\N__17378\;
    \this_vram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18175\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18849\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_3\ <= \this_vram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_2\ <= \this_vram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_1_physical_RADDR_wire\ <= \N__12389\&\N__12233\&\N__12053\&\N__12569\&\N__11654\&\N__13877\&\N__9896\&\N__8120\&\N__10292\&\N__10484\&\N__10706\;
    \this_vram.mem_mem_6_1_physical_WADDR_wire\ <= \N__17222\&\N__16523\&\N__17564\&\N__16655\&\N__17801\&\N__16790\&\N__16922\&\N__17054\&\N__16178\&\N__16322\&\N__17372\;
    \this_vram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19417\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20830\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_1\ <= \this_vram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_0\ <= \this_vram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_0_physical_RADDR_wire\ <= \N__12383\&\N__12227\&\N__12047\&\N__12563\&\N__11648\&\N__13871\&\N__9890\&\N__8114\&\N__10286\&\N__10478\&\N__10700\;
    \this_vram.mem_mem_7_0_physical_WADDR_wire\ <= \N__17216\&\N__16517\&\N__17558\&\N__16649\&\N__17795\&\N__16784\&\N__16916\&\N__17048\&\N__16172\&\N__16316\&\N__17366\;
    \this_vram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18176\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18865\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_3\ <= \this_vram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_2\ <= \this_vram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_1_physical_RADDR_wire\ <= \N__12377\&\N__12221\&\N__12041\&\N__12557\&\N__11642\&\N__13865\&\N__9884\&\N__8108\&\N__10280\&\N__10472\&\N__10694\;
    \this_vram.mem_mem_7_1_physical_WADDR_wire\ <= \N__17210\&\N__16511\&\N__17552\&\N__16643\&\N__17789\&\N__16778\&\N__16910\&\N__17042\&\N__16166\&\N__16310\&\N__17360\;
    \this_vram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19430\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20843\&'0'&'0'&'0';

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21570\,
            RE => \N__20438\,
            WCLKE => \N__18574\,
            WCLK => \N__21571\,
            WE => \N__20436\
        );

    \this_vram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21572\,
            RE => \N__20437\,
            WCLKE => \N__18575\,
            WCLK => \N__21573\,
            WE => \N__20435\
        );

    \this_vram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21574\,
            RE => \N__20420\,
            WCLKE => \N__18650\,
            WCLK => \N__21575\,
            WE => \N__20427\
        );

    \this_vram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21576\,
            RE => \N__20419\,
            WCLKE => \N__18646\,
            WCLK => \N__21577\,
            WE => \N__20434\
        );

    \this_vram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21581\,
            RE => \N__20394\,
            WCLKE => \N__18623\,
            WCLK => \N__21580\,
            WE => \N__20415\
        );

    \this_vram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21585\,
            RE => \N__20393\,
            WCLKE => \N__18622\,
            WCLK => \N__21586\,
            WE => \N__20414\
        );

    \this_vram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21593\,
            RE => \N__20362\,
            WCLKE => \N__18668\,
            WCLK => \N__21594\,
            WE => \N__20382\
        );

    \this_vram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21611\,
            RE => \N__20361\,
            WCLKE => \N__18661\,
            WCLK => \N__21612\,
            WE => \N__20381\
        );

    \this_vram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21621\,
            RE => \N__20324\,
            WCLKE => \N__19087\,
            WCLK => \N__21622\,
            WE => \N__20344\
        );

    \this_vram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21630\,
            RE => \N__20323\,
            WCLKE => \N__19091\,
            WCLK => \N__21631\,
            WE => \N__20343\
        );

    \this_vram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21635\,
            RE => \N__20271\,
            WCLKE => \N__19369\,
            WCLK => \N__21636\,
            WE => \N__20294\
        );

    \this_vram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21640\,
            RE => \N__20188\,
            WCLKE => \N__19370\,
            WCLK => \N__21641\,
            WE => \N__20149\
        );

    \this_vram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21644\,
            RE => \N__20180\,
            WCLKE => \N__20455\,
            WCLK => \N__21645\,
            WE => \N__20207\
        );

    \this_vram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21646\,
            RE => \N__20322\,
            WCLKE => \N__20459\,
            WCLK => \N__21647\,
            WE => \N__20234\
        );

    \this_vram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21649\,
            RE => \N__20305\,
            WCLKE => \N__20782\,
            WCLK => \N__21650\,
            WE => \N__20307\
        );

    \this_vram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21652\,
            RE => \N__20306\,
            WCLKE => \N__20783\,
            WCLK => \N__21653\,
            WE => \N__20308\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__22314\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22316\,
            DIN => \N__22315\,
            DOUT => \N__22314\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22316\,
            PADOUT => \N__22315\,
            PADIN => \N__22314\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22305\,
            DIN => \N__22304\,
            DOUT => \N__22303\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22305\,
            PADOUT => \N__22304\,
            PADIN => \N__22303\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7793\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22296\,
            DIN => \N__22295\,
            DOUT => \N__22294\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22296\,
            PADOUT => \N__22295\,
            PADIN => \N__22294\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11609\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22287\,
            DIN => \N__22286\,
            DOUT => \N__22285\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22287\,
            PADOUT => \N__22286\,
            PADIN => \N__22285\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7937\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22278\,
            DIN => \N__22277\,
            DOUT => \N__22276\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22278\,
            PADOUT => \N__22277\,
            PADIN => \N__22276\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7814\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22269\,
            DIN => \N__22268\,
            DOUT => \N__22267\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22269\,
            PADOUT => \N__22268\,
            PADIN => \N__22267\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__19901\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13580\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22260\,
            DIN => \N__22259\,
            DOUT => \N__22258\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22260\,
            PADOUT => \N__22259\,
            PADIN => \N__22258\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__19877\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13636\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22251\,
            DIN => \N__22250\,
            DOUT => \N__22249\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22251\,
            PADOUT => \N__22250\,
            PADIN => \N__22249\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__19853\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13616\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22242\,
            DIN => \N__22241\,
            DOUT => \N__22240\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22242\,
            PADOUT => \N__22241\,
            PADIN => \N__22240\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__19823\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13640\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22233\,
            DIN => \N__22232\,
            DOUT => \N__22231\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22233\,
            PADOUT => \N__22232\,
            PADIN => \N__22231\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__19799\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13624\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22224\,
            DIN => \N__22223\,
            DOUT => \N__22222\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22224\,
            PADOUT => \N__22223\,
            PADIN => \N__22222\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__21173\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13593\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22215\,
            DIN => \N__22214\,
            DOUT => \N__22213\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22215\,
            PADOUT => \N__22214\,
            PADIN => \N__22213\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__21152\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13623\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22206\,
            DIN => \N__22205\,
            DOUT => \N__22204\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22206\,
            PADOUT => \N__22205\,
            PADIN => \N__22204\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__21131\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13658\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22197\,
            DIN => \N__22196\,
            DOUT => \N__22195\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22197\,
            PADOUT => \N__22196\,
            PADIN => \N__22195\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21050\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13615\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22188\,
            DIN => \N__22187\,
            DOUT => \N__22186\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22188\,
            PADOUT => \N__22187\,
            PADIN => \N__22186\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21020\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13647\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22179\,
            DIN => \N__22178\,
            DOUT => \N__22177\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22179\,
            PADOUT => \N__22178\,
            PADIN => \N__22177\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21002\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13625\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22170\,
            DIN => \N__22169\,
            DOUT => \N__22168\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22170\,
            PADOUT => \N__22169\,
            PADIN => \N__22168\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21908\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13594\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22161\,
            DIN => \N__22160\,
            DOUT => \N__22159\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22161\,
            PADOUT => \N__22160\,
            PADIN => \N__22159\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21884\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13641\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22152\,
            DIN => \N__22151\,
            DOUT => \N__22150\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22152\,
            PADOUT => \N__22151\,
            PADIN => \N__22150\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21677\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13654\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22143\,
            DIN => \N__22142\,
            DOUT => \N__22141\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22143\,
            PADOUT => \N__22142\,
            PADIN => \N__22141\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21104\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13497\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22134\,
            DIN => \N__22133\,
            DOUT => \N__22132\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22134\,
            PADOUT => \N__22133\,
            PADIN => \N__22132\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21071\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13635\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22125\,
            DIN => \N__22124\,
            DOUT => \N__22123\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22125\,
            PADOUT => \N__22124\,
            PADIN => \N__22123\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22116\,
            DIN => \N__22115\,
            DOUT => \N__22114\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22116\,
            PADOUT => \N__22115\,
            PADIN => \N__22114\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22107\,
            DIN => \N__22106\,
            DOUT => \N__22105\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22107\,
            PADOUT => \N__22106\,
            PADIN => \N__22105\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22098\,
            DIN => \N__22097\,
            DOUT => \N__22096\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22098\,
            PADOUT => \N__22097\,
            PADIN => \N__22096\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22089\,
            DIN => \N__22088\,
            DOUT => \N__22087\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22089\,
            PADOUT => \N__22088\,
            PADIN => \N__22087\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22080\,
            DIN => \N__22079\,
            DOUT => \N__22078\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22080\,
            PADOUT => \N__22079\,
            PADIN => \N__22078\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22071\,
            DIN => \N__22070\,
            DOUT => \N__22069\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22071\,
            PADOUT => \N__22070\,
            PADIN => \N__22069\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22062\,
            DIN => \N__22061\,
            DOUT => \N__22060\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22062\,
            PADOUT => \N__22061\,
            PADIN => \N__22060\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22053\,
            DIN => \N__22052\,
            DOUT => \N__22051\,
            PACKAGEPIN => port_data_wire(7)
        );

    \port_data_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22053\,
            PADOUT => \N__22052\,
            PADIN => \N__22051\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22044\,
            DIN => \N__22043\,
            DOUT => \N__22042\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22044\,
            PADOUT => \N__22043\,
            PADIN => \N__22042\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7430\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22035\,
            DIN => \N__22034\,
            DOUT => \N__22033\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22035\,
            PADOUT => \N__22034\,
            PADIN => \N__22033\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14888\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22026\,
            DIN => \N__22025\,
            DOUT => \N__22024\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22026\,
            PADOUT => \N__22025\,
            PADIN => \N__22024\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22017\,
            DIN => \N__22016\,
            DOUT => \N__22015\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22017\,
            PADOUT => \N__22016\,
            PADIN => \N__22015\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7553\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22008\,
            DIN => \N__22007\,
            DOUT => \N__22006\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22008\,
            PADOUT => \N__22007\,
            PADIN => \N__22006\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__20392\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13592\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21999\,
            DIN => \N__21998\,
            DOUT => \N__21997\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21999\,
            PADOUT => \N__21998\,
            PADIN => \N__21997\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7526\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21990\,
            DIN => \N__21989\,
            DOUT => \N__21988\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21990\,
            PADOUT => \N__21989\,
            PADIN => \N__21988\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7493\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21981\,
            DIN => \N__21980\,
            DOUT => \N__21979\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21981\,
            PADOUT => \N__21980\,
            PADIN => \N__21979\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7745\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21972\,
            DIN => \N__21971\,
            DOUT => \N__21970\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21972\,
            PADOUT => \N__21971\,
            PADIN => \N__21970\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7646\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21963\,
            DIN => \N__21962\,
            DOUT => \N__21961\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21963\,
            PADOUT => \N__21962\,
            PADIN => \N__21961\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7616\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21954\,
            DIN => \N__21953\,
            DOUT => \N__21952\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21954\,
            PADOUT => \N__21953\,
            PADIN => \N__21952\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7460\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21945\,
            DIN => \N__21944\,
            DOUT => \N__21943\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__21945\,
            PADOUT => \N__21944\,
            PADIN => \N__21943\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21936\,
            DIN => \N__21935\,
            DOUT => \N__21934\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21936\,
            PADOUT => \N__21935\,
            PADIN => \N__21934\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7577\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21927\,
            DIN => \N__21926\,
            DOUT => \N__21925\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__21927\,
            PADOUT => \N__21926\,
            PADIN => \N__21925\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11750\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__5365\ : IoInMux
    port map (
            O => \N__21908\,
            I => \N__21905\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__21905\,
            I => \N__21902\
        );

    \I__5363\ : IoSpan4Mux
    port map (
            O => \N__21902\,
            I => \N__21899\
        );

    \I__5362\ : Sp12to4
    port map (
            O => \N__21899\,
            I => \N__21895\
        );

    \I__5361\ : InMux
    port map (
            O => \N__21898\,
            I => \N__21892\
        );

    \I__5360\ : Odrv12
    port map (
            O => \N__21895\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__21892\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__5358\ : InMux
    port map (
            O => \N__21887\,
            I => \un1_M_this_external_address_q_cry_12\
        );

    \I__5357\ : IoInMux
    port map (
            O => \N__21884\,
            I => \N__21881\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__21881\,
            I => \N__21878\
        );

    \I__5355\ : Span4Mux_s2_h
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__5354\ : Sp12to4
    port map (
            O => \N__21875\,
            I => \N__21871\
        );

    \I__5353\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21868\
        );

    \I__5352\ : Odrv12
    port map (
            O => \N__21871\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__21868\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__5350\ : InMux
    port map (
            O => \N__21863\,
            I => \un1_M_this_external_address_q_cry_13\
        );

    \I__5349\ : InMux
    port map (
            O => \N__21860\,
            I => \N__21830\
        );

    \I__5348\ : InMux
    port map (
            O => \N__21859\,
            I => \N__21830\
        );

    \I__5347\ : InMux
    port map (
            O => \N__21858\,
            I => \N__21821\
        );

    \I__5346\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21821\
        );

    \I__5345\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21821\
        );

    \I__5344\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21821\
        );

    \I__5343\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21810\
        );

    \I__5342\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21810\
        );

    \I__5341\ : InMux
    port map (
            O => \N__21852\,
            I => \N__21810\
        );

    \I__5340\ : InMux
    port map (
            O => \N__21851\,
            I => \N__21810\
        );

    \I__5339\ : InMux
    port map (
            O => \N__21850\,
            I => \N__21801\
        );

    \I__5338\ : InMux
    port map (
            O => \N__21849\,
            I => \N__21801\
        );

    \I__5337\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21801\
        );

    \I__5336\ : InMux
    port map (
            O => \N__21847\,
            I => \N__21801\
        );

    \I__5335\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21792\
        );

    \I__5334\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21792\
        );

    \I__5333\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21792\
        );

    \I__5332\ : InMux
    port map (
            O => \N__21843\,
            I => \N__21792\
        );

    \I__5331\ : InMux
    port map (
            O => \N__21842\,
            I => \N__21783\
        );

    \I__5330\ : InMux
    port map (
            O => \N__21841\,
            I => \N__21783\
        );

    \I__5329\ : InMux
    port map (
            O => \N__21840\,
            I => \N__21783\
        );

    \I__5328\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21783\
        );

    \I__5327\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21775\
        );

    \I__5326\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21775\
        );

    \I__5325\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21775\
        );

    \I__5324\ : InMux
    port map (
            O => \N__21835\,
            I => \N__21772\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__21830\,
            I => \N__21767\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__21821\,
            I => \N__21767\
        );

    \I__5321\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21762\
        );

    \I__5320\ : InMux
    port map (
            O => \N__21819\,
            I => \N__21762\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__21810\,
            I => \N__21758\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__21801\,
            I => \N__21751\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__21792\,
            I => \N__21751\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__21783\,
            I => \N__21751\
        );

    \I__5315\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21748\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__21775\,
            I => \N__21743\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__21772\,
            I => \N__21736\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__21767\,
            I => \N__21736\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__21762\,
            I => \N__21736\
        );

    \I__5310\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21733\
        );

    \I__5309\ : Span4Mux_v
    port map (
            O => \N__21758\,
            I => \N__21728\
        );

    \I__5308\ : Span4Mux_v
    port map (
            O => \N__21751\,
            I => \N__21728\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__21748\,
            I => \N__21724\
        );

    \I__5306\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21719\
        );

    \I__5305\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21719\
        );

    \I__5304\ : Span4Mux_v
    port map (
            O => \N__21743\,
            I => \N__21714\
        );

    \I__5303\ : Span4Mux_v
    port map (
            O => \N__21736\,
            I => \N__21711\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__21733\,
            I => \N__21706\
        );

    \I__5301\ : Sp12to4
    port map (
            O => \N__21728\,
            I => \N__21706\
        );

    \I__5300\ : InMux
    port map (
            O => \N__21727\,
            I => \N__21703\
        );

    \I__5299\ : Span4Mux_h
    port map (
            O => \N__21724\,
            I => \N__21698\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__21719\,
            I => \N__21698\
        );

    \I__5297\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21693\
        );

    \I__5296\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21693\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__21714\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__21711\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__5293\ : Odrv12
    port map (
            O => \N__21706\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__21703\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__5291\ : Odrv4
    port map (
            O => \N__21698\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__21693\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__5289\ : InMux
    port map (
            O => \N__21680\,
            I => \un1_M_this_external_address_q_cry_14\
        );

    \I__5288\ : IoInMux
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__5286\ : Span4Mux_s2_h
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__5285\ : Sp12to4
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__5284\ : Span12Mux_v
    port map (
            O => \N__21665\,
            I => \N__21661\
        );

    \I__5283\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21658\
        );

    \I__5282\ : Odrv12
    port map (
            O => \N__21661\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__21658\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__5280\ : ClkMux
    port map (
            O => \N__21653\,
            I => \N__21401\
        );

    \I__5279\ : ClkMux
    port map (
            O => \N__21652\,
            I => \N__21401\
        );

    \I__5278\ : ClkMux
    port map (
            O => \N__21651\,
            I => \N__21401\
        );

    \I__5277\ : ClkMux
    port map (
            O => \N__21650\,
            I => \N__21401\
        );

    \I__5276\ : ClkMux
    port map (
            O => \N__21649\,
            I => \N__21401\
        );

    \I__5275\ : ClkMux
    port map (
            O => \N__21648\,
            I => \N__21401\
        );

    \I__5274\ : ClkMux
    port map (
            O => \N__21647\,
            I => \N__21401\
        );

    \I__5273\ : ClkMux
    port map (
            O => \N__21646\,
            I => \N__21401\
        );

    \I__5272\ : ClkMux
    port map (
            O => \N__21645\,
            I => \N__21401\
        );

    \I__5271\ : ClkMux
    port map (
            O => \N__21644\,
            I => \N__21401\
        );

    \I__5270\ : ClkMux
    port map (
            O => \N__21643\,
            I => \N__21401\
        );

    \I__5269\ : ClkMux
    port map (
            O => \N__21642\,
            I => \N__21401\
        );

    \I__5268\ : ClkMux
    port map (
            O => \N__21641\,
            I => \N__21401\
        );

    \I__5267\ : ClkMux
    port map (
            O => \N__21640\,
            I => \N__21401\
        );

    \I__5266\ : ClkMux
    port map (
            O => \N__21639\,
            I => \N__21401\
        );

    \I__5265\ : ClkMux
    port map (
            O => \N__21638\,
            I => \N__21401\
        );

    \I__5264\ : ClkMux
    port map (
            O => \N__21637\,
            I => \N__21401\
        );

    \I__5263\ : ClkMux
    port map (
            O => \N__21636\,
            I => \N__21401\
        );

    \I__5262\ : ClkMux
    port map (
            O => \N__21635\,
            I => \N__21401\
        );

    \I__5261\ : ClkMux
    port map (
            O => \N__21634\,
            I => \N__21401\
        );

    \I__5260\ : ClkMux
    port map (
            O => \N__21633\,
            I => \N__21401\
        );

    \I__5259\ : ClkMux
    port map (
            O => \N__21632\,
            I => \N__21401\
        );

    \I__5258\ : ClkMux
    port map (
            O => \N__21631\,
            I => \N__21401\
        );

    \I__5257\ : ClkMux
    port map (
            O => \N__21630\,
            I => \N__21401\
        );

    \I__5256\ : ClkMux
    port map (
            O => \N__21629\,
            I => \N__21401\
        );

    \I__5255\ : ClkMux
    port map (
            O => \N__21628\,
            I => \N__21401\
        );

    \I__5254\ : ClkMux
    port map (
            O => \N__21627\,
            I => \N__21401\
        );

    \I__5253\ : ClkMux
    port map (
            O => \N__21626\,
            I => \N__21401\
        );

    \I__5252\ : ClkMux
    port map (
            O => \N__21625\,
            I => \N__21401\
        );

    \I__5251\ : ClkMux
    port map (
            O => \N__21624\,
            I => \N__21401\
        );

    \I__5250\ : ClkMux
    port map (
            O => \N__21623\,
            I => \N__21401\
        );

    \I__5249\ : ClkMux
    port map (
            O => \N__21622\,
            I => \N__21401\
        );

    \I__5248\ : ClkMux
    port map (
            O => \N__21621\,
            I => \N__21401\
        );

    \I__5247\ : ClkMux
    port map (
            O => \N__21620\,
            I => \N__21401\
        );

    \I__5246\ : ClkMux
    port map (
            O => \N__21619\,
            I => \N__21401\
        );

    \I__5245\ : ClkMux
    port map (
            O => \N__21618\,
            I => \N__21401\
        );

    \I__5244\ : ClkMux
    port map (
            O => \N__21617\,
            I => \N__21401\
        );

    \I__5243\ : ClkMux
    port map (
            O => \N__21616\,
            I => \N__21401\
        );

    \I__5242\ : ClkMux
    port map (
            O => \N__21615\,
            I => \N__21401\
        );

    \I__5241\ : ClkMux
    port map (
            O => \N__21614\,
            I => \N__21401\
        );

    \I__5240\ : ClkMux
    port map (
            O => \N__21613\,
            I => \N__21401\
        );

    \I__5239\ : ClkMux
    port map (
            O => \N__21612\,
            I => \N__21401\
        );

    \I__5238\ : ClkMux
    port map (
            O => \N__21611\,
            I => \N__21401\
        );

    \I__5237\ : ClkMux
    port map (
            O => \N__21610\,
            I => \N__21401\
        );

    \I__5236\ : ClkMux
    port map (
            O => \N__21609\,
            I => \N__21401\
        );

    \I__5235\ : ClkMux
    port map (
            O => \N__21608\,
            I => \N__21401\
        );

    \I__5234\ : ClkMux
    port map (
            O => \N__21607\,
            I => \N__21401\
        );

    \I__5233\ : ClkMux
    port map (
            O => \N__21606\,
            I => \N__21401\
        );

    \I__5232\ : ClkMux
    port map (
            O => \N__21605\,
            I => \N__21401\
        );

    \I__5231\ : ClkMux
    port map (
            O => \N__21604\,
            I => \N__21401\
        );

    \I__5230\ : ClkMux
    port map (
            O => \N__21603\,
            I => \N__21401\
        );

    \I__5229\ : ClkMux
    port map (
            O => \N__21602\,
            I => \N__21401\
        );

    \I__5228\ : ClkMux
    port map (
            O => \N__21601\,
            I => \N__21401\
        );

    \I__5227\ : ClkMux
    port map (
            O => \N__21600\,
            I => \N__21401\
        );

    \I__5226\ : ClkMux
    port map (
            O => \N__21599\,
            I => \N__21401\
        );

    \I__5225\ : ClkMux
    port map (
            O => \N__21598\,
            I => \N__21401\
        );

    \I__5224\ : ClkMux
    port map (
            O => \N__21597\,
            I => \N__21401\
        );

    \I__5223\ : ClkMux
    port map (
            O => \N__21596\,
            I => \N__21401\
        );

    \I__5222\ : ClkMux
    port map (
            O => \N__21595\,
            I => \N__21401\
        );

    \I__5221\ : ClkMux
    port map (
            O => \N__21594\,
            I => \N__21401\
        );

    \I__5220\ : ClkMux
    port map (
            O => \N__21593\,
            I => \N__21401\
        );

    \I__5219\ : ClkMux
    port map (
            O => \N__21592\,
            I => \N__21401\
        );

    \I__5218\ : ClkMux
    port map (
            O => \N__21591\,
            I => \N__21401\
        );

    \I__5217\ : ClkMux
    port map (
            O => \N__21590\,
            I => \N__21401\
        );

    \I__5216\ : ClkMux
    port map (
            O => \N__21589\,
            I => \N__21401\
        );

    \I__5215\ : ClkMux
    port map (
            O => \N__21588\,
            I => \N__21401\
        );

    \I__5214\ : ClkMux
    port map (
            O => \N__21587\,
            I => \N__21401\
        );

    \I__5213\ : ClkMux
    port map (
            O => \N__21586\,
            I => \N__21401\
        );

    \I__5212\ : ClkMux
    port map (
            O => \N__21585\,
            I => \N__21401\
        );

    \I__5211\ : ClkMux
    port map (
            O => \N__21584\,
            I => \N__21401\
        );

    \I__5210\ : ClkMux
    port map (
            O => \N__21583\,
            I => \N__21401\
        );

    \I__5209\ : ClkMux
    port map (
            O => \N__21582\,
            I => \N__21401\
        );

    \I__5208\ : ClkMux
    port map (
            O => \N__21581\,
            I => \N__21401\
        );

    \I__5207\ : ClkMux
    port map (
            O => \N__21580\,
            I => \N__21401\
        );

    \I__5206\ : ClkMux
    port map (
            O => \N__21579\,
            I => \N__21401\
        );

    \I__5205\ : ClkMux
    port map (
            O => \N__21578\,
            I => \N__21401\
        );

    \I__5204\ : ClkMux
    port map (
            O => \N__21577\,
            I => \N__21401\
        );

    \I__5203\ : ClkMux
    port map (
            O => \N__21576\,
            I => \N__21401\
        );

    \I__5202\ : ClkMux
    port map (
            O => \N__21575\,
            I => \N__21401\
        );

    \I__5201\ : ClkMux
    port map (
            O => \N__21574\,
            I => \N__21401\
        );

    \I__5200\ : ClkMux
    port map (
            O => \N__21573\,
            I => \N__21401\
        );

    \I__5199\ : ClkMux
    port map (
            O => \N__21572\,
            I => \N__21401\
        );

    \I__5198\ : ClkMux
    port map (
            O => \N__21571\,
            I => \N__21401\
        );

    \I__5197\ : ClkMux
    port map (
            O => \N__21570\,
            I => \N__21401\
        );

    \I__5196\ : GlobalMux
    port map (
            O => \N__21401\,
            I => \N__21398\
        );

    \I__5195\ : gio2CtrlBuf
    port map (
            O => \N__21398\,
            I => clk_0_c_g
        );

    \I__5194\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21381\
        );

    \I__5193\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21378\
        );

    \I__5192\ : InMux
    port map (
            O => \N__21393\,
            I => \N__21375\
        );

    \I__5191\ : InMux
    port map (
            O => \N__21392\,
            I => \N__21372\
        );

    \I__5190\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21369\
        );

    \I__5189\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21366\
        );

    \I__5188\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21359\
        );

    \I__5187\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21359\
        );

    \I__5186\ : InMux
    port map (
            O => \N__21387\,
            I => \N__21359\
        );

    \I__5185\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21354\
        );

    \I__5184\ : InMux
    port map (
            O => \N__21385\,
            I => \N__21354\
        );

    \I__5183\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21351\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__21381\,
            I => \N__21337\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__21378\,
            I => \N__21334\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__21375\,
            I => \N__21331\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__21372\,
            I => \N__21328\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__21369\,
            I => \N__21325\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__21366\,
            I => \N__21322\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__21359\,
            I => \N__21319\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__21354\,
            I => \N__21316\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__21351\,
            I => \N__21313\
        );

    \I__5173\ : SRMux
    port map (
            O => \N__21350\,
            I => \N__21272\
        );

    \I__5172\ : SRMux
    port map (
            O => \N__21349\,
            I => \N__21272\
        );

    \I__5171\ : SRMux
    port map (
            O => \N__21348\,
            I => \N__21272\
        );

    \I__5170\ : SRMux
    port map (
            O => \N__21347\,
            I => \N__21272\
        );

    \I__5169\ : SRMux
    port map (
            O => \N__21346\,
            I => \N__21272\
        );

    \I__5168\ : SRMux
    port map (
            O => \N__21345\,
            I => \N__21272\
        );

    \I__5167\ : SRMux
    port map (
            O => \N__21344\,
            I => \N__21272\
        );

    \I__5166\ : SRMux
    port map (
            O => \N__21343\,
            I => \N__21272\
        );

    \I__5165\ : SRMux
    port map (
            O => \N__21342\,
            I => \N__21272\
        );

    \I__5164\ : SRMux
    port map (
            O => \N__21341\,
            I => \N__21272\
        );

    \I__5163\ : SRMux
    port map (
            O => \N__21340\,
            I => \N__21272\
        );

    \I__5162\ : Glb2LocalMux
    port map (
            O => \N__21337\,
            I => \N__21272\
        );

    \I__5161\ : Glb2LocalMux
    port map (
            O => \N__21334\,
            I => \N__21272\
        );

    \I__5160\ : Glb2LocalMux
    port map (
            O => \N__21331\,
            I => \N__21272\
        );

    \I__5159\ : Glb2LocalMux
    port map (
            O => \N__21328\,
            I => \N__21272\
        );

    \I__5158\ : Glb2LocalMux
    port map (
            O => \N__21325\,
            I => \N__21272\
        );

    \I__5157\ : Glb2LocalMux
    port map (
            O => \N__21322\,
            I => \N__21272\
        );

    \I__5156\ : Glb2LocalMux
    port map (
            O => \N__21319\,
            I => \N__21272\
        );

    \I__5155\ : Glb2LocalMux
    port map (
            O => \N__21316\,
            I => \N__21272\
        );

    \I__5154\ : Glb2LocalMux
    port map (
            O => \N__21313\,
            I => \N__21272\
        );

    \I__5153\ : GlobalMux
    port map (
            O => \N__21272\,
            I => \N__21269\
        );

    \I__5152\ : gio2CtrlBuf
    port map (
            O => \N__21269\,
            I => \M_this_state_q_nss_g_0\
        );

    \I__5151\ : InMux
    port map (
            O => \N__21266\,
            I => \N__21263\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__5149\ : Span4Mux_v
    port map (
            O => \N__21260\,
            I => \N__21257\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__21257\,
            I => port_address_in_5
        );

    \I__5147\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__5145\ : Span12Mux_v
    port map (
            O => \N__21248\,
            I => \N__21245\
        );

    \I__5144\ : Odrv12
    port map (
            O => \N__21245\,
            I => port_address_in_6
        );

    \I__5143\ : CascadeMux
    port map (
            O => \N__21242\,
            I => \N__21239\
        );

    \I__5142\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21236\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__21236\,
            I => \N__21233\
        );

    \I__5140\ : Span4Mux_v
    port map (
            O => \N__21233\,
            I => \N__21230\
        );

    \I__5139\ : Span4Mux_v
    port map (
            O => \N__21230\,
            I => \N__21227\
        );

    \I__5138\ : Span4Mux_v
    port map (
            O => \N__21227\,
            I => \N__21224\
        );

    \I__5137\ : Span4Mux_v
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__5136\ : Odrv4
    port map (
            O => \N__21221\,
            I => port_address_in_7
        );

    \I__5135\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21212\
        );

    \I__5133\ : IoSpan4Mux
    port map (
            O => \N__21212\,
            I => \N__21209\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__21209\,
            I => port_address_in_4
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__21206\,
            I => \N__21202\
        );

    \I__5130\ : CascadeMux
    port map (
            O => \N__21205\,
            I => \N__21198\
        );

    \I__5129\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21188\
        );

    \I__5128\ : InMux
    port map (
            O => \N__21201\,
            I => \N__21188\
        );

    \I__5127\ : InMux
    port map (
            O => \N__21198\,
            I => \N__21188\
        );

    \I__5126\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21188\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__21188\,
            I => \N__21185\
        );

    \I__5124\ : Span12Mux_v
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__5123\ : Span12Mux_h
    port map (
            O => \N__21182\,
            I => \N__21179\
        );

    \I__5122\ : Odrv12
    port map (
            O => \N__21179\,
            I => \this_start_data_delay.M_this_state_d27Z0Z_6\
        );

    \I__5121\ : InMux
    port map (
            O => \N__21176\,
            I => \un1_M_this_external_address_q_cry_3\
        );

    \I__5120\ : IoInMux
    port map (
            O => \N__21173\,
            I => \N__21170\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__21170\,
            I => \N__21167\
        );

    \I__5118\ : Span4Mux_s2_h
    port map (
            O => \N__21167\,
            I => \N__21163\
        );

    \I__5117\ : InMux
    port map (
            O => \N__21166\,
            I => \N__21160\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__21163\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__21160\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__5114\ : InMux
    port map (
            O => \N__21155\,
            I => \un1_M_this_external_address_q_cry_4\
        );

    \I__5113\ : IoInMux
    port map (
            O => \N__21152\,
            I => \N__21149\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__21149\,
            I => \N__21146\
        );

    \I__5111\ : Span12Mux_s2_h
    port map (
            O => \N__21146\,
            I => \N__21142\
        );

    \I__5110\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21139\
        );

    \I__5109\ : Odrv12
    port map (
            O => \N__21142\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__21139\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__5107\ : InMux
    port map (
            O => \N__21134\,
            I => \un1_M_this_external_address_q_cry_5\
        );

    \I__5106\ : IoInMux
    port map (
            O => \N__21131\,
            I => \N__21128\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__21128\,
            I => \N__21125\
        );

    \I__5104\ : Span4Mux_s2_h
    port map (
            O => \N__21125\,
            I => \N__21122\
        );

    \I__5103\ : Sp12to4
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__5102\ : Span12Mux_v
    port map (
            O => \N__21119\,
            I => \N__21115\
        );

    \I__5101\ : InMux
    port map (
            O => \N__21118\,
            I => \N__21112\
        );

    \I__5100\ : Odrv12
    port map (
            O => \N__21115\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__21112\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__5098\ : InMux
    port map (
            O => \N__21107\,
            I => \un1_M_this_external_address_q_cry_6\
        );

    \I__5097\ : IoInMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__5095\ : IoSpan4Mux
    port map (
            O => \N__21098\,
            I => \N__21095\
        );

    \I__5094\ : Span4Mux_s2_v
    port map (
            O => \N__21095\,
            I => \N__21092\
        );

    \I__5093\ : Sp12to4
    port map (
            O => \N__21092\,
            I => \N__21089\
        );

    \I__5092\ : Span12Mux_s8_v
    port map (
            O => \N__21089\,
            I => \N__21086\
        );

    \I__5091\ : Span12Mux_h
    port map (
            O => \N__21086\,
            I => \N__21082\
        );

    \I__5090\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21079\
        );

    \I__5089\ : Odrv12
    port map (
            O => \N__21082\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__21079\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__5087\ : InMux
    port map (
            O => \N__21074\,
            I => \bfn_30_24_0_\
        );

    \I__5086\ : IoInMux
    port map (
            O => \N__21071\,
            I => \N__21068\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__21068\,
            I => \N__21065\
        );

    \I__5084\ : Span12Mux_s8_v
    port map (
            O => \N__21065\,
            I => \N__21061\
        );

    \I__5083\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21058\
        );

    \I__5082\ : Odrv12
    port map (
            O => \N__21061\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__21058\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__5080\ : InMux
    port map (
            O => \N__21053\,
            I => \un1_M_this_external_address_q_cry_8\
        );

    \I__5079\ : IoInMux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__21047\,
            I => \N__21044\
        );

    \I__5077\ : Span4Mux_s2_v
    port map (
            O => \N__21044\,
            I => \N__21041\
        );

    \I__5076\ : Span4Mux_h
    port map (
            O => \N__21041\,
            I => \N__21038\
        );

    \I__5075\ : Sp12to4
    port map (
            O => \N__21038\,
            I => \N__21035\
        );

    \I__5074\ : Span12Mux_s8_v
    port map (
            O => \N__21035\,
            I => \N__21031\
        );

    \I__5073\ : InMux
    port map (
            O => \N__21034\,
            I => \N__21028\
        );

    \I__5072\ : Odrv12
    port map (
            O => \N__21031\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__21028\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__5070\ : InMux
    port map (
            O => \N__21023\,
            I => \un1_M_this_external_address_q_cry_9\
        );

    \I__5069\ : IoInMux
    port map (
            O => \N__21020\,
            I => \N__21017\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__21017\,
            I => \N__21013\
        );

    \I__5067\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21010\
        );

    \I__5066\ : Odrv12
    port map (
            O => \N__21013\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__21010\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__5064\ : InMux
    port map (
            O => \N__21005\,
            I => \un1_M_this_external_address_q_cry_10\
        );

    \I__5063\ : IoInMux
    port map (
            O => \N__21002\,
            I => \N__20999\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20995\
        );

    \I__5061\ : InMux
    port map (
            O => \N__20998\,
            I => \N__20992\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__20995\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__20992\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__5058\ : InMux
    port map (
            O => \N__20987\,
            I => \un1_M_this_external_address_q_cry_11\
        );

    \I__5057\ : CascadeMux
    port map (
            O => \N__20984\,
            I => \N__20981\
        );

    \I__5056\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20978\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__20978\,
            I => \N__20974\
        );

    \I__5054\ : CascadeMux
    port map (
            O => \N__20977\,
            I => \N__20971\
        );

    \I__5053\ : Span4Mux_h
    port map (
            O => \N__20974\,
            I => \N__20967\
        );

    \I__5052\ : InMux
    port map (
            O => \N__20971\,
            I => \N__20964\
        );

    \I__5051\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20961\
        );

    \I__5050\ : Span4Mux_h
    port map (
            O => \N__20967\,
            I => \N__20958\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__20964\,
            I => \N__20953\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__20961\,
            I => \N__20953\
        );

    \I__5047\ : Sp12to4
    port map (
            O => \N__20958\,
            I => \N__20950\
        );

    \I__5046\ : Span12Mux_h
    port map (
            O => \N__20953\,
            I => \N__20947\
        );

    \I__5045\ : Odrv12
    port map (
            O => \N__20950\,
            I => port_data_c_2
        );

    \I__5044\ : Odrv12
    port map (
            O => \N__20947\,
            I => port_data_c_2
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__20942\,
            I => \N__20939\
        );

    \I__5042\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20935\
        );

    \I__5041\ : CascadeMux
    port map (
            O => \N__20938\,
            I => \N__20932\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__20935\,
            I => \N__20929\
        );

    \I__5039\ : InMux
    port map (
            O => \N__20932\,
            I => \N__20926\
        );

    \I__5038\ : Span4Mux_h
    port map (
            O => \N__20929\,
            I => \N__20921\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__20926\,
            I => \N__20921\
        );

    \I__5036\ : Span4Mux_h
    port map (
            O => \N__20921\,
            I => \N__20917\
        );

    \I__5035\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20914\
        );

    \I__5034\ : Sp12to4
    port map (
            O => \N__20917\,
            I => \N__20909\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__20914\,
            I => \N__20909\
        );

    \I__5032\ : Span12Mux_v
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__5031\ : Odrv12
    port map (
            O => \N__20906\,
            I => port_data_c_6
        );

    \I__5030\ : CascadeMux
    port map (
            O => \N__20903\,
            I => \N__20898\
        );

    \I__5029\ : InMux
    port map (
            O => \N__20902\,
            I => \N__20895\
        );

    \I__5028\ : InMux
    port map (
            O => \N__20901\,
            I => \N__20892\
        );

    \I__5027\ : InMux
    port map (
            O => \N__20898\,
            I => \N__20889\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__20895\,
            I => \N__20886\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__20892\,
            I => \M_this_vram_write_data_0_sqmuxa\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__20889\,
            I => \M_this_vram_write_data_0_sqmuxa\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__20886\,
            I => \M_this_vram_write_data_0_sqmuxa\
        );

    \I__5022\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20873\
        );

    \I__5021\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20870\
        );

    \I__5020\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20867\
        );

    \I__5019\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20864\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__20873\,
            I => \this_start_data_delay.un1_M_this_state_q_0\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__20870\,
            I => \this_start_data_delay.un1_M_this_state_q_0\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__20867\,
            I => \this_start_data_delay.un1_M_this_state_q_0\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__20864\,
            I => \this_start_data_delay.un1_M_this_state_q_0\
        );

    \I__5014\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20852\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__20852\,
            I => \N__20848\
        );

    \I__5012\ : InMux
    port map (
            O => \N__20851\,
            I => \N__20845\
        );

    \I__5011\ : Span4Mux_v
    port map (
            O => \N__20848\,
            I => \N__20838\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__20845\,
            I => \N__20838\
        );

    \I__5009\ : InMux
    port map (
            O => \N__20844\,
            I => \N__20835\
        );

    \I__5008\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20831\
        );

    \I__5007\ : Span4Mux_v
    port map (
            O => \N__20838\,
            I => \N__20825\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__20835\,
            I => \N__20825\
        );

    \I__5005\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20822\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__20831\,
            I => \N__20819\
        );

    \I__5003\ : InMux
    port map (
            O => \N__20830\,
            I => \N__20816\
        );

    \I__5002\ : Span4Mux_v
    port map (
            O => \N__20825\,
            I => \N__20810\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__20822\,
            I => \N__20810\
        );

    \I__5000\ : Span4Mux_v
    port map (
            O => \N__20819\,
            I => \N__20805\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__20816\,
            I => \N__20805\
        );

    \I__4998\ : InMux
    port map (
            O => \N__20815\,
            I => \N__20802\
        );

    \I__4997\ : Span4Mux_v
    port map (
            O => \N__20810\,
            I => \N__20798\
        );

    \I__4996\ : Span4Mux_v
    port map (
            O => \N__20805\,
            I => \N__20793\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__20802\,
            I => \N__20793\
        );

    \I__4994\ : InMux
    port map (
            O => \N__20801\,
            I => \N__20790\
        );

    \I__4993\ : Odrv4
    port map (
            O => \N__20798\,
            I => \M_this_vram_write_data_0_i_2\
        );

    \I__4992\ : Odrv4
    port map (
            O => \N__20793\,
            I => \M_this_vram_write_data_0_i_2\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__20790\,
            I => \M_this_vram_write_data_0_i_2\
        );

    \I__4990\ : CEMux
    port map (
            O => \N__20783\,
            I => \N__20779\
        );

    \I__4989\ : CEMux
    port map (
            O => \N__20782\,
            I => \N__20776\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__20779\,
            I => \N__20771\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__20776\,
            I => \N__20771\
        );

    \I__4986\ : Span4Mux_s3_v
    port map (
            O => \N__20771\,
            I => \N__20768\
        );

    \I__4985\ : Span4Mux_v
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__20765\,
            I => \this_vram.mem_WE_0\
        );

    \I__4983\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20752\
        );

    \I__4982\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20752\
        );

    \I__4981\ : InMux
    port map (
            O => \N__20760\,
            I => \N__20752\
        );

    \I__4980\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20746\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__20752\,
            I => \N__20743\
        );

    \I__4978\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20740\
        );

    \I__4977\ : InMux
    port map (
            O => \N__20750\,
            I => \N__20735\
        );

    \I__4976\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20735\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__20746\,
            I => \N__20731\
        );

    \I__4974\ : Span4Mux_v
    port map (
            O => \N__20743\,
            I => \N__20725\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__20740\,
            I => \N__20725\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__20735\,
            I => \N__20722\
        );

    \I__4971\ : InMux
    port map (
            O => \N__20734\,
            I => \N__20719\
        );

    \I__4970\ : Span4Mux_v
    port map (
            O => \N__20731\,
            I => \N__20716\
        );

    \I__4969\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20713\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__20725\,
            I => \N__20707\
        );

    \I__4967\ : Span4Mux_h
    port map (
            O => \N__20722\,
            I => \N__20707\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__20719\,
            I => \N__20704\
        );

    \I__4965\ : Span4Mux_v
    port map (
            O => \N__20716\,
            I => \N__20699\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__20713\,
            I => \N__20699\
        );

    \I__4963\ : InMux
    port map (
            O => \N__20712\,
            I => \N__20696\
        );

    \I__4962\ : Odrv4
    port map (
            O => \N__20707\,
            I => \M_this_internal_address_qZ0Z_12\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__20704\,
            I => \M_this_internal_address_qZ0Z_12\
        );

    \I__4960\ : Odrv4
    port map (
            O => \N__20699\,
            I => \M_this_internal_address_qZ0Z_12\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__20696\,
            I => \M_this_internal_address_qZ0Z_12\
        );

    \I__4958\ : CascadeMux
    port map (
            O => \N__20687\,
            I => \N__20682\
        );

    \I__4957\ : CascadeMux
    port map (
            O => \N__20686\,
            I => \N__20676\
        );

    \I__4956\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20672\
        );

    \I__4955\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20665\
        );

    \I__4954\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20665\
        );

    \I__4953\ : InMux
    port map (
            O => \N__20680\,
            I => \N__20665\
        );

    \I__4952\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20660\
        );

    \I__4951\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20655\
        );

    \I__4950\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20655\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__20672\,
            I => \N__20650\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__20665\,
            I => \N__20650\
        );

    \I__4947\ : CascadeMux
    port map (
            O => \N__20664\,
            I => \N__20647\
        );

    \I__4946\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20644\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__20660\,
            I => \N__20641\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__20655\,
            I => \N__20638\
        );

    \I__4943\ : Span4Mux_h
    port map (
            O => \N__20650\,
            I => \N__20635\
        );

    \I__4942\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20631\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__20644\,
            I => \N__20628\
        );

    \I__4940\ : Span4Mux_v
    port map (
            O => \N__20641\,
            I => \N__20623\
        );

    \I__4939\ : Span4Mux_v
    port map (
            O => \N__20638\,
            I => \N__20623\
        );

    \I__4938\ : Span4Mux_v
    port map (
            O => \N__20635\,
            I => \N__20620\
        );

    \I__4937\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20617\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__20631\,
            I => \N__20614\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__20628\,
            I => \N__20609\
        );

    \I__4934\ : Span4Mux_h
    port map (
            O => \N__20623\,
            I => \N__20609\
        );

    \I__4933\ : Span4Mux_h
    port map (
            O => \N__20620\,
            I => \N__20606\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__20617\,
            I => \M_this_internal_address_qZ0Z_11\
        );

    \I__4931\ : Odrv12
    port map (
            O => \N__20614\,
            I => \M_this_internal_address_qZ0Z_11\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__20609\,
            I => \M_this_internal_address_qZ0Z_11\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__20606\,
            I => \M_this_internal_address_qZ0Z_11\
        );

    \I__4928\ : CascadeMux
    port map (
            O => \N__20597\,
            I => \N__20591\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__20596\,
            I => \N__20587\
        );

    \I__4926\ : CascadeMux
    port map (
            O => \N__20595\,
            I => \N__20584\
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__20594\,
            I => \N__20581\
        );

    \I__4924\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20574\
        );

    \I__4923\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20574\
        );

    \I__4922\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20574\
        );

    \I__4921\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20571\
        );

    \I__4920\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20568\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20561\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__20571\,
            I => \N__20561\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__20568\,
            I => \N__20558\
        );

    \I__4916\ : InMux
    port map (
            O => \N__20567\,
            I => \N__20555\
        );

    \I__4915\ : CascadeMux
    port map (
            O => \N__20566\,
            I => \N__20551\
        );

    \I__4914\ : Span4Mux_v
    port map (
            O => \N__20561\,
            I => \N__20543\
        );

    \I__4913\ : Span4Mux_h
    port map (
            O => \N__20558\,
            I => \N__20543\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__20555\,
            I => \N__20543\
        );

    \I__4911\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20538\
        );

    \I__4910\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20538\
        );

    \I__4909\ : InMux
    port map (
            O => \N__20550\,
            I => \N__20535\
        );

    \I__4908\ : Span4Mux_v
    port map (
            O => \N__20543\,
            I => \N__20530\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__20538\,
            I => \N__20530\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__20535\,
            I => \N__20527\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__20530\,
            I => \N__20521\
        );

    \I__4904\ : Span4Mux_v
    port map (
            O => \N__20527\,
            I => \N__20521\
        );

    \I__4903\ : InMux
    port map (
            O => \N__20526\,
            I => \N__20518\
        );

    \I__4902\ : Odrv4
    port map (
            O => \N__20521\,
            I => \M_this_internal_address_qZ0Z_13\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__20518\,
            I => \M_this_internal_address_qZ0Z_13\
        );

    \I__4900\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20503\
        );

    \I__4899\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20503\
        );

    \I__4898\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20503\
        );

    \I__4897\ : InMux
    port map (
            O => \N__20510\,
            I => \N__20499\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__20503\,
            I => \N__20496\
        );

    \I__4895\ : InMux
    port map (
            O => \N__20502\,
            I => \N__20493\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__20499\,
            I => \N__20490\
        );

    \I__4893\ : Span4Mux_v
    port map (
            O => \N__20496\,
            I => \N__20484\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__20493\,
            I => \N__20481\
        );

    \I__4891\ : Span4Mux_h
    port map (
            O => \N__20490\,
            I => \N__20478\
        );

    \I__4890\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20475\
        );

    \I__4889\ : InMux
    port map (
            O => \N__20488\,
            I => \N__20470\
        );

    \I__4888\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20470\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__20484\,
            I => \M_this_vram_write_en_0_0\
        );

    \I__4886\ : Odrv12
    port map (
            O => \N__20481\,
            I => \M_this_vram_write_en_0_0\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__20478\,
            I => \M_this_vram_write_en_0_0\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__20475\,
            I => \M_this_vram_write_en_0_0\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__20470\,
            I => \M_this_vram_write_en_0_0\
        );

    \I__4882\ : CEMux
    port map (
            O => \N__20459\,
            I => \N__20456\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__20456\,
            I => \N__20452\
        );

    \I__4880\ : CEMux
    port map (
            O => \N__20455\,
            I => \N__20449\
        );

    \I__4879\ : Span4Mux_v
    port map (
            O => \N__20452\,
            I => \N__20444\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__20449\,
            I => \N__20444\
        );

    \I__4877\ : Span4Mux_v
    port map (
            O => \N__20444\,
            I => \N__20441\
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__20441\,
            I => \this_vram.mem_WE_2\
        );

    \I__4875\ : SRMux
    port map (
            O => \N__20438\,
            I => \N__20431\
        );

    \I__4874\ : SRMux
    port map (
            O => \N__20437\,
            I => \N__20428\
        );

    \I__4873\ : SRMux
    port map (
            O => \N__20436\,
            I => \N__20424\
        );

    \I__4872\ : SRMux
    port map (
            O => \N__20435\,
            I => \N__20421\
        );

    \I__4871\ : SRMux
    port map (
            O => \N__20434\,
            I => \N__20416\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__20431\,
            I => \N__20409\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__20428\,
            I => \N__20409\
        );

    \I__4868\ : SRMux
    port map (
            O => \N__20427\,
            I => \N__20406\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__20424\,
            I => \N__20401\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__20421\,
            I => \N__20401\
        );

    \I__4865\ : SRMux
    port map (
            O => \N__20420\,
            I => \N__20398\
        );

    \I__4864\ : SRMux
    port map (
            O => \N__20419\,
            I => \N__20395\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__20416\,
            I => \N__20389\
        );

    \I__4862\ : SRMux
    port map (
            O => \N__20415\,
            I => \N__20386\
        );

    \I__4861\ : SRMux
    port map (
            O => \N__20414\,
            I => \N__20383\
        );

    \I__4860\ : Span4Mux_s3_v
    port map (
            O => \N__20409\,
            I => \N__20376\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__20406\,
            I => \N__20376\
        );

    \I__4858\ : Span4Mux_s3_v
    port map (
            O => \N__20401\,
            I => \N__20369\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__20398\,
            I => \N__20369\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__20395\,
            I => \N__20369\
        );

    \I__4855\ : SRMux
    port map (
            O => \N__20394\,
            I => \N__20366\
        );

    \I__4854\ : SRMux
    port map (
            O => \N__20393\,
            I => \N__20363\
        );

    \I__4853\ : IoInMux
    port map (
            O => \N__20392\,
            I => \N__20357\
        );

    \I__4852\ : Span4Mux_h
    port map (
            O => \N__20389\,
            I => \N__20351\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__20386\,
            I => \N__20351\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__20383\,
            I => \N__20348\
        );

    \I__4849\ : SRMux
    port map (
            O => \N__20382\,
            I => \N__20345\
        );

    \I__4848\ : SRMux
    port map (
            O => \N__20381\,
            I => \N__20340\
        );

    \I__4847\ : Span4Mux_v
    port map (
            O => \N__20376\,
            I => \N__20331\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__20369\,
            I => \N__20331\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__20366\,
            I => \N__20331\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20331\
        );

    \I__4843\ : SRMux
    port map (
            O => \N__20362\,
            I => \N__20328\
        );

    \I__4842\ : SRMux
    port map (
            O => \N__20361\,
            I => \N__20325\
        );

    \I__4841\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20319\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__20357\,
            I => \N__20313\
        );

    \I__4839\ : CascadeMux
    port map (
            O => \N__20356\,
            I => \N__20309\
        );

    \I__4838\ : Span4Mux_v
    port map (
            O => \N__20351\,
            I => \N__20298\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__20348\,
            I => \N__20298\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__20345\,
            I => \N__20298\
        );

    \I__4835\ : SRMux
    port map (
            O => \N__20344\,
            I => \N__20295\
        );

    \I__4834\ : SRMux
    port map (
            O => \N__20343\,
            I => \N__20291\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__20340\,
            I => \N__20288\
        );

    \I__4832\ : Span4Mux_v
    port map (
            O => \N__20331\,
            I => \N__20281\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__20328\,
            I => \N__20281\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__20325\,
            I => \N__20281\
        );

    \I__4829\ : SRMux
    port map (
            O => \N__20324\,
            I => \N__20278\
        );

    \I__4828\ : SRMux
    port map (
            O => \N__20323\,
            I => \N__20275\
        );

    \I__4827\ : SRMux
    port map (
            O => \N__20322\,
            I => \N__20272\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__20319\,
            I => \N__20268\
        );

    \I__4825\ : CascadeMux
    port map (
            O => \N__20318\,
            I => \N__20264\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__20317\,
            I => \N__20260\
        );

    \I__4823\ : CascadeMux
    port map (
            O => \N__20316\,
            I => \N__20256\
        );

    \I__4822\ : IoSpan4Mux
    port map (
            O => \N__20313\,
            I => \N__20252\
        );

    \I__4821\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20247\
        );

    \I__4820\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20247\
        );

    \I__4819\ : SRMux
    port map (
            O => \N__20308\,
            I => \N__20244\
        );

    \I__4818\ : SRMux
    port map (
            O => \N__20307\,
            I => \N__20241\
        );

    \I__4817\ : SRMux
    port map (
            O => \N__20306\,
            I => \N__20238\
        );

    \I__4816\ : SRMux
    port map (
            O => \N__20305\,
            I => \N__20235\
        );

    \I__4815\ : Span4Mux_v
    port map (
            O => \N__20298\,
            I => \N__20229\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__20295\,
            I => \N__20229\
        );

    \I__4813\ : SRMux
    port map (
            O => \N__20294\,
            I => \N__20226\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__20291\,
            I => \N__20223\
        );

    \I__4811\ : Span4Mux_h
    port map (
            O => \N__20288\,
            I => \N__20214\
        );

    \I__4810\ : Span4Mux_v
    port map (
            O => \N__20281\,
            I => \N__20214\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__20278\,
            I => \N__20214\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__20275\,
            I => \N__20214\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__20272\,
            I => \N__20211\
        );

    \I__4806\ : SRMux
    port map (
            O => \N__20271\,
            I => \N__20208\
        );

    \I__4805\ : Span4Mux_h
    port map (
            O => \N__20268\,
            I => \N__20204\
        );

    \I__4804\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20189\
        );

    \I__4803\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20189\
        );

    \I__4802\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20189\
        );

    \I__4801\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20189\
        );

    \I__4800\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20189\
        );

    \I__4799\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20189\
        );

    \I__4798\ : InMux
    port map (
            O => \N__20255\,
            I => \N__20189\
        );

    \I__4797\ : Span4Mux_s2_h
    port map (
            O => \N__20252\,
            I => \N__20185\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__20247\,
            I => \N__20182\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__20244\,
            I => \N__20175\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__20241\,
            I => \N__20175\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__20238\,
            I => \N__20170\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__20235\,
            I => \N__20170\
        );

    \I__4791\ : SRMux
    port map (
            O => \N__20234\,
            I => \N__20167\
        );

    \I__4790\ : Span4Mux_v
    port map (
            O => \N__20229\,
            I => \N__20162\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__20226\,
            I => \N__20162\
        );

    \I__4788\ : Span4Mux_h
    port map (
            O => \N__20223\,
            I => \N__20153\
        );

    \I__4787\ : Span4Mux_v
    port map (
            O => \N__20214\,
            I => \N__20153\
        );

    \I__4786\ : Span4Mux_v
    port map (
            O => \N__20211\,
            I => \N__20153\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__20208\,
            I => \N__20153\
        );

    \I__4784\ : SRMux
    port map (
            O => \N__20207\,
            I => \N__20150\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__20204\,
            I => \N__20144\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__20189\,
            I => \N__20144\
        );

    \I__4781\ : SRMux
    port map (
            O => \N__20188\,
            I => \N__20141\
        );

    \I__4780\ : Span4Mux_h
    port map (
            O => \N__20185\,
            I => \N__20136\
        );

    \I__4779\ : Span4Mux_v
    port map (
            O => \N__20182\,
            I => \N__20136\
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__20181\,
            I => \N__20132\
        );

    \I__4777\ : SRMux
    port map (
            O => \N__20180\,
            I => \N__20128\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__20175\,
            I => \N__20115\
        );

    \I__4775\ : Span4Mux_v
    port map (
            O => \N__20170\,
            I => \N__20115\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__20167\,
            I => \N__20115\
        );

    \I__4773\ : Span4Mux_v
    port map (
            O => \N__20162\,
            I => \N__20115\
        );

    \I__4772\ : Span4Mux_v
    port map (
            O => \N__20153\,
            I => \N__20115\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__20150\,
            I => \N__20115\
        );

    \I__4770\ : SRMux
    port map (
            O => \N__20149\,
            I => \N__20112\
        );

    \I__4769\ : Span4Mux_v
    port map (
            O => \N__20144\,
            I => \N__20109\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__20141\,
            I => \N__20106\
        );

    \I__4767\ : Sp12to4
    port map (
            O => \N__20136\,
            I => \N__20103\
        );

    \I__4766\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20096\
        );

    \I__4765\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20096\
        );

    \I__4764\ : InMux
    port map (
            O => \N__20131\,
            I => \N__20096\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__20128\,
            I => \N__20093\
        );

    \I__4762\ : Span4Mux_v
    port map (
            O => \N__20115\,
            I => \N__20088\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__20112\,
            I => \N__20088\
        );

    \I__4760\ : Span4Mux_h
    port map (
            O => \N__20109\,
            I => \N__20083\
        );

    \I__4759\ : Span4Mux_h
    port map (
            O => \N__20106\,
            I => \N__20083\
        );

    \I__4758\ : Span12Mux_h
    port map (
            O => \N__20103\,
            I => \N__20078\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__20096\,
            I => \N__20078\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__20093\,
            I => \N__20075\
        );

    \I__4755\ : Sp12to4
    port map (
            O => \N__20088\,
            I => \N__20072\
        );

    \I__4754\ : Span4Mux_h
    port map (
            O => \N__20083\,
            I => \N__20069\
        );

    \I__4753\ : Odrv12
    port map (
            O => \N__20078\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4752\ : Odrv4
    port map (
            O => \N__20075\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4751\ : Odrv12
    port map (
            O => \N__20072\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4750\ : Odrv4
    port map (
            O => \N__20069\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4749\ : CascadeMux
    port map (
            O => \N__20060\,
            I => \N__20056\
        );

    \I__4748\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20044\
        );

    \I__4747\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20041\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__20055\,
            I => \N__20036\
        );

    \I__4745\ : CascadeMux
    port map (
            O => \N__20054\,
            I => \N__20033\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__20053\,
            I => \N__20030\
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__20052\,
            I => \N__20027\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__20051\,
            I => \N__20024\
        );

    \I__4741\ : CascadeMux
    port map (
            O => \N__20050\,
            I => \N__20020\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__20049\,
            I => \N__20016\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__20048\,
            I => \N__20012\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__20047\,
            I => \N__20008\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__20044\,
            I => \N__20003\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__20041\,
            I => \N__20003\
        );

    \I__4735\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20000\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__20039\,
            I => \N__19997\
        );

    \I__4733\ : InMux
    port map (
            O => \N__20036\,
            I => \N__19990\
        );

    \I__4732\ : InMux
    port map (
            O => \N__20033\,
            I => \N__19990\
        );

    \I__4731\ : InMux
    port map (
            O => \N__20030\,
            I => \N__19983\
        );

    \I__4730\ : InMux
    port map (
            O => \N__20027\,
            I => \N__19983\
        );

    \I__4729\ : InMux
    port map (
            O => \N__20024\,
            I => \N__19983\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20023\,
            I => \N__19966\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20020\,
            I => \N__19966\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20019\,
            I => \N__19966\
        );

    \I__4725\ : InMux
    port map (
            O => \N__20016\,
            I => \N__19966\
        );

    \I__4724\ : InMux
    port map (
            O => \N__20015\,
            I => \N__19966\
        );

    \I__4723\ : InMux
    port map (
            O => \N__20012\,
            I => \N__19966\
        );

    \I__4722\ : InMux
    port map (
            O => \N__20011\,
            I => \N__19966\
        );

    \I__4721\ : InMux
    port map (
            O => \N__20008\,
            I => \N__19966\
        );

    \I__4720\ : Span4Mux_s2_h
    port map (
            O => \N__20003\,
            I => \N__19962\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__20000\,
            I => \N__19959\
        );

    \I__4718\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19956\
        );

    \I__4717\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19951\
        );

    \I__4716\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19951\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__19990\,
            I => \N__19944\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__19983\,
            I => \N__19944\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__19966\,
            I => \N__19944\
        );

    \I__4712\ : InMux
    port map (
            O => \N__19965\,
            I => \N__19940\
        );

    \I__4711\ : Span4Mux_h
    port map (
            O => \N__19962\,
            I => \N__19937\
        );

    \I__4710\ : Span4Mux_v
    port map (
            O => \N__19959\,
            I => \N__19932\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__19956\,
            I => \N__19932\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__19951\,
            I => \N__19927\
        );

    \I__4707\ : Span4Mux_v
    port map (
            O => \N__19944\,
            I => \N__19927\
        );

    \I__4706\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19924\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__19940\,
            I => \N__19921\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__19937\,
            I => \N__19918\
        );

    \I__4703\ : Span4Mux_h
    port map (
            O => \N__19932\,
            I => \N__19911\
        );

    \I__4702\ : Span4Mux_h
    port map (
            O => \N__19927\,
            I => \N__19911\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__19924\,
            I => \N__19911\
        );

    \I__4700\ : Span4Mux_h
    port map (
            O => \N__19921\,
            I => \N__19908\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__19918\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4698\ : Odrv4
    port map (
            O => \N__19911\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__19908\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4696\ : IoInMux
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__4694\ : Span4Mux_s1_v
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__4693\ : Sp12to4
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__4692\ : Span12Mux_h
    port map (
            O => \N__19889\,
            I => \N__19885\
        );

    \I__4691\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19882\
        );

    \I__4690\ : Odrv12
    port map (
            O => \N__19885\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__19882\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__4688\ : IoInMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__4686\ : IoSpan4Mux
    port map (
            O => \N__19871\,
            I => \N__19868\
        );

    \I__4685\ : Sp12to4
    port map (
            O => \N__19868\,
            I => \N__19864\
        );

    \I__4684\ : InMux
    port map (
            O => \N__19867\,
            I => \N__19861\
        );

    \I__4683\ : Odrv12
    port map (
            O => \N__19864\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__19861\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__4681\ : InMux
    port map (
            O => \N__19856\,
            I => \un1_M_this_external_address_q_cry_0\
        );

    \I__4680\ : IoInMux
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__4678\ : IoSpan4Mux
    port map (
            O => \N__19847\,
            I => \N__19844\
        );

    \I__4677\ : IoSpan4Mux
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__4676\ : Span4Mux_s2_v
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__4675\ : Span4Mux_v
    port map (
            O => \N__19838\,
            I => \N__19834\
        );

    \I__4674\ : InMux
    port map (
            O => \N__19837\,
            I => \N__19831\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__19834\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__19831\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__4671\ : InMux
    port map (
            O => \N__19826\,
            I => \un1_M_this_external_address_q_cry_1\
        );

    \I__4670\ : IoInMux
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__4668\ : Span4Mux_s2_h
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__4667\ : Span4Mux_v
    port map (
            O => \N__19814\,
            I => \N__19810\
        );

    \I__4666\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19807\
        );

    \I__4665\ : Odrv4
    port map (
            O => \N__19810\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__19807\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__4663\ : InMux
    port map (
            O => \N__19802\,
            I => \un1_M_this_external_address_q_cry_2\
        );

    \I__4662\ : IoInMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__19796\,
            I => \N__19792\
        );

    \I__4660\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19789\
        );

    \I__4659\ : Odrv4
    port map (
            O => \N__19792\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__19789\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__4657\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__19778\,
            I => \this_vram.mem_out_bus5_1\
        );

    \I__4654\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__19769\,
            I => \this_vram.mem_mem_1_0_RNISSK11Z0Z_0\
        );

    \I__4651\ : InMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__4649\ : Span4Mux_v
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__19757\,
            I => \this_vram.mem_out_bus5_2\
        );

    \I__4647\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__4645\ : Span4Mux_v
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__4644\ : Span4Mux_v
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__4643\ : Odrv4
    port map (
            O => \N__19742\,
            I => \this_vram.mem_out_bus1_2\
        );

    \I__4642\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__19736\,
            I => \this_vram.mem_mem_1_1_RNIUSKZ0Z11\
        );

    \I__4640\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__4637\ : Sp12to4
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__4636\ : Odrv12
    port map (
            O => \N__19721\,
            I => \this_vram.mem_out_bus7_2\
        );

    \I__4635\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__4633\ : Span4Mux_h
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__4632\ : Odrv4
    port map (
            O => \N__19709\,
            I => \this_vram.mem_out_bus3_2\
        );

    \I__4631\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__19703\,
            I => \this_vram.mem_mem_3_1_RNI25PZ0Z11\
        );

    \I__4629\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19697\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__4627\ : Span4Mux_v
    port map (
            O => \N__19694\,
            I => \N__19691\
        );

    \I__4626\ : Span4Mux_v
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__4625\ : Odrv4
    port map (
            O => \N__19688\,
            I => \this_vram.mem_out_bus7_0\
        );

    \I__4624\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19682\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__4622\ : Span4Mux_v
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__19673\,
            I => \this_vram.mem_out_bus3_0\
        );

    \I__4619\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__19667\,
            I => \this_vram.mem_mem_3_0_RNI05PZ0Z11\
        );

    \I__4617\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__4615\ : Span4Mux_v
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__4614\ : Odrv4
    port map (
            O => \N__19655\,
            I => \this_vram.mem_out_bus2_2\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__4612\ : InMux
    port map (
            O => \N__19649\,
            I => \N__19646\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__4610\ : Sp12to4
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__4609\ : Odrv12
    port map (
            O => \N__19640\,
            I => \this_vram.mem_out_bus6_2\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__4607\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__19631\,
            I => \this_vram.mem_mem_2_1_RNI01NZ0Z11\
        );

    \I__4605\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19612\
        );

    \I__4604\ : InMux
    port map (
            O => \N__19627\,
            I => \N__19601\
        );

    \I__4603\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19601\
        );

    \I__4602\ : InMux
    port map (
            O => \N__19625\,
            I => \N__19601\
        );

    \I__4601\ : InMux
    port map (
            O => \N__19624\,
            I => \N__19601\
        );

    \I__4600\ : InMux
    port map (
            O => \N__19623\,
            I => \N__19601\
        );

    \I__4599\ : InMux
    port map (
            O => \N__19622\,
            I => \N__19598\
        );

    \I__4598\ : InMux
    port map (
            O => \N__19621\,
            I => \N__19593\
        );

    \I__4597\ : InMux
    port map (
            O => \N__19620\,
            I => \N__19593\
        );

    \I__4596\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19590\
        );

    \I__4595\ : InMux
    port map (
            O => \N__19618\,
            I => \N__19587\
        );

    \I__4594\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19580\
        );

    \I__4593\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19580\
        );

    \I__4592\ : InMux
    port map (
            O => \N__19615\,
            I => \N__19580\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__19612\,
            I => \N__19571\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__19601\,
            I => \N__19571\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19571\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__19593\,
            I => \N__19571\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__19590\,
            I => \N__19564\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__19587\,
            I => \N__19564\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__19580\,
            I => \N__19564\
        );

    \I__4584\ : Span4Mux_v
    port map (
            O => \N__19571\,
            I => \N__19561\
        );

    \I__4583\ : Span4Mux_h
    port map (
            O => \N__19564\,
            I => \N__19558\
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__19561\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__4581\ : Odrv4
    port map (
            O => \N__19558\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__4580\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19550\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__4578\ : Odrv4
    port map (
            O => \N__19547\,
            I => \this_vram.mem_out_bus5_0\
        );

    \I__4577\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__4575\ : Span4Mux_v
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__4574\ : Span4Mux_v
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__4573\ : Span4Mux_v
    port map (
            O => \N__19532\,
            I => \N__19529\
        );

    \I__4572\ : Odrv4
    port map (
            O => \N__19529\,
            I => \this_vram.mem_out_bus1_0\
        );

    \I__4571\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__19523\,
            I => \this_vram.mem_mem_1_0_RNISSKZ0Z11\
        );

    \I__4569\ : CascadeMux
    port map (
            O => \N__19520\,
            I => \N__19516\
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__19519\,
            I => \N__19513\
        );

    \I__4567\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19510\
        );

    \I__4566\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19507\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__19510\,
            I => \N__19503\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__19507\,
            I => \N__19500\
        );

    \I__4563\ : InMux
    port map (
            O => \N__19506\,
            I => \N__19497\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__19503\,
            I => \N__19494\
        );

    \I__4561\ : Span4Mux_h
    port map (
            O => \N__19500\,
            I => \N__19491\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__19497\,
            I => \N__19488\
        );

    \I__4559\ : Sp12to4
    port map (
            O => \N__19494\,
            I => \N__19485\
        );

    \I__4558\ : Span4Mux_h
    port map (
            O => \N__19491\,
            I => \N__19480\
        );

    \I__4557\ : Span4Mux_v
    port map (
            O => \N__19488\,
            I => \N__19480\
        );

    \I__4556\ : Span12Mux_h
    port map (
            O => \N__19485\,
            I => \N__19477\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__19480\,
            I => \N__19474\
        );

    \I__4554\ : Span12Mux_v
    port map (
            O => \N__19477\,
            I => \N__19471\
        );

    \I__4553\ : Sp12to4
    port map (
            O => \N__19474\,
            I => \N__19468\
        );

    \I__4552\ : Odrv12
    port map (
            O => \N__19471\,
            I => port_data_c_3
        );

    \I__4551\ : Odrv12
    port map (
            O => \N__19468\,
            I => port_data_c_3
        );

    \I__4550\ : CascadeMux
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__4549\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19457\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__19457\,
            I => \N__19454\
        );

    \I__4547\ : Span4Mux_h
    port map (
            O => \N__19454\,
            I => \N__19451\
        );

    \I__4546\ : Sp12to4
    port map (
            O => \N__19451\,
            I => \N__19448\
        );

    \I__4545\ : Span12Mux_v
    port map (
            O => \N__19448\,
            I => \N__19445\
        );

    \I__4544\ : Odrv12
    port map (
            O => \N__19445\,
            I => port_data_c_7
        );

    \I__4543\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19439\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__19439\,
            I => \N__19435\
        );

    \I__4541\ : InMux
    port map (
            O => \N__19438\,
            I => \N__19432\
        );

    \I__4540\ : Span4Mux_v
    port map (
            O => \N__19435\,
            I => \N__19425\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__19432\,
            I => \N__19425\
        );

    \I__4538\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19422\
        );

    \I__4537\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19418\
        );

    \I__4536\ : Span4Mux_v
    port map (
            O => \N__19425\,
            I => \N__19412\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__19422\,
            I => \N__19412\
        );

    \I__4534\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19409\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__19418\,
            I => \N__19406\
        );

    \I__4532\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19403\
        );

    \I__4531\ : Span4Mux_v
    port map (
            O => \N__19412\,
            I => \N__19397\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__19409\,
            I => \N__19397\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__19406\,
            I => \N__19392\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__19403\,
            I => \N__19392\
        );

    \I__4527\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19389\
        );

    \I__4526\ : Span4Mux_v
    port map (
            O => \N__19397\,
            I => \N__19385\
        );

    \I__4525\ : Span4Mux_v
    port map (
            O => \N__19392\,
            I => \N__19380\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__19389\,
            I => \N__19380\
        );

    \I__4523\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19377\
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__19385\,
            I => \M_this_vram_write_data_0_i_3\
        );

    \I__4521\ : Odrv4
    port map (
            O => \N__19380\,
            I => \M_this_vram_write_data_0_i_3\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__19377\,
            I => \M_this_vram_write_data_0_i_3\
        );

    \I__4519\ : CEMux
    port map (
            O => \N__19370\,
            I => \N__19366\
        );

    \I__4518\ : CEMux
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__19366\,
            I => \N__19360\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__19363\,
            I => \N__19357\
        );

    \I__4515\ : Span4Mux_v
    port map (
            O => \N__19360\,
            I => \N__19354\
        );

    \I__4514\ : Span4Mux_h
    port map (
            O => \N__19357\,
            I => \N__19351\
        );

    \I__4513\ : Span4Mux_h
    port map (
            O => \N__19354\,
            I => \N__19348\
        );

    \I__4512\ : Span4Mux_h
    port map (
            O => \N__19351\,
            I => \N__19345\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__19348\,
            I => \this_vram.mem_WE_4\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__19345\,
            I => \this_vram.mem_WE_4\
        );

    \I__4509\ : InMux
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__4507\ : Odrv4
    port map (
            O => \N__19334\,
            I => \this_vram.mem_mem_0_1_RNISOIZ0Z11\
        );

    \I__4506\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19328\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__19328\,
            I => \N__19325\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__19325\,
            I => \N__19322\
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__19322\,
            I => \this_vram.mem_out_bus5_3\
        );

    \I__4502\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__4500\ : Span4Mux_v
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__4499\ : Span4Mux_v
    port map (
            O => \N__19310\,
            I => \N__19307\
        );

    \I__4498\ : Odrv4
    port map (
            O => \N__19307\,
            I => \this_vram.mem_out_bus1_3\
        );

    \I__4497\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__19301\,
            I => \N__19298\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__19298\,
            I => \this_vram.mem_out_bus3_3\
        );

    \I__4494\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__4492\ : Sp12to4
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__4491\ : Span12Mux_v
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__4490\ : Odrv12
    port map (
            O => \N__19283\,
            I => \this_vram.mem_out_bus7_3\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__19280\,
            I => \this_vram.mem_DOUT_6_i_m2_ns_1_3_cascade_\
        );

    \I__4488\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__19274\,
            I => \this_vram.mem_N_102\
        );

    \I__4486\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__4484\ : Span4Mux_h
    port map (
            O => \N__19265\,
            I => \N__19262\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__19262\,
            I => \this_vram.mem_out_bus4_3\
        );

    \I__4482\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19256\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__19256\,
            I => \N__19253\
        );

    \I__4480\ : Sp12to4
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__4479\ : Span12Mux_v
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__4478\ : Odrv12
    port map (
            O => \N__19247\,
            I => \this_vram.mem_out_bus0_3\
        );

    \I__4477\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19241\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__4475\ : Span4Mux_v
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__4474\ : Span4Mux_v
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__19232\,
            I => \this_vram.mem_out_bus6_3\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19229\,
            I => \N__19226\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__4470\ : Span4Mux_v
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__4469\ : Odrv4
    port map (
            O => \N__19220\,
            I => \this_vram.mem_out_bus2_3\
        );

    \I__4468\ : CascadeMux
    port map (
            O => \N__19217\,
            I => \this_vram.mem_DOUT_3_i_m2_ns_1_3_cascade_\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__19214\,
            I => \N__19206\
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__19213\,
            I => \N__19203\
        );

    \I__4465\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19200\
        );

    \I__4464\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19196\
        );

    \I__4463\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19187\
        );

    \I__4462\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19187\
        );

    \I__4461\ : InMux
    port map (
            O => \N__19206\,
            I => \N__19187\
        );

    \I__4460\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19187\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__19200\,
            I => \N__19184\
        );

    \I__4458\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19181\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__19196\,
            I => \N__19178\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__19187\,
            I => \N__19175\
        );

    \I__4455\ : Span4Mux_h
    port map (
            O => \N__19184\,
            I => \N__19172\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__19181\,
            I => \N__19165\
        );

    \I__4453\ : Span4Mux_v
    port map (
            O => \N__19178\,
            I => \N__19165\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__19175\,
            I => \N__19165\
        );

    \I__4451\ : Odrv4
    port map (
            O => \N__19172\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__4450\ : Odrv4
    port map (
            O => \N__19165\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__4449\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__19157\,
            I => \this_vram.mem_N_105\
        );

    \I__4447\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__4445\ : Sp12to4
    port map (
            O => \N__19148\,
            I => \N__19145\
        );

    \I__4444\ : Span12Mux_v
    port map (
            O => \N__19145\,
            I => \N__19142\
        );

    \I__4443\ : Odrv12
    port map (
            O => \N__19142\,
            I => \this_vram.mem_out_bus0_0\
        );

    \I__4442\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__19136\,
            I => \this_vram.mem_out_bus4_0\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__19133\,
            I => \N__19130\
        );

    \I__4439\ : InMux
    port map (
            O => \N__19130\,
            I => \N__19127\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__19127\,
            I => \this_vram.mem_mem_0_0_RNIQOIZ0Z11\
        );

    \I__4437\ : InMux
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__4435\ : Sp12to4
    port map (
            O => \N__19118\,
            I => \N__19115\
        );

    \I__4434\ : Odrv12
    port map (
            O => \N__19115\,
            I => \this_vram.mem_out_bus6_0\
        );

    \I__4433\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__19109\,
            I => \N__19106\
        );

    \I__4431\ : Span4Mux_v
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__4430\ : Span4Mux_v
    port map (
            O => \N__19103\,
            I => \N__19100\
        );

    \I__4429\ : Odrv4
    port map (
            O => \N__19100\,
            I => \this_vram.mem_out_bus2_0\
        );

    \I__4428\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__19094\,
            I => \this_vram.mem_mem_2_0_RNIU0NZ0Z11\
        );

    \I__4426\ : CEMux
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__19088\,
            I => \N__19084\
        );

    \I__4424\ : CEMux
    port map (
            O => \N__19087\,
            I => \N__19081\
        );

    \I__4423\ : Span4Mux_h
    port map (
            O => \N__19084\,
            I => \N__19078\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__19081\,
            I => \N__19075\
        );

    \I__4421\ : Odrv4
    port map (
            O => \N__19078\,
            I => \this_vram.mem_WE_6\
        );

    \I__4420\ : Odrv12
    port map (
            O => \N__19075\,
            I => \this_vram.mem_WE_6\
        );

    \I__4419\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__4417\ : Sp12to4
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__4416\ : Span12Mux_v
    port map (
            O => \N__19061\,
            I => \N__19058\
        );

    \I__4415\ : Odrv12
    port map (
            O => \N__19058\,
            I => \this_vram.mem_out_bus1_1\
        );

    \I__4414\ : InMux
    port map (
            O => \N__19055\,
            I => \N__19048\
        );

    \I__4413\ : InMux
    port map (
            O => \N__19054\,
            I => \N__19048\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__19053\,
            I => \N__19045\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__19048\,
            I => \N__19042\
        );

    \I__4410\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19039\
        );

    \I__4409\ : Span4Mux_h
    port map (
            O => \N__19042\,
            I => \N__19036\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__19039\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__19036\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4406\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19027\
        );

    \I__4405\ : InMux
    port map (
            O => \N__19030\,
            I => \N__19024\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__19027\,
            I => \N__19020\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19024\,
            I => \N__19016\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19023\,
            I => \N__19011\
        );

    \I__4401\ : Span4Mux_v
    port map (
            O => \N__19020\,
            I => \N__19008\
        );

    \I__4400\ : InMux
    port map (
            O => \N__19019\,
            I => \N__19005\
        );

    \I__4399\ : Span4Mux_v
    port map (
            O => \N__19016\,
            I => \N__19002\
        );

    \I__4398\ : InMux
    port map (
            O => \N__19015\,
            I => \N__18999\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19014\,
            I => \N__18996\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__19011\,
            I => \N__18989\
        );

    \I__4395\ : Sp12to4
    port map (
            O => \N__19008\,
            I => \N__18989\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__19005\,
            I => \N__18989\
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__19002\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__18999\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__18996\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4390\ : Odrv12
    port map (
            O => \N__18989\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__18980\,
            I => \N__18976\
        );

    \I__4388\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18972\
        );

    \I__4387\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18969\
        );

    \I__4386\ : InMux
    port map (
            O => \N__18975\,
            I => \N__18966\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__18972\,
            I => \N__18963\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__18969\,
            I => \N__18960\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__18966\,
            I => \N__18957\
        );

    \I__4382\ : Span4Mux_v
    port map (
            O => \N__18963\,
            I => \N__18952\
        );

    \I__4381\ : Span4Mux_v
    port map (
            O => \N__18960\,
            I => \N__18952\
        );

    \I__4380\ : Span4Mux_v
    port map (
            O => \N__18957\,
            I => \N__18949\
        );

    \I__4379\ : Sp12to4
    port map (
            O => \N__18952\,
            I => \N__18944\
        );

    \I__4378\ : Sp12to4
    port map (
            O => \N__18949\,
            I => \N__18944\
        );

    \I__4377\ : Span12Mux_h
    port map (
            O => \N__18944\,
            I => \N__18941\
        );

    \I__4376\ : Odrv12
    port map (
            O => \N__18941\,
            I => port_data_c_0
        );

    \I__4375\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18934\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__18937\,
            I => \N__18930\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__18934\,
            I => \N__18927\
        );

    \I__4372\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18924\
        );

    \I__4371\ : InMux
    port map (
            O => \N__18930\,
            I => \N__18921\
        );

    \I__4370\ : Span4Mux_v
    port map (
            O => \N__18927\,
            I => \N__18918\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__18924\,
            I => \N__18915\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__18921\,
            I => \N__18912\
        );

    \I__4367\ : Span4Mux_h
    port map (
            O => \N__18918\,
            I => \N__18907\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__18915\,
            I => \N__18907\
        );

    \I__4365\ : Span12Mux_v
    port map (
            O => \N__18912\,
            I => \N__18904\
        );

    \I__4364\ : Span4Mux_v
    port map (
            O => \N__18907\,
            I => \N__18901\
        );

    \I__4363\ : Span12Mux_h
    port map (
            O => \N__18904\,
            I => \N__18898\
        );

    \I__4362\ : Sp12to4
    port map (
            O => \N__18901\,
            I => \N__18895\
        );

    \I__4361\ : Odrv12
    port map (
            O => \N__18898\,
            I => port_data_c_4
        );

    \I__4360\ : Odrv12
    port map (
            O => \N__18895\,
            I => port_data_c_4
        );

    \I__4359\ : CascadeMux
    port map (
            O => \N__18890\,
            I => \M_this_vram_write_data_0_sqmuxa_cascade_\
        );

    \I__4358\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__18884\,
            I => \N__18880\
        );

    \I__4356\ : InMux
    port map (
            O => \N__18883\,
            I => \N__18877\
        );

    \I__4355\ : Span4Mux_h
    port map (
            O => \N__18880\,
            I => \N__18873\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__18877\,
            I => \N__18870\
        );

    \I__4353\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18867\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__18873\,
            I => \N__18860\
        );

    \I__4351\ : Span4Mux_h
    port map (
            O => \N__18870\,
            I => \N__18860\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__18867\,
            I => \N__18857\
        );

    \I__4349\ : InMux
    port map (
            O => \N__18866\,
            I => \N__18854\
        );

    \I__4348\ : InMux
    port map (
            O => \N__18865\,
            I => \N__18850\
        );

    \I__4347\ : Span4Mux_v
    port map (
            O => \N__18860\,
            I => \N__18844\
        );

    \I__4346\ : Span4Mux_h
    port map (
            O => \N__18857\,
            I => \N__18844\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__18854\,
            I => \N__18841\
        );

    \I__4344\ : InMux
    port map (
            O => \N__18853\,
            I => \N__18838\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__18850\,
            I => \N__18835\
        );

    \I__4342\ : InMux
    port map (
            O => \N__18849\,
            I => \N__18832\
        );

    \I__4341\ : Span4Mux_v
    port map (
            O => \N__18844\,
            I => \N__18826\
        );

    \I__4340\ : Span4Mux_h
    port map (
            O => \N__18841\,
            I => \N__18826\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__18838\,
            I => \N__18823\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__18835\,
            I => \N__18818\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__18832\,
            I => \N__18818\
        );

    \I__4336\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18815\
        );

    \I__4335\ : Span4Mux_v
    port map (
            O => \N__18826\,
            I => \N__18810\
        );

    \I__4334\ : Span4Mux_h
    port map (
            O => \N__18823\,
            I => \N__18810\
        );

    \I__4333\ : Span4Mux_v
    port map (
            O => \N__18818\,
            I => \N__18805\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__18815\,
            I => \N__18805\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__18810\,
            I => \M_this_vram_write_data_0_i_0\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__18805\,
            I => \M_this_vram_write_data_0_i_0\
        );

    \I__4329\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18787\
        );

    \I__4328\ : InMux
    port map (
            O => \N__18799\,
            I => \N__18784\
        );

    \I__4327\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18780\
        );

    \I__4326\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18777\
        );

    \I__4325\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18772\
        );

    \I__4324\ : InMux
    port map (
            O => \N__18795\,
            I => \N__18772\
        );

    \I__4323\ : InMux
    port map (
            O => \N__18794\,
            I => \N__18764\
        );

    \I__4322\ : InMux
    port map (
            O => \N__18793\,
            I => \N__18764\
        );

    \I__4321\ : InMux
    port map (
            O => \N__18792\,
            I => \N__18764\
        );

    \I__4320\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18756\
        );

    \I__4319\ : InMux
    port map (
            O => \N__18790\,
            I => \N__18756\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__18787\,
            I => \N__18751\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__18784\,
            I => \N__18751\
        );

    \I__4316\ : InMux
    port map (
            O => \N__18783\,
            I => \N__18748\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__18780\,
            I => \N__18741\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__18777\,
            I => \N__18741\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__18772\,
            I => \N__18741\
        );

    \I__4312\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18733\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__18764\,
            I => \N__18730\
        );

    \I__4310\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18725\
        );

    \I__4309\ : InMux
    port map (
            O => \N__18762\,
            I => \N__18725\
        );

    \I__4308\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18722\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__18756\,
            I => \N__18717\
        );

    \I__4306\ : Span12Mux_h
    port map (
            O => \N__18751\,
            I => \N__18717\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__18748\,
            I => \N__18712\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__18741\,
            I => \N__18712\
        );

    \I__4303\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18709\
        );

    \I__4302\ : InMux
    port map (
            O => \N__18739\,
            I => \N__18700\
        );

    \I__4301\ : InMux
    port map (
            O => \N__18738\,
            I => \N__18700\
        );

    \I__4300\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18700\
        );

    \I__4299\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18700\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__18733\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4297\ : Odrv4
    port map (
            O => \N__18730\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__18725\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__18722\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4294\ : Odrv12
    port map (
            O => \N__18717\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__18712\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__18709\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__18700\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4290\ : InMux
    port map (
            O => \N__18683\,
            I => \N__18679\
        );

    \I__4289\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18676\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__18679\,
            I => \N__18673\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__18676\,
            I => \this_start_data_delay.N_351_0\
        );

    \I__4286\ : Odrv12
    port map (
            O => \N__18673\,
            I => \this_start_data_delay.N_351_0\
        );

    \I__4285\ : CEMux
    port map (
            O => \N__18668\,
            I => \N__18665\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__18665\,
            I => \N__18662\
        );

    \I__4283\ : Span12Mux_s8_h
    port map (
            O => \N__18662\,
            I => \N__18658\
        );

    \I__4282\ : CEMux
    port map (
            O => \N__18661\,
            I => \N__18655\
        );

    \I__4281\ : Odrv12
    port map (
            O => \N__18658\,
            I => \this_vram.mem_WE_8\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__18655\,
            I => \this_vram.mem_WE_8\
        );

    \I__4279\ : CEMux
    port map (
            O => \N__18650\,
            I => \N__18647\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__18647\,
            I => \N__18643\
        );

    \I__4277\ : CEMux
    port map (
            O => \N__18646\,
            I => \N__18640\
        );

    \I__4276\ : Span4Mux_v
    port map (
            O => \N__18643\,
            I => \N__18637\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__18640\,
            I => \N__18634\
        );

    \I__4274\ : Span4Mux_v
    port map (
            O => \N__18637\,
            I => \N__18631\
        );

    \I__4273\ : Span12Mux_s8_h
    port map (
            O => \N__18634\,
            I => \N__18628\
        );

    \I__4272\ : Odrv4
    port map (
            O => \N__18631\,
            I => \this_vram.mem_WE_12\
        );

    \I__4271\ : Odrv12
    port map (
            O => \N__18628\,
            I => \this_vram.mem_WE_12\
        );

    \I__4270\ : CEMux
    port map (
            O => \N__18623\,
            I => \N__18619\
        );

    \I__4269\ : CEMux
    port map (
            O => \N__18622\,
            I => \N__18616\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__18619\,
            I => \N__18613\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__18616\,
            I => \N__18610\
        );

    \I__4266\ : Span4Mux_v
    port map (
            O => \N__18613\,
            I => \N__18605\
        );

    \I__4265\ : Span4Mux_h
    port map (
            O => \N__18610\,
            I => \N__18605\
        );

    \I__4264\ : Odrv4
    port map (
            O => \N__18605\,
            I => \this_vram.mem_WE_10\
        );

    \I__4263\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18599\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__4261\ : Span4Mux_h
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__18593\,
            I => \this_vram.mem_out_bus4_2\
        );

    \I__4259\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18587\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__18587\,
            I => \N__18584\
        );

    \I__4257\ : Sp12to4
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__4256\ : Span12Mux_v
    port map (
            O => \N__18581\,
            I => \N__18578\
        );

    \I__4255\ : Odrv12
    port map (
            O => \N__18578\,
            I => \this_vram.mem_out_bus0_2\
        );

    \I__4254\ : CEMux
    port map (
            O => \N__18575\,
            I => \N__18571\
        );

    \I__4253\ : CEMux
    port map (
            O => \N__18574\,
            I => \N__18568\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__18571\,
            I => \N__18565\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__18568\,
            I => \N__18562\
        );

    \I__4250\ : Span4Mux_h
    port map (
            O => \N__18565\,
            I => \N__18559\
        );

    \I__4249\ : Span4Mux_h
    port map (
            O => \N__18562\,
            I => \N__18556\
        );

    \I__4248\ : Span4Mux_v
    port map (
            O => \N__18559\,
            I => \N__18553\
        );

    \I__4247\ : Sp12to4
    port map (
            O => \N__18556\,
            I => \N__18550\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__18553\,
            I => \N__18547\
        );

    \I__4245\ : Odrv12
    port map (
            O => \N__18550\,
            I => \this_vram.mem_WE_14\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__18547\,
            I => \this_vram.mem_WE_14\
        );

    \I__4243\ : InMux
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__18536\,
            I => \N__18533\
        );

    \I__4240\ : Span4Mux_v
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__4239\ : Odrv4
    port map (
            O => \N__18530\,
            I => \this_vram.mem_out_bus6_1\
        );

    \I__4238\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__4236\ : Span4Mux_v
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__4234\ : Odrv4
    port map (
            O => \N__18515\,
            I => \this_vram.mem_out_bus2_1\
        );

    \I__4233\ : InMux
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__18509\,
            I => \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0\
        );

    \I__4231\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__4228\ : Span4Mux_v
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__4227\ : Span4Mux_v
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__4226\ : Odrv4
    port map (
            O => \N__18491\,
            I => \this_vram.mem_out_bus7_1\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__4223\ : Span4Mux_v
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__4222\ : Span4Mux_v
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__18476\,
            I => \this_vram.mem_out_bus3_1\
        );

    \I__4220\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__18470\,
            I => \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__18467\,
            I => \N__18463\
        );

    \I__4217\ : InMux
    port map (
            O => \N__18466\,
            I => \N__18456\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18463\,
            I => \N__18451\
        );

    \I__4215\ : InMux
    port map (
            O => \N__18462\,
            I => \N__18451\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18444\
        );

    \I__4213\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18444\
        );

    \I__4212\ : InMux
    port map (
            O => \N__18459\,
            I => \N__18444\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__18456\,
            I => \N__18441\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__18451\,
            I => \N__18436\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__18444\,
            I => \N__18436\
        );

    \I__4208\ : Span4Mux_v
    port map (
            O => \N__18441\,
            I => \N__18431\
        );

    \I__4207\ : Span4Mux_v
    port map (
            O => \N__18436\,
            I => \N__18431\
        );

    \I__4206\ : Sp12to4
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__4205\ : Span12Mux_h
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__4204\ : Odrv12
    port map (
            O => \N__18425\,
            I => \M_this_vram_read_data_3\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__18422\,
            I => \this_vram.mem_DOUT_7_i_m2_ns_1_2_cascade_\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__18419\,
            I => \N__18414\
        );

    \I__4201\ : CascadeMux
    port map (
            O => \N__18418\,
            I => \N__18409\
        );

    \I__4200\ : CascadeMux
    port map (
            O => \N__18417\,
            I => \N__18406\
        );

    \I__4199\ : InMux
    port map (
            O => \N__18414\,
            I => \N__18403\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__18413\,
            I => \N__18400\
        );

    \I__4197\ : InMux
    port map (
            O => \N__18412\,
            I => \N__18393\
        );

    \I__4196\ : InMux
    port map (
            O => \N__18409\,
            I => \N__18393\
        );

    \I__4195\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18393\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__18403\,
            I => \N__18390\
        );

    \I__4193\ : InMux
    port map (
            O => \N__18400\,
            I => \N__18387\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__18393\,
            I => \N__18384\
        );

    \I__4191\ : Span12Mux_s10_h
    port map (
            O => \N__18390\,
            I => \N__18381\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__18387\,
            I => \N__18376\
        );

    \I__4189\ : Span12Mux_s5_h
    port map (
            O => \N__18384\,
            I => \N__18376\
        );

    \I__4188\ : Span12Mux_h
    port map (
            O => \N__18381\,
            I => \N__18373\
        );

    \I__4187\ : Span12Mux_h
    port map (
            O => \N__18376\,
            I => \N__18370\
        );

    \I__4186\ : Odrv12
    port map (
            O => \N__18373\,
            I => \M_this_vram_read_data_2\
        );

    \I__4185\ : Odrv12
    port map (
            O => \N__18370\,
            I => \M_this_vram_read_data_2\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__18365\,
            I => \N__18360\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__18364\,
            I => \N__18356\
        );

    \I__4182\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18352\
        );

    \I__4181\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18347\
        );

    \I__4180\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18340\
        );

    \I__4179\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18340\
        );

    \I__4178\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18340\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__18352\,
            I => \N__18337\
        );

    \I__4176\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18332\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18332\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__18347\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__18340\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__18337\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__18332\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__4170\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__18320\,
            I => \this_vram.mem_DOUT_7_i_m2_ns_1_0\
        );

    \I__4168\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18314\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__18314\,
            I => \N__18311\
        );

    \I__4166\ : Span4Mux_v
    port map (
            O => \N__18311\,
            I => \N__18303\
        );

    \I__4165\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18296\
        );

    \I__4164\ : InMux
    port map (
            O => \N__18309\,
            I => \N__18296\
        );

    \I__4163\ : InMux
    port map (
            O => \N__18308\,
            I => \N__18296\
        );

    \I__4162\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18291\
        );

    \I__4161\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18291\
        );

    \I__4160\ : Sp12to4
    port map (
            O => \N__18303\,
            I => \N__18284\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__18296\,
            I => \N__18284\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__18291\,
            I => \N__18284\
        );

    \I__4157\ : Span12Mux_s11_h
    port map (
            O => \N__18284\,
            I => \N__18281\
        );

    \I__4156\ : Odrv12
    port map (
            O => \N__18281\,
            I => \M_this_vram_read_data_0\
        );

    \I__4155\ : CascadeMux
    port map (
            O => \N__18278\,
            I => \N__18275\
        );

    \I__4154\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18271\
        );

    \I__4153\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18267\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__18271\,
            I => \N__18264\
        );

    \I__4151\ : CascadeMux
    port map (
            O => \N__18270\,
            I => \N__18261\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__18267\,
            I => \N__18258\
        );

    \I__4149\ : Span4Mux_v
    port map (
            O => \N__18264\,
            I => \N__18255\
        );

    \I__4148\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18252\
        );

    \I__4147\ : Span4Mux_v
    port map (
            O => \N__18258\,
            I => \N__18249\
        );

    \I__4146\ : Span4Mux_h
    port map (
            O => \N__18255\,
            I => \N__18244\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__18252\,
            I => \N__18244\
        );

    \I__4144\ : Span4Mux_v
    port map (
            O => \N__18249\,
            I => \N__18241\
        );

    \I__4143\ : Span4Mux_v
    port map (
            O => \N__18244\,
            I => \N__18238\
        );

    \I__4142\ : Sp12to4
    port map (
            O => \N__18241\,
            I => \N__18233\
        );

    \I__4141\ : Sp12to4
    port map (
            O => \N__18238\,
            I => \N__18233\
        );

    \I__4140\ : Span12Mux_h
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__4139\ : Odrv12
    port map (
            O => \N__18230\,
            I => port_data_c_1
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__18227\,
            I => \N__18223\
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__18226\,
            I => \N__18220\
        );

    \I__4136\ : InMux
    port map (
            O => \N__18223\,
            I => \N__18216\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18220\,
            I => \N__18213\
        );

    \I__4134\ : CascadeMux
    port map (
            O => \N__18219\,
            I => \N__18210\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__18216\,
            I => \N__18205\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__18213\,
            I => \N__18205\
        );

    \I__4131\ : InMux
    port map (
            O => \N__18210\,
            I => \N__18202\
        );

    \I__4130\ : Span4Mux_v
    port map (
            O => \N__18205\,
            I => \N__18199\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__18202\,
            I => \N__18196\
        );

    \I__4128\ : Span4Mux_h
    port map (
            O => \N__18199\,
            I => \N__18191\
        );

    \I__4127\ : Span4Mux_v
    port map (
            O => \N__18196\,
            I => \N__18191\
        );

    \I__4126\ : Sp12to4
    port map (
            O => \N__18191\,
            I => \N__18188\
        );

    \I__4125\ : Odrv12
    port map (
            O => \N__18188\,
            I => port_data_c_5
        );

    \I__4124\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18181\
        );

    \I__4123\ : InMux
    port map (
            O => \N__18184\,
            I => \N__18177\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__18181\,
            I => \N__18172\
        );

    \I__4121\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18168\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__18177\,
            I => \N__18165\
        );

    \I__4119\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18161\
        );

    \I__4118\ : InMux
    port map (
            O => \N__18175\,
            I => \N__18158\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__18172\,
            I => \N__18155\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18171\,
            I => \N__18152\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__18168\,
            I => \N__18149\
        );

    \I__4114\ : Span4Mux_h
    port map (
            O => \N__18165\,
            I => \N__18146\
        );

    \I__4113\ : InMux
    port map (
            O => \N__18164\,
            I => \N__18143\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__18161\,
            I => \N__18140\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__18158\,
            I => \N__18137\
        );

    \I__4110\ : Span4Mux_v
    port map (
            O => \N__18155\,
            I => \N__18132\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__18152\,
            I => \N__18132\
        );

    \I__4108\ : Span12Mux_s9_h
    port map (
            O => \N__18149\,
            I => \N__18128\
        );

    \I__4107\ : Sp12to4
    port map (
            O => \N__18146\,
            I => \N__18125\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__18143\,
            I => \N__18122\
        );

    \I__4105\ : Span4Mux_v
    port map (
            O => \N__18140\,
            I => \N__18119\
        );

    \I__4104\ : Span4Mux_h
    port map (
            O => \N__18137\,
            I => \N__18116\
        );

    \I__4103\ : Span4Mux_h
    port map (
            O => \N__18132\,
            I => \N__18113\
        );

    \I__4102\ : InMux
    port map (
            O => \N__18131\,
            I => \N__18110\
        );

    \I__4101\ : Span12Mux_v
    port map (
            O => \N__18128\,
            I => \N__18107\
        );

    \I__4100\ : Span12Mux_s8_v
    port map (
            O => \N__18125\,
            I => \N__18102\
        );

    \I__4099\ : Span12Mux_s9_h
    port map (
            O => \N__18122\,
            I => \N__18102\
        );

    \I__4098\ : Span4Mux_v
    port map (
            O => \N__18119\,
            I => \N__18093\
        );

    \I__4097\ : Span4Mux_v
    port map (
            O => \N__18116\,
            I => \N__18093\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__18113\,
            I => \N__18093\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__18110\,
            I => \N__18093\
        );

    \I__4094\ : Odrv12
    port map (
            O => \N__18107\,
            I => \M_this_vram_write_data_0_i_1\
        );

    \I__4093\ : Odrv12
    port map (
            O => \N__18102\,
            I => \M_this_vram_write_data_0_i_1\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__18093\,
            I => \M_this_vram_write_data_0_i_1\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__18086\,
            I => \N__18077\
        );

    \I__4090\ : CascadeMux
    port map (
            O => \N__18085\,
            I => \N__18074\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__18084\,
            I => \N__18070\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__18083\,
            I => \N__18066\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__18082\,
            I => \N__18063\
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__18081\,
            I => \N__18060\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__18080\,
            I => \N__18057\
        );

    \I__4084\ : InMux
    port map (
            O => \N__18077\,
            I => \N__18052\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18052\
        );

    \I__4082\ : CascadeMux
    port map (
            O => \N__18073\,
            I => \N__18047\
        );

    \I__4081\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18042\
        );

    \I__4080\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18035\
        );

    \I__4079\ : InMux
    port map (
            O => \N__18066\,
            I => \N__18035\
        );

    \I__4078\ : InMux
    port map (
            O => \N__18063\,
            I => \N__18035\
        );

    \I__4077\ : InMux
    port map (
            O => \N__18060\,
            I => \N__18032\
        );

    \I__4076\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18029\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__18052\,
            I => \N__18026\
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__18051\,
            I => \N__18023\
        );

    \I__4073\ : InMux
    port map (
            O => \N__18050\,
            I => \N__18014\
        );

    \I__4072\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18014\
        );

    \I__4071\ : InMux
    port map (
            O => \N__18046\,
            I => \N__18014\
        );

    \I__4070\ : InMux
    port map (
            O => \N__18045\,
            I => \N__18014\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__18042\,
            I => \N__18008\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__18035\,
            I => \N__18008\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__18032\,
            I => \N__18001\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__18029\,
            I => \N__18001\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__18026\,
            I => \N__18001\
        );

    \I__4064\ : InMux
    port map (
            O => \N__18023\,
            I => \N__17998\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__18014\,
            I => \N__17995\
        );

    \I__4062\ : InMux
    port map (
            O => \N__18013\,
            I => \N__17992\
        );

    \I__4061\ : Span4Mux_h
    port map (
            O => \N__18008\,
            I => \N__17989\
        );

    \I__4060\ : Span4Mux_v
    port map (
            O => \N__18001\,
            I => \N__17986\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__17998\,
            I => \N__17981\
        );

    \I__4058\ : Span12Mux_h
    port map (
            O => \N__17995\,
            I => \N__17981\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__17992\,
            I => \M_this_internal_address_q_3_sm0_0\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__17989\,
            I => \M_this_internal_address_q_3_sm0_0\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__17986\,
            I => \M_this_internal_address_q_3_sm0_0\
        );

    \I__4054\ : Odrv12
    port map (
            O => \N__17981\,
            I => \M_this_internal_address_q_3_sm0_0\
        );

    \I__4053\ : InMux
    port map (
            O => \N__17972\,
            I => \N__17969\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__17969\,
            I => \N__17966\
        );

    \I__4051\ : Odrv4
    port map (
            O => \N__17966\,
            I => \this_vram.mem_out_bus4_1\
        );

    \I__4050\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17960\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__17960\,
            I => \N__17957\
        );

    \I__4048\ : Span12Mux_h
    port map (
            O => \N__17957\,
            I => \N__17954\
        );

    \I__4047\ : Span12Mux_v
    port map (
            O => \N__17954\,
            I => \N__17951\
        );

    \I__4046\ : Odrv12
    port map (
            O => \N__17951\,
            I => \this_vram.mem_out_bus0_1\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__17948\,
            I => \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_\
        );

    \I__4044\ : InMux
    port map (
            O => \N__17945\,
            I => \N__17942\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__17942\,
            I => \N__17939\
        );

    \I__4042\ : Odrv12
    port map (
            O => \N__17939\,
            I => \M_this_vga_signals_address_11\
        );

    \I__4041\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17933\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__17933\,
            I => \this_vram.mem_DOUT_7_i_m2_ns_1_1\
        );

    \I__4039\ : CascadeMux
    port map (
            O => \N__17930\,
            I => \N__17927\
        );

    \I__4038\ : InMux
    port map (
            O => \N__17927\,
            I => \N__17915\
        );

    \I__4037\ : InMux
    port map (
            O => \N__17926\,
            I => \N__17915\
        );

    \I__4036\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17915\
        );

    \I__4035\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17912\
        );

    \I__4034\ : InMux
    port map (
            O => \N__17923\,
            I => \N__17907\
        );

    \I__4033\ : InMux
    port map (
            O => \N__17922\,
            I => \N__17907\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__17915\,
            I => \N__17904\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__17912\,
            I => \N__17899\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__17907\,
            I => \N__17899\
        );

    \I__4029\ : Span4Mux_v
    port map (
            O => \N__17904\,
            I => \N__17896\
        );

    \I__4028\ : Span4Mux_v
    port map (
            O => \N__17899\,
            I => \N__17893\
        );

    \I__4027\ : Span4Mux_h
    port map (
            O => \N__17896\,
            I => \N__17890\
        );

    \I__4026\ : Sp12to4
    port map (
            O => \N__17893\,
            I => \N__17885\
        );

    \I__4025\ : Sp12to4
    port map (
            O => \N__17890\,
            I => \N__17885\
        );

    \I__4024\ : Span12Mux_h
    port map (
            O => \N__17885\,
            I => \N__17882\
        );

    \I__4023\ : Odrv12
    port map (
            O => \N__17882\,
            I => \M_this_vram_read_data_1\
        );

    \I__4022\ : CascadeMux
    port map (
            O => \N__17879\,
            I => \N__17876\
        );

    \I__4021\ : CascadeBuf
    port map (
            O => \N__17876\,
            I => \N__17873\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__17873\,
            I => \N__17870\
        );

    \I__4019\ : CascadeBuf
    port map (
            O => \N__17870\,
            I => \N__17867\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__17867\,
            I => \N__17864\
        );

    \I__4017\ : CascadeBuf
    port map (
            O => \N__17864\,
            I => \N__17861\
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__17861\,
            I => \N__17858\
        );

    \I__4015\ : CascadeBuf
    port map (
            O => \N__17858\,
            I => \N__17855\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__17855\,
            I => \N__17852\
        );

    \I__4013\ : CascadeBuf
    port map (
            O => \N__17852\,
            I => \N__17849\
        );

    \I__4012\ : CascadeMux
    port map (
            O => \N__17849\,
            I => \N__17846\
        );

    \I__4011\ : CascadeBuf
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__17843\,
            I => \N__17840\
        );

    \I__4009\ : CascadeBuf
    port map (
            O => \N__17840\,
            I => \N__17837\
        );

    \I__4008\ : CascadeMux
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__4007\ : CascadeBuf
    port map (
            O => \N__17834\,
            I => \N__17831\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__17831\,
            I => \N__17828\
        );

    \I__4005\ : CascadeBuf
    port map (
            O => \N__17828\,
            I => \N__17825\
        );

    \I__4004\ : CascadeMux
    port map (
            O => \N__17825\,
            I => \N__17822\
        );

    \I__4003\ : CascadeBuf
    port map (
            O => \N__17822\,
            I => \N__17819\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__17819\,
            I => \N__17816\
        );

    \I__4001\ : CascadeBuf
    port map (
            O => \N__17816\,
            I => \N__17813\
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__17813\,
            I => \N__17810\
        );

    \I__3999\ : CascadeBuf
    port map (
            O => \N__17810\,
            I => \N__17807\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__17807\,
            I => \N__17804\
        );

    \I__3997\ : CascadeBuf
    port map (
            O => \N__17804\,
            I => \N__17801\
        );

    \I__3996\ : CascadeMux
    port map (
            O => \N__17801\,
            I => \N__17798\
        );

    \I__3995\ : CascadeBuf
    port map (
            O => \N__17798\,
            I => \N__17795\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__3993\ : CascadeBuf
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__17789\,
            I => \N__17786\
        );

    \I__3991\ : InMux
    port map (
            O => \N__17786\,
            I => \N__17783\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__17783\,
            I => \N__17780\
        );

    \I__3989\ : Span4Mux_v
    port map (
            O => \N__17780\,
            I => \N__17777\
        );

    \I__3988\ : Span4Mux_h
    port map (
            O => \N__17777\,
            I => \N__17772\
        );

    \I__3987\ : InMux
    port map (
            O => \N__17776\,
            I => \N__17769\
        );

    \I__3986\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17766\
        );

    \I__3985\ : Span4Mux_v
    port map (
            O => \N__17772\,
            I => \N__17763\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__17769\,
            I => \M_this_internal_address_qZ0Z_6\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__17766\,
            I => \M_this_internal_address_qZ0Z_6\
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__17763\,
            I => \M_this_internal_address_qZ0Z_6\
        );

    \I__3981\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17753\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__17753\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_6\
        );

    \I__3979\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17742\
        );

    \I__3978\ : InMux
    port map (
            O => \N__17749\,
            I => \N__17738\
        );

    \I__3977\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17727\
        );

    \I__3976\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17727\
        );

    \I__3975\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17727\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__17745\,
            I => \N__17723\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__17742\,
            I => \N__17716\
        );

    \I__3972\ : InMux
    port map (
            O => \N__17741\,
            I => \N__17713\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__17738\,
            I => \N__17710\
        );

    \I__3970\ : InMux
    port map (
            O => \N__17737\,
            I => \N__17707\
        );

    \I__3969\ : InMux
    port map (
            O => \N__17736\,
            I => \N__17700\
        );

    \I__3968\ : InMux
    port map (
            O => \N__17735\,
            I => \N__17700\
        );

    \I__3967\ : InMux
    port map (
            O => \N__17734\,
            I => \N__17700\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__17727\,
            I => \N__17697\
        );

    \I__3965\ : InMux
    port map (
            O => \N__17726\,
            I => \N__17694\
        );

    \I__3964\ : InMux
    port map (
            O => \N__17723\,
            I => \N__17691\
        );

    \I__3963\ : InMux
    port map (
            O => \N__17722\,
            I => \N__17688\
        );

    \I__3962\ : InMux
    port map (
            O => \N__17721\,
            I => \N__17685\
        );

    \I__3961\ : InMux
    port map (
            O => \N__17720\,
            I => \N__17680\
        );

    \I__3960\ : InMux
    port map (
            O => \N__17719\,
            I => \N__17680\
        );

    \I__3959\ : Span4Mux_v
    port map (
            O => \N__17716\,
            I => \N__17677\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__17713\,
            I => \N__17674\
        );

    \I__3957\ : Span4Mux_h
    port map (
            O => \N__17710\,
            I => \N__17671\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__17707\,
            I => \N__17666\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__17700\,
            I => \N__17666\
        );

    \I__3954\ : Span4Mux_v
    port map (
            O => \N__17697\,
            I => \N__17661\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__17694\,
            I => \N__17661\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__17691\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__17688\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__17685\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__17680\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3948\ : Odrv4
    port map (
            O => \N__17677\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__17674\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__17671\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__17666\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__17661\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__17642\,
            I => \N__17639\
        );

    \I__3942\ : CascadeBuf
    port map (
            O => \N__17639\,
            I => \N__17636\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__17636\,
            I => \N__17633\
        );

    \I__3940\ : CascadeBuf
    port map (
            O => \N__17633\,
            I => \N__17630\
        );

    \I__3939\ : CascadeMux
    port map (
            O => \N__17630\,
            I => \N__17627\
        );

    \I__3938\ : CascadeBuf
    port map (
            O => \N__17627\,
            I => \N__17624\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__17624\,
            I => \N__17621\
        );

    \I__3936\ : CascadeBuf
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__17618\,
            I => \N__17615\
        );

    \I__3934\ : CascadeBuf
    port map (
            O => \N__17615\,
            I => \N__17612\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__17612\,
            I => \N__17609\
        );

    \I__3932\ : CascadeBuf
    port map (
            O => \N__17609\,
            I => \N__17606\
        );

    \I__3931\ : CascadeMux
    port map (
            O => \N__17606\,
            I => \N__17603\
        );

    \I__3930\ : CascadeBuf
    port map (
            O => \N__17603\,
            I => \N__17600\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__17600\,
            I => \N__17597\
        );

    \I__3928\ : CascadeBuf
    port map (
            O => \N__17597\,
            I => \N__17594\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__17594\,
            I => \N__17591\
        );

    \I__3926\ : CascadeBuf
    port map (
            O => \N__17591\,
            I => \N__17588\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__17588\,
            I => \N__17585\
        );

    \I__3924\ : CascadeBuf
    port map (
            O => \N__17585\,
            I => \N__17582\
        );

    \I__3923\ : CascadeMux
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__3922\ : CascadeBuf
    port map (
            O => \N__17579\,
            I => \N__17576\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__3920\ : CascadeBuf
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__3919\ : CascadeMux
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__3918\ : CascadeBuf
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__3916\ : CascadeBuf
    port map (
            O => \N__17561\,
            I => \N__17558\
        );

    \I__3915\ : CascadeMux
    port map (
            O => \N__17558\,
            I => \N__17555\
        );

    \I__3914\ : CascadeBuf
    port map (
            O => \N__17555\,
            I => \N__17552\
        );

    \I__3913\ : CascadeMux
    port map (
            O => \N__17552\,
            I => \N__17549\
        );

    \I__3912\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17546\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__3910\ : Span4Mux_s2_v
    port map (
            O => \N__17543\,
            I => \N__17540\
        );

    \I__3909\ : Span4Mux_v
    port map (
            O => \N__17540\,
            I => \N__17535\
        );

    \I__3908\ : InMux
    port map (
            O => \N__17539\,
            I => \N__17532\
        );

    \I__3907\ : InMux
    port map (
            O => \N__17538\,
            I => \N__17529\
        );

    \I__3906\ : Span4Mux_v
    port map (
            O => \N__17535\,
            I => \N__17526\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__17532\,
            I => \M_this_internal_address_qZ0Z_8\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__17529\,
            I => \M_this_internal_address_qZ0Z_8\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__17526\,
            I => \M_this_internal_address_qZ0Z_8\
        );

    \I__3902\ : InMux
    port map (
            O => \N__17519\,
            I => \N__17516\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__17516\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_8\
        );

    \I__3900\ : InMux
    port map (
            O => \N__17513\,
            I => \N__17510\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__17510\,
            I => \N__17507\
        );

    \I__3898\ : Span12Mux_h
    port map (
            O => \N__17507\,
            I => \N__17504\
        );

    \I__3897\ : Odrv12
    port map (
            O => \N__17504\,
            I => port_address_in_3
        );

    \I__3896\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17498\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__17498\,
            I => \N__17495\
        );

    \I__3894\ : Odrv12
    port map (
            O => \N__17495\,
            I => port_address_in_2
        );

    \I__3893\ : InMux
    port map (
            O => \N__17492\,
            I => \N__17480\
        );

    \I__3892\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17480\
        );

    \I__3891\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17480\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17480\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__17480\,
            I => \N__17477\
        );

    \I__3888\ : Span4Mux_v
    port map (
            O => \N__17477\,
            I => \N__17474\
        );

    \I__3887\ : Odrv4
    port map (
            O => \N__17474\,
            I => \this_start_data_delay.M_this_state_d27Z0Z_2\
        );

    \I__3886\ : InMux
    port map (
            O => \N__17471\,
            I => \N__17468\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__17468\,
            I => \N__17465\
        );

    \I__3884\ : Span4Mux_h
    port map (
            O => \N__17465\,
            I => \N__17462\
        );

    \I__3883\ : Odrv4
    port map (
            O => \N__17462\,
            I => \un1_M_this_internal_address_q_cry_10_c_RNI6I0DZ0\
        );

    \I__3882\ : InMux
    port map (
            O => \N__17459\,
            I => \un1_M_this_internal_address_q_cry_10\
        );

    \I__3881\ : InMux
    port map (
            O => \N__17456\,
            I => \un1_M_this_internal_address_q_cry_11\
        );

    \I__3880\ : InMux
    port map (
            O => \N__17453\,
            I => \un1_M_this_internal_address_q_cry_12\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__17450\,
            I => \N__17447\
        );

    \I__3878\ : CascadeBuf
    port map (
            O => \N__17447\,
            I => \N__17444\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__17444\,
            I => \N__17441\
        );

    \I__3876\ : CascadeBuf
    port map (
            O => \N__17441\,
            I => \N__17438\
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__17438\,
            I => \N__17435\
        );

    \I__3874\ : CascadeBuf
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__17432\,
            I => \N__17429\
        );

    \I__3872\ : CascadeBuf
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__3871\ : CascadeMux
    port map (
            O => \N__17426\,
            I => \N__17423\
        );

    \I__3870\ : CascadeBuf
    port map (
            O => \N__17423\,
            I => \N__17420\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__17420\,
            I => \N__17417\
        );

    \I__3868\ : CascadeBuf
    port map (
            O => \N__17417\,
            I => \N__17414\
        );

    \I__3867\ : CascadeMux
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__3866\ : CascadeBuf
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__3865\ : CascadeMux
    port map (
            O => \N__17408\,
            I => \N__17405\
        );

    \I__3864\ : CascadeBuf
    port map (
            O => \N__17405\,
            I => \N__17402\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__17402\,
            I => \N__17399\
        );

    \I__3862\ : CascadeBuf
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__17396\,
            I => \N__17393\
        );

    \I__3860\ : CascadeBuf
    port map (
            O => \N__17393\,
            I => \N__17390\
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__17390\,
            I => \N__17387\
        );

    \I__3858\ : CascadeBuf
    port map (
            O => \N__17387\,
            I => \N__17384\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__17384\,
            I => \N__17381\
        );

    \I__3856\ : CascadeBuf
    port map (
            O => \N__17381\,
            I => \N__17378\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__17378\,
            I => \N__17375\
        );

    \I__3854\ : CascadeBuf
    port map (
            O => \N__17375\,
            I => \N__17372\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__17372\,
            I => \N__17369\
        );

    \I__3852\ : CascadeBuf
    port map (
            O => \N__17369\,
            I => \N__17366\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__17366\,
            I => \N__17363\
        );

    \I__3850\ : CascadeBuf
    port map (
            O => \N__17363\,
            I => \N__17360\
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__17360\,
            I => \N__17357\
        );

    \I__3848\ : InMux
    port map (
            O => \N__17357\,
            I => \N__17353\
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__17356\,
            I => \N__17350\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__17353\,
            I => \N__17347\
        );

    \I__3845\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17344\
        );

    \I__3844\ : Span12Mux_h
    port map (
            O => \N__17347\,
            I => \N__17340\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17344\,
            I => \N__17337\
        );

    \I__3842\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17334\
        );

    \I__3841\ : Span12Mux_v
    port map (
            O => \N__17340\,
            I => \N__17331\
        );

    \I__3840\ : Odrv4
    port map (
            O => \N__17337\,
            I => \M_this_internal_address_qZ0Z_0\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__17334\,
            I => \M_this_internal_address_qZ0Z_0\
        );

    \I__3838\ : Odrv12
    port map (
            O => \N__17331\,
            I => \M_this_internal_address_qZ0Z_0\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__17324\,
            I => \N__17321\
        );

    \I__3836\ : InMux
    port map (
            O => \N__17321\,
            I => \N__17318\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__17318\,
            I => \N__17315\
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__17315\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_0\
        );

    \I__3833\ : InMux
    port map (
            O => \N__17312\,
            I => \N__17309\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__17309\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_10\
        );

    \I__3831\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17303\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__17303\,
            I => \un1_M_this_internal_address_q_cry_9_c_RNITQCIZ0\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__17300\,
            I => \N__17297\
        );

    \I__3828\ : CascadeBuf
    port map (
            O => \N__17297\,
            I => \N__17294\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__17294\,
            I => \N__17291\
        );

    \I__3826\ : CascadeBuf
    port map (
            O => \N__17291\,
            I => \N__17288\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__17288\,
            I => \N__17285\
        );

    \I__3824\ : CascadeBuf
    port map (
            O => \N__17285\,
            I => \N__17282\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__17282\,
            I => \N__17279\
        );

    \I__3822\ : CascadeBuf
    port map (
            O => \N__17279\,
            I => \N__17276\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__17276\,
            I => \N__17273\
        );

    \I__3820\ : CascadeBuf
    port map (
            O => \N__17273\,
            I => \N__17270\
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__17270\,
            I => \N__17267\
        );

    \I__3818\ : CascadeBuf
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__17264\,
            I => \N__17261\
        );

    \I__3816\ : CascadeBuf
    port map (
            O => \N__17261\,
            I => \N__17258\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__17258\,
            I => \N__17255\
        );

    \I__3814\ : CascadeBuf
    port map (
            O => \N__17255\,
            I => \N__17252\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__17252\,
            I => \N__17249\
        );

    \I__3812\ : CascadeBuf
    port map (
            O => \N__17249\,
            I => \N__17246\
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__17246\,
            I => \N__17243\
        );

    \I__3810\ : CascadeBuf
    port map (
            O => \N__17243\,
            I => \N__17240\
        );

    \I__3809\ : CascadeMux
    port map (
            O => \N__17240\,
            I => \N__17237\
        );

    \I__3808\ : CascadeBuf
    port map (
            O => \N__17237\,
            I => \N__17234\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__17234\,
            I => \N__17231\
        );

    \I__3806\ : CascadeBuf
    port map (
            O => \N__17231\,
            I => \N__17228\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__17228\,
            I => \N__17225\
        );

    \I__3804\ : CascadeBuf
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__17222\,
            I => \N__17219\
        );

    \I__3802\ : CascadeBuf
    port map (
            O => \N__17219\,
            I => \N__17216\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__17216\,
            I => \N__17213\
        );

    \I__3800\ : CascadeBuf
    port map (
            O => \N__17213\,
            I => \N__17210\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__17210\,
            I => \N__17207\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17204\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__17204\,
            I => \N__17201\
        );

    \I__3796\ : Span4Mux_s2_v
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__3795\ : Span4Mux_h
    port map (
            O => \N__17198\,
            I => \N__17193\
        );

    \I__3794\ : InMux
    port map (
            O => \N__17197\,
            I => \N__17190\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17196\,
            I => \N__17187\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__17193\,
            I => \N__17184\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__17190\,
            I => \M_this_internal_address_qZ0Z_10\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__17187\,
            I => \M_this_internal_address_qZ0Z_10\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__17184\,
            I => \M_this_internal_address_qZ0Z_10\
        );

    \I__3788\ : InMux
    port map (
            O => \N__17177\,
            I => \N__17174\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__17174\,
            I => \N__17171\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__17171\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_12\
        );

    \I__3785\ : InMux
    port map (
            O => \N__17168\,
            I => \N__17165\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__17165\,
            I => \un1_M_this_internal_address_q_cry_11_c_RNI8L1DZ0\
        );

    \I__3783\ : InMux
    port map (
            O => \N__17162\,
            I => \N__17159\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__17159\,
            I => \un1_M_this_internal_address_q_cry_5_c_RNIE50JZ0\
        );

    \I__3781\ : InMux
    port map (
            O => \N__17156\,
            I => \N__17153\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__17153\,
            I => \N__17150\
        );

    \I__3779\ : Span4Mux_h
    port map (
            O => \N__17150\,
            I => \N__17147\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__17147\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_13\
        );

    \I__3777\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17141\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__17141\,
            I => \un1_M_this_internal_address_q_cry_12_c_RNIAO2DZ0\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17138\,
            I => \N__17135\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__17135\,
            I => \un1_M_this_internal_address_q_cry_7_c_RNIIB2JZ0\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__17132\,
            I => \N__17129\
        );

    \I__3772\ : CascadeBuf
    port map (
            O => \N__17129\,
            I => \N__17126\
        );

    \I__3771\ : CascadeMux
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__3770\ : CascadeBuf
    port map (
            O => \N__17123\,
            I => \N__17120\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__17120\,
            I => \N__17117\
        );

    \I__3768\ : CascadeBuf
    port map (
            O => \N__17117\,
            I => \N__17114\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__17114\,
            I => \N__17111\
        );

    \I__3766\ : CascadeBuf
    port map (
            O => \N__17111\,
            I => \N__17108\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__17108\,
            I => \N__17105\
        );

    \I__3764\ : CascadeBuf
    port map (
            O => \N__17105\,
            I => \N__17102\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__17102\,
            I => \N__17099\
        );

    \I__3762\ : CascadeBuf
    port map (
            O => \N__17099\,
            I => \N__17096\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__17096\,
            I => \N__17093\
        );

    \I__3760\ : CascadeBuf
    port map (
            O => \N__17093\,
            I => \N__17090\
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__17090\,
            I => \N__17087\
        );

    \I__3758\ : CascadeBuf
    port map (
            O => \N__17087\,
            I => \N__17084\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__17084\,
            I => \N__17081\
        );

    \I__3756\ : CascadeBuf
    port map (
            O => \N__17081\,
            I => \N__17078\
        );

    \I__3755\ : CascadeMux
    port map (
            O => \N__17078\,
            I => \N__17075\
        );

    \I__3754\ : CascadeBuf
    port map (
            O => \N__17075\,
            I => \N__17072\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__17072\,
            I => \N__17069\
        );

    \I__3752\ : CascadeBuf
    port map (
            O => \N__17069\,
            I => \N__17066\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__17066\,
            I => \N__17063\
        );

    \I__3750\ : CascadeBuf
    port map (
            O => \N__17063\,
            I => \N__17060\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__17060\,
            I => \N__17057\
        );

    \I__3748\ : CascadeBuf
    port map (
            O => \N__17057\,
            I => \N__17054\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__17054\,
            I => \N__17051\
        );

    \I__3746\ : CascadeBuf
    port map (
            O => \N__17051\,
            I => \N__17048\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__17048\,
            I => \N__17045\
        );

    \I__3744\ : CascadeBuf
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__3742\ : InMux
    port map (
            O => \N__17039\,
            I => \N__17036\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__17036\,
            I => \N__17032\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17035\,
            I => \N__17028\
        );

    \I__3739\ : Span12Mux_h
    port map (
            O => \N__17032\,
            I => \N__17025\
        );

    \I__3738\ : InMux
    port map (
            O => \N__17031\,
            I => \N__17022\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__17028\,
            I => \N__17017\
        );

    \I__3736\ : Span12Mux_v
    port map (
            O => \N__17025\,
            I => \N__17017\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__17022\,
            I => \M_this_internal_address_qZ0Z_3\
        );

    \I__3734\ : Odrv12
    port map (
            O => \N__17017\,
            I => \M_this_internal_address_qZ0Z_3\
        );

    \I__3733\ : CascadeMux
    port map (
            O => \N__17012\,
            I => \N__17009\
        );

    \I__3732\ : InMux
    port map (
            O => \N__17009\,
            I => \N__17006\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__17006\,
            I => \un1_M_this_internal_address_q_cry_2_c_RNI8SSIZ0\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17003\,
            I => \un1_M_this_internal_address_q_cry_2\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__17000\,
            I => \N__16997\
        );

    \I__3728\ : CascadeBuf
    port map (
            O => \N__16997\,
            I => \N__16994\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__16994\,
            I => \N__16991\
        );

    \I__3726\ : CascadeBuf
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__16988\,
            I => \N__16985\
        );

    \I__3724\ : CascadeBuf
    port map (
            O => \N__16985\,
            I => \N__16982\
        );

    \I__3723\ : CascadeMux
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__3722\ : CascadeBuf
    port map (
            O => \N__16979\,
            I => \N__16976\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__16976\,
            I => \N__16973\
        );

    \I__3720\ : CascadeBuf
    port map (
            O => \N__16973\,
            I => \N__16970\
        );

    \I__3719\ : CascadeMux
    port map (
            O => \N__16970\,
            I => \N__16967\
        );

    \I__3718\ : CascadeBuf
    port map (
            O => \N__16967\,
            I => \N__16964\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__16964\,
            I => \N__16961\
        );

    \I__3716\ : CascadeBuf
    port map (
            O => \N__16961\,
            I => \N__16958\
        );

    \I__3715\ : CascadeMux
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__3714\ : CascadeBuf
    port map (
            O => \N__16955\,
            I => \N__16952\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__16952\,
            I => \N__16949\
        );

    \I__3712\ : CascadeBuf
    port map (
            O => \N__16949\,
            I => \N__16946\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__16946\,
            I => \N__16943\
        );

    \I__3710\ : CascadeBuf
    port map (
            O => \N__16943\,
            I => \N__16940\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__16940\,
            I => \N__16937\
        );

    \I__3708\ : CascadeBuf
    port map (
            O => \N__16937\,
            I => \N__16934\
        );

    \I__3707\ : CascadeMux
    port map (
            O => \N__16934\,
            I => \N__16931\
        );

    \I__3706\ : CascadeBuf
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__16928\,
            I => \N__16925\
        );

    \I__3704\ : CascadeBuf
    port map (
            O => \N__16925\,
            I => \N__16922\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__16922\,
            I => \N__16919\
        );

    \I__3702\ : CascadeBuf
    port map (
            O => \N__16919\,
            I => \N__16916\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__3700\ : CascadeBuf
    port map (
            O => \N__16913\,
            I => \N__16910\
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__16910\,
            I => \N__16907\
        );

    \I__3698\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16904\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__16904\,
            I => \N__16901\
        );

    \I__3696\ : Span4Mux_h
    port map (
            O => \N__16901\,
            I => \N__16898\
        );

    \I__3695\ : Span4Mux_h
    port map (
            O => \N__16898\,
            I => \N__16893\
        );

    \I__3694\ : InMux
    port map (
            O => \N__16897\,
            I => \N__16890\
        );

    \I__3693\ : InMux
    port map (
            O => \N__16896\,
            I => \N__16887\
        );

    \I__3692\ : Sp12to4
    port map (
            O => \N__16893\,
            I => \N__16884\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__16890\,
            I => \M_this_internal_address_qZ0Z_4\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__16887\,
            I => \M_this_internal_address_qZ0Z_4\
        );

    \I__3689\ : Odrv12
    port map (
            O => \N__16884\,
            I => \M_this_internal_address_qZ0Z_4\
        );

    \I__3688\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16874\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__16874\,
            I => \un1_M_this_internal_address_q_cry_3_c_RNIAVTIZ0\
        );

    \I__3686\ : InMux
    port map (
            O => \N__16871\,
            I => \un1_M_this_internal_address_q_cry_3\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__16868\,
            I => \N__16865\
        );

    \I__3684\ : CascadeBuf
    port map (
            O => \N__16865\,
            I => \N__16862\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__16862\,
            I => \N__16859\
        );

    \I__3682\ : CascadeBuf
    port map (
            O => \N__16859\,
            I => \N__16856\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__16856\,
            I => \N__16853\
        );

    \I__3680\ : CascadeBuf
    port map (
            O => \N__16853\,
            I => \N__16850\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__16850\,
            I => \N__16847\
        );

    \I__3678\ : CascadeBuf
    port map (
            O => \N__16847\,
            I => \N__16844\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__16844\,
            I => \N__16841\
        );

    \I__3676\ : CascadeBuf
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__3674\ : CascadeBuf
    port map (
            O => \N__16835\,
            I => \N__16832\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__16832\,
            I => \N__16829\
        );

    \I__3672\ : CascadeBuf
    port map (
            O => \N__16829\,
            I => \N__16826\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__16826\,
            I => \N__16823\
        );

    \I__3670\ : CascadeBuf
    port map (
            O => \N__16823\,
            I => \N__16820\
        );

    \I__3669\ : CascadeMux
    port map (
            O => \N__16820\,
            I => \N__16817\
        );

    \I__3668\ : CascadeBuf
    port map (
            O => \N__16817\,
            I => \N__16814\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__16814\,
            I => \N__16811\
        );

    \I__3666\ : CascadeBuf
    port map (
            O => \N__16811\,
            I => \N__16808\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__16808\,
            I => \N__16805\
        );

    \I__3664\ : CascadeBuf
    port map (
            O => \N__16805\,
            I => \N__16802\
        );

    \I__3663\ : CascadeMux
    port map (
            O => \N__16802\,
            I => \N__16799\
        );

    \I__3662\ : CascadeBuf
    port map (
            O => \N__16799\,
            I => \N__16796\
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__16796\,
            I => \N__16793\
        );

    \I__3660\ : CascadeBuf
    port map (
            O => \N__16793\,
            I => \N__16790\
        );

    \I__3659\ : CascadeMux
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__3658\ : CascadeBuf
    port map (
            O => \N__16787\,
            I => \N__16784\
        );

    \I__3657\ : CascadeMux
    port map (
            O => \N__16784\,
            I => \N__16781\
        );

    \I__3656\ : CascadeBuf
    port map (
            O => \N__16781\,
            I => \N__16778\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__16778\,
            I => \N__16775\
        );

    \I__3654\ : InMux
    port map (
            O => \N__16775\,
            I => \N__16772\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__16772\,
            I => \N__16769\
        );

    \I__3652\ : Span4Mux_s2_v
    port map (
            O => \N__16769\,
            I => \N__16766\
        );

    \I__3651\ : Sp12to4
    port map (
            O => \N__16766\,
            I => \N__16761\
        );

    \I__3650\ : InMux
    port map (
            O => \N__16765\,
            I => \N__16758\
        );

    \I__3649\ : InMux
    port map (
            O => \N__16764\,
            I => \N__16755\
        );

    \I__3648\ : Span12Mux_h
    port map (
            O => \N__16761\,
            I => \N__16752\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__16758\,
            I => \M_this_internal_address_qZ0Z_5\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__16755\,
            I => \M_this_internal_address_qZ0Z_5\
        );

    \I__3645\ : Odrv12
    port map (
            O => \N__16752\,
            I => \M_this_internal_address_qZ0Z_5\
        );

    \I__3644\ : InMux
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__16742\,
            I => \un1_M_this_internal_address_q_cry_4_c_RNIC2VIZ0\
        );

    \I__3642\ : InMux
    port map (
            O => \N__16739\,
            I => \un1_M_this_internal_address_q_cry_4\
        );

    \I__3641\ : InMux
    port map (
            O => \N__16736\,
            I => \un1_M_this_internal_address_q_cry_5\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__16733\,
            I => \N__16730\
        );

    \I__3639\ : CascadeBuf
    port map (
            O => \N__16730\,
            I => \N__16727\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__16727\,
            I => \N__16724\
        );

    \I__3637\ : CascadeBuf
    port map (
            O => \N__16724\,
            I => \N__16721\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__16721\,
            I => \N__16718\
        );

    \I__3635\ : CascadeBuf
    port map (
            O => \N__16718\,
            I => \N__16715\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__16715\,
            I => \N__16712\
        );

    \I__3633\ : CascadeBuf
    port map (
            O => \N__16712\,
            I => \N__16709\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__16709\,
            I => \N__16706\
        );

    \I__3631\ : CascadeBuf
    port map (
            O => \N__16706\,
            I => \N__16703\
        );

    \I__3630\ : CascadeMux
    port map (
            O => \N__16703\,
            I => \N__16700\
        );

    \I__3629\ : CascadeBuf
    port map (
            O => \N__16700\,
            I => \N__16697\
        );

    \I__3628\ : CascadeMux
    port map (
            O => \N__16697\,
            I => \N__16694\
        );

    \I__3627\ : CascadeBuf
    port map (
            O => \N__16694\,
            I => \N__16691\
        );

    \I__3626\ : CascadeMux
    port map (
            O => \N__16691\,
            I => \N__16688\
        );

    \I__3625\ : CascadeBuf
    port map (
            O => \N__16688\,
            I => \N__16685\
        );

    \I__3624\ : CascadeMux
    port map (
            O => \N__16685\,
            I => \N__16682\
        );

    \I__3623\ : CascadeBuf
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__16679\,
            I => \N__16676\
        );

    \I__3621\ : CascadeBuf
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__3620\ : CascadeMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__3619\ : CascadeBuf
    port map (
            O => \N__16670\,
            I => \N__16667\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__3617\ : CascadeBuf
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__3615\ : CascadeBuf
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__3613\ : CascadeBuf
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3611\ : CascadeBuf
    port map (
            O => \N__16646\,
            I => \N__16643\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__16643\,
            I => \N__16640\
        );

    \I__3609\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16637\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__16637\,
            I => \N__16634\
        );

    \I__3607\ : Span12Mux_s10_h
    port map (
            O => \N__16634\,
            I => \N__16629\
        );

    \I__3606\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16626\
        );

    \I__3605\ : InMux
    port map (
            O => \N__16632\,
            I => \N__16623\
        );

    \I__3604\ : Span12Mux_v
    port map (
            O => \N__16629\,
            I => \N__16620\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__16626\,
            I => \M_this_internal_address_qZ0Z_7\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__16623\,
            I => \M_this_internal_address_qZ0Z_7\
        );

    \I__3601\ : Odrv12
    port map (
            O => \N__16620\,
            I => \M_this_internal_address_qZ0Z_7\
        );

    \I__3600\ : InMux
    port map (
            O => \N__16613\,
            I => \N__16610\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__16610\,
            I => \un1_M_this_internal_address_q_cry_6_c_RNIG81JZ0\
        );

    \I__3598\ : InMux
    port map (
            O => \N__16607\,
            I => \un1_M_this_internal_address_q_cry_6\
        );

    \I__3597\ : InMux
    port map (
            O => \N__16604\,
            I => \bfn_20_22_0_\
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__16601\,
            I => \N__16598\
        );

    \I__3595\ : CascadeBuf
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__3593\ : CascadeBuf
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__16589\,
            I => \N__16586\
        );

    \I__3591\ : CascadeBuf
    port map (
            O => \N__16586\,
            I => \N__16583\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__3589\ : CascadeBuf
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__16577\,
            I => \N__16574\
        );

    \I__3587\ : CascadeBuf
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__16571\,
            I => \N__16568\
        );

    \I__3585\ : CascadeBuf
    port map (
            O => \N__16568\,
            I => \N__16565\
        );

    \I__3584\ : CascadeMux
    port map (
            O => \N__16565\,
            I => \N__16562\
        );

    \I__3583\ : CascadeBuf
    port map (
            O => \N__16562\,
            I => \N__16559\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__16559\,
            I => \N__16556\
        );

    \I__3581\ : CascadeBuf
    port map (
            O => \N__16556\,
            I => \N__16553\
        );

    \I__3580\ : CascadeMux
    port map (
            O => \N__16553\,
            I => \N__16550\
        );

    \I__3579\ : CascadeBuf
    port map (
            O => \N__16550\,
            I => \N__16547\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__16547\,
            I => \N__16544\
        );

    \I__3577\ : CascadeBuf
    port map (
            O => \N__16544\,
            I => \N__16541\
        );

    \I__3576\ : CascadeMux
    port map (
            O => \N__16541\,
            I => \N__16538\
        );

    \I__3575\ : CascadeBuf
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__16535\,
            I => \N__16532\
        );

    \I__3573\ : CascadeBuf
    port map (
            O => \N__16532\,
            I => \N__16529\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__16529\,
            I => \N__16526\
        );

    \I__3571\ : CascadeBuf
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__3569\ : CascadeBuf
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__3567\ : CascadeBuf
    port map (
            O => \N__16514\,
            I => \N__16511\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__16511\,
            I => \N__16508\
        );

    \I__3565\ : InMux
    port map (
            O => \N__16508\,
            I => \N__16505\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__3563\ : Span4Mux_s3_v
    port map (
            O => \N__16502\,
            I => \N__16499\
        );

    \I__3562\ : Sp12to4
    port map (
            O => \N__16499\,
            I => \N__16494\
        );

    \I__3561\ : InMux
    port map (
            O => \N__16498\,
            I => \N__16491\
        );

    \I__3560\ : InMux
    port map (
            O => \N__16497\,
            I => \N__16488\
        );

    \I__3559\ : Span12Mux_h
    port map (
            O => \N__16494\,
            I => \N__16485\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__16491\,
            I => \M_this_internal_address_qZ0Z_9\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__16488\,
            I => \M_this_internal_address_qZ0Z_9\
        );

    \I__3556\ : Odrv12
    port map (
            O => \N__16485\,
            I => \M_this_internal_address_qZ0Z_9\
        );

    \I__3555\ : InMux
    port map (
            O => \N__16478\,
            I => \N__16475\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__16475\,
            I => \un1_M_this_internal_address_q_cry_8_c_RNIKE3JZ0\
        );

    \I__3553\ : InMux
    port map (
            O => \N__16472\,
            I => \un1_M_this_internal_address_q_cry_8\
        );

    \I__3552\ : InMux
    port map (
            O => \N__16469\,
            I => \un1_M_this_internal_address_q_cry_9\
        );

    \I__3551\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__16463\,
            I => \N__16460\
        );

    \I__3549\ : Odrv12
    port map (
            O => \N__16460\,
            I => \M_this_vga_signals_address_13\
        );

    \I__3548\ : InMux
    port map (
            O => \N__16457\,
            I => \N__16454\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__16454\,
            I => \N__16451\
        );

    \I__3546\ : Sp12to4
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__3545\ : Odrv12
    port map (
            O => \N__16448\,
            I => \M_this_vga_signals_address_12\
        );

    \I__3544\ : InMux
    port map (
            O => \N__16445\,
            I => \N__16442\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__16442\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_5\
        );

    \I__3542\ : InMux
    port map (
            O => \N__16439\,
            I => \N__16436\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__16436\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_3\
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__16433\,
            I => \N__16430\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16430\,
            I => \N__16427\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__16427\,
            I => \N__16424\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__16424\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_7\
        );

    \I__3536\ : CascadeMux
    port map (
            O => \N__16421\,
            I => \N__16417\
        );

    \I__3535\ : InMux
    port map (
            O => \N__16420\,
            I => \N__16414\
        );

    \I__3534\ : InMux
    port map (
            O => \N__16417\,
            I => \N__16411\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__16414\,
            I => \N_346_0\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16411\,
            I => \N_346_0\
        );

    \I__3531\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__16403\,
            I => \M_this_internal_address_q_RNI6EA12Z0Z_0\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__16400\,
            I => \N__16397\
        );

    \I__3528\ : CascadeBuf
    port map (
            O => \N__16397\,
            I => \N__16394\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__16394\,
            I => \N__16391\
        );

    \I__3526\ : CascadeBuf
    port map (
            O => \N__16391\,
            I => \N__16388\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__16388\,
            I => \N__16385\
        );

    \I__3524\ : CascadeBuf
    port map (
            O => \N__16385\,
            I => \N__16382\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__16382\,
            I => \N__16379\
        );

    \I__3522\ : CascadeBuf
    port map (
            O => \N__16379\,
            I => \N__16376\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__16376\,
            I => \N__16373\
        );

    \I__3520\ : CascadeBuf
    port map (
            O => \N__16373\,
            I => \N__16370\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__16370\,
            I => \N__16367\
        );

    \I__3518\ : CascadeBuf
    port map (
            O => \N__16367\,
            I => \N__16364\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__16364\,
            I => \N__16361\
        );

    \I__3516\ : CascadeBuf
    port map (
            O => \N__16361\,
            I => \N__16358\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__16358\,
            I => \N__16355\
        );

    \I__3514\ : CascadeBuf
    port map (
            O => \N__16355\,
            I => \N__16352\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__16352\,
            I => \N__16349\
        );

    \I__3512\ : CascadeBuf
    port map (
            O => \N__16349\,
            I => \N__16346\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__16346\,
            I => \N__16343\
        );

    \I__3510\ : CascadeBuf
    port map (
            O => \N__16343\,
            I => \N__16340\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__16340\,
            I => \N__16337\
        );

    \I__3508\ : CascadeBuf
    port map (
            O => \N__16337\,
            I => \N__16334\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__16334\,
            I => \N__16331\
        );

    \I__3506\ : CascadeBuf
    port map (
            O => \N__16331\,
            I => \N__16328\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__16328\,
            I => \N__16325\
        );

    \I__3504\ : CascadeBuf
    port map (
            O => \N__16325\,
            I => \N__16322\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__16322\,
            I => \N__16319\
        );

    \I__3502\ : CascadeBuf
    port map (
            O => \N__16319\,
            I => \N__16316\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__16316\,
            I => \N__16313\
        );

    \I__3500\ : CascadeBuf
    port map (
            O => \N__16313\,
            I => \N__16310\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__16310\,
            I => \N__16307\
        );

    \I__3498\ : InMux
    port map (
            O => \N__16307\,
            I => \N__16304\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__16304\,
            I => \N__16300\
        );

    \I__3496\ : InMux
    port map (
            O => \N__16303\,
            I => \N__16297\
        );

    \I__3495\ : Span4Mux_s3_v
    port map (
            O => \N__16300\,
            I => \N__16294\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__16297\,
            I => \N__16291\
        );

    \I__3493\ : Span4Mux_h
    port map (
            O => \N__16294\,
            I => \N__16287\
        );

    \I__3492\ : Span4Mux_h
    port map (
            O => \N__16291\,
            I => \N__16284\
        );

    \I__3491\ : InMux
    port map (
            O => \N__16290\,
            I => \N__16281\
        );

    \I__3490\ : Span4Mux_v
    port map (
            O => \N__16287\,
            I => \N__16278\
        );

    \I__3489\ : Odrv4
    port map (
            O => \N__16284\,
            I => \M_this_internal_address_qZ0Z_1\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__16281\,
            I => \M_this_internal_address_qZ0Z_1\
        );

    \I__3487\ : Odrv4
    port map (
            O => \N__16278\,
            I => \M_this_internal_address_qZ0Z_1\
        );

    \I__3486\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16268\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__16268\,
            I => \N__16265\
        );

    \I__3484\ : Span4Mux_v
    port map (
            O => \N__16265\,
            I => \N__16262\
        );

    \I__3483\ : Odrv4
    port map (
            O => \N__16262\,
            I => \un1_M_this_internal_address_q_cry_0_c_RNI4MQIZ0\
        );

    \I__3482\ : InMux
    port map (
            O => \N__16259\,
            I => \un1_M_this_internal_address_q_cry_0\
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__16256\,
            I => \N__16253\
        );

    \I__3480\ : CascadeBuf
    port map (
            O => \N__16253\,
            I => \N__16250\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__16250\,
            I => \N__16247\
        );

    \I__3478\ : CascadeBuf
    port map (
            O => \N__16247\,
            I => \N__16244\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__16244\,
            I => \N__16241\
        );

    \I__3476\ : CascadeBuf
    port map (
            O => \N__16241\,
            I => \N__16238\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__16238\,
            I => \N__16235\
        );

    \I__3474\ : CascadeBuf
    port map (
            O => \N__16235\,
            I => \N__16232\
        );

    \I__3473\ : CascadeMux
    port map (
            O => \N__16232\,
            I => \N__16229\
        );

    \I__3472\ : CascadeBuf
    port map (
            O => \N__16229\,
            I => \N__16226\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__16226\,
            I => \N__16223\
        );

    \I__3470\ : CascadeBuf
    port map (
            O => \N__16223\,
            I => \N__16220\
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__16220\,
            I => \N__16217\
        );

    \I__3468\ : CascadeBuf
    port map (
            O => \N__16217\,
            I => \N__16214\
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__16214\,
            I => \N__16211\
        );

    \I__3466\ : CascadeBuf
    port map (
            O => \N__16211\,
            I => \N__16208\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__16208\,
            I => \N__16205\
        );

    \I__3464\ : CascadeBuf
    port map (
            O => \N__16205\,
            I => \N__16202\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__16202\,
            I => \N__16199\
        );

    \I__3462\ : CascadeBuf
    port map (
            O => \N__16199\,
            I => \N__16196\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__16196\,
            I => \N__16193\
        );

    \I__3460\ : CascadeBuf
    port map (
            O => \N__16193\,
            I => \N__16190\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__16190\,
            I => \N__16187\
        );

    \I__3458\ : CascadeBuf
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__16184\,
            I => \N__16181\
        );

    \I__3456\ : CascadeBuf
    port map (
            O => \N__16181\,
            I => \N__16178\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__16178\,
            I => \N__16175\
        );

    \I__3454\ : CascadeBuf
    port map (
            O => \N__16175\,
            I => \N__16172\
        );

    \I__3453\ : CascadeMux
    port map (
            O => \N__16172\,
            I => \N__16169\
        );

    \I__3452\ : CascadeBuf
    port map (
            O => \N__16169\,
            I => \N__16166\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__16166\,
            I => \N__16163\
        );

    \I__3450\ : InMux
    port map (
            O => \N__16163\,
            I => \N__16160\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__16160\,
            I => \N__16157\
        );

    \I__3448\ : Span4Mux_h
    port map (
            O => \N__16157\,
            I => \N__16154\
        );

    \I__3447\ : Sp12to4
    port map (
            O => \N__16154\,
            I => \N__16149\
        );

    \I__3446\ : InMux
    port map (
            O => \N__16153\,
            I => \N__16146\
        );

    \I__3445\ : InMux
    port map (
            O => \N__16152\,
            I => \N__16143\
        );

    \I__3444\ : Span12Mux_s10_v
    port map (
            O => \N__16149\,
            I => \N__16140\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__16146\,
            I => \M_this_internal_address_qZ0Z_2\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__16143\,
            I => \M_this_internal_address_qZ0Z_2\
        );

    \I__3441\ : Odrv12
    port map (
            O => \N__16140\,
            I => \M_this_internal_address_qZ0Z_2\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__16133\,
            I => \N__16130\
        );

    \I__3439\ : InMux
    port map (
            O => \N__16130\,
            I => \N__16127\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__16127\,
            I => \N__16124\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__16124\,
            I => \un1_M_this_internal_address_q_cry_1_c_RNI6PRIZ0\
        );

    \I__3436\ : InMux
    port map (
            O => \N__16121\,
            I => \un1_M_this_internal_address_q_cry_1\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16115\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__16115\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_9\
        );

    \I__3433\ : InMux
    port map (
            O => \N__16112\,
            I => \N__16109\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__16109\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_2\
        );

    \I__3431\ : InMux
    port map (
            O => \N__16106\,
            I => \N__16102\
        );

    \I__3430\ : InMux
    port map (
            O => \N__16105\,
            I => \N__16099\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__16102\,
            I => \this_start_data_delay.N_407\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__16099\,
            I => \this_start_data_delay.N_407\
        );

    \I__3427\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16087\
        );

    \I__3426\ : InMux
    port map (
            O => \N__16093\,
            I => \N__16087\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16092\,
            I => \N__16084\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__16087\,
            I => \this_start_data_delay.N_398\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__16084\,
            I => \this_start_data_delay.N_398\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16079\,
            I => \N__16076\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__16076\,
            I => \this_start_data_delay.M_this_state_dZ0Z29\
        );

    \I__3420\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16070\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__16070\,
            I => \N__16067\
        );

    \I__3418\ : Span4Mux_v
    port map (
            O => \N__16067\,
            I => \N__16064\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__16064\,
            I => \this_start_data_delay.N_396\
        );

    \I__3416\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16058\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__16058\,
            I => \this_start_data_delay.M_this_state_dZ0Z27\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__16055\,
            I => \N__16049\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__16054\,
            I => \N__16046\
        );

    \I__3412\ : InMux
    port map (
            O => \N__16053\,
            I => \N__16041\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16052\,
            I => \N__16041\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16049\,
            I => \N__16036\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16036\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__16041\,
            I => \N__16031\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__16036\,
            I => \N__16031\
        );

    \I__3406\ : Span12Mux_h
    port map (
            O => \N__16031\,
            I => \N__16028\
        );

    \I__3405\ : Odrv12
    port map (
            O => \N__16028\,
            I => port_address_in_0
        );

    \I__3404\ : InMux
    port map (
            O => \N__16025\,
            I => \N__16017\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16024\,
            I => \N__16017\
        );

    \I__3402\ : InMux
    port map (
            O => \N__16023\,
            I => \N__16012\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16012\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__16017\,
            I => \N__16007\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__16012\,
            I => \N__16007\
        );

    \I__3398\ : Span12Mux_h
    port map (
            O => \N__16007\,
            I => \N__16004\
        );

    \I__3397\ : Odrv12
    port map (
            O => \N__16004\,
            I => port_address_in_1
        );

    \I__3396\ : InMux
    port map (
            O => \N__16001\,
            I => \N__15998\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__15998\,
            I => \this_start_data_delay.M_this_state_dZ0Z28\
        );

    \I__3394\ : InMux
    port map (
            O => \N__15995\,
            I => \N__15991\
        );

    \I__3393\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15988\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__15991\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__15988\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__3390\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15980\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__15980\,
            I => \N__15972\
        );

    \I__3388\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15967\
        );

    \I__3387\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15967\
        );

    \I__3386\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15964\
        );

    \I__3385\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15959\
        );

    \I__3384\ : InMux
    port map (
            O => \N__15975\,
            I => \N__15959\
        );

    \I__3383\ : Span4Mux_v
    port map (
            O => \N__15972\,
            I => \N__15956\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__15967\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__15964\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__15959\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__15956\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__15947\,
            I => \N__15942\
        );

    \I__3377\ : InMux
    port map (
            O => \N__15946\,
            I => \N__15939\
        );

    \I__3376\ : InMux
    port map (
            O => \N__15945\,
            I => \N__15936\
        );

    \I__3375\ : InMux
    port map (
            O => \N__15942\,
            I => \N__15933\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__15939\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__15936\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__15933\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__3371\ : InMux
    port map (
            O => \N__15926\,
            I => \N__15923\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__15923\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_4\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__15920\,
            I => \N__15917\
        );

    \I__3368\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15914\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__15914\,
            I => \N__15911\
        );

    \I__3366\ : Span12Mux_s11_v
    port map (
            O => \N__15911\,
            I => \N__15908\
        );

    \I__3365\ : Span12Mux_h
    port map (
            O => \N__15908\,
            I => \N__15904\
        );

    \I__3364\ : InMux
    port map (
            O => \N__15907\,
            I => \N__15901\
        );

    \I__3363\ : Odrv12
    port map (
            O => \N__15904\,
            I => port_rw_in
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__15901\,
            I => port_rw_in
        );

    \I__3361\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15893\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__15893\,
            I => \this_start_data_delay.M_this_state_q_srsts_0_a2_1_4\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__15890\,
            I => \this_start_data_delay.N_352_0_cascade_\
        );

    \I__3358\ : InMux
    port map (
            O => \N__15887\,
            I => \N__15884\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__15884\,
            I => \N__15881\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__15881\,
            I => \this_start_data_delay.M_this_state_q_srsts_0_0_4\
        );

    \I__3355\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15866\
        );

    \I__3354\ : InMux
    port map (
            O => \N__15877\,
            I => \N__15866\
        );

    \I__3353\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15866\
        );

    \I__3352\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15866\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15863\
        );

    \I__3350\ : Span12Mux_v
    port map (
            O => \N__15863\,
            I => \N__15860\
        );

    \I__3349\ : Span12Mux_h
    port map (
            O => \N__15860\,
            I => \N__15857\
        );

    \I__3348\ : Odrv12
    port map (
            O => \N__15857\,
            I => port_enb_c
        );

    \I__3347\ : InMux
    port map (
            O => \N__15854\,
            I => \N__15842\
        );

    \I__3346\ : InMux
    port map (
            O => \N__15853\,
            I => \N__15842\
        );

    \I__3345\ : InMux
    port map (
            O => \N__15852\,
            I => \N__15842\
        );

    \I__3344\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15842\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__15842\,
            I => \M_this_delay_clk_out_0\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__15839\,
            I => \N__15836\
        );

    \I__3341\ : InMux
    port map (
            O => \N__15836\,
            I => \N__15827\
        );

    \I__3340\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15827\
        );

    \I__3339\ : InMux
    port map (
            O => \N__15834\,
            I => \N__15827\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__15827\,
            I => \this_start_data_delay.M_last_qZ0\
        );

    \I__3337\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15821\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__15821\,
            I => \this_start_data_delay.N_352_0\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__15818\,
            I => \this_start_data_delay.N_407_cascade_\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__15815\,
            I => \N__15812\
        );

    \I__3333\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15809\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__15809\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_1\
        );

    \I__3331\ : InMux
    port map (
            O => \N__15806\,
            I => \N__15803\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__15803\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__3329\ : InMux
    port map (
            O => \N__15800\,
            I => \N__15788\
        );

    \I__3328\ : InMux
    port map (
            O => \N__15799\,
            I => \N__15788\
        );

    \I__3327\ : InMux
    port map (
            O => \N__15798\,
            I => \N__15788\
        );

    \I__3326\ : InMux
    port map (
            O => \N__15797\,
            I => \N__15788\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__15788\,
            I => \N__15785\
        );

    \I__3324\ : Span12Mux_v
    port map (
            O => \N__15785\,
            I => \N__15782\
        );

    \I__3323\ : Span12Mux_v
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__3322\ : Odrv12
    port map (
            O => \N__15779\,
            I => rst_n_c
        );

    \I__3321\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__15773\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__3319\ : IoInMux
    port map (
            O => \N__15770\,
            I => \N__15767\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__15767\,
            I => \N__15763\
        );

    \I__3317\ : InMux
    port map (
            O => \N__15766\,
            I => \N__15760\
        );

    \I__3316\ : Span4Mux_s3_v
    port map (
            O => \N__15763\,
            I => \N__15757\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__15760\,
            I => \N__15752\
        );

    \I__3314\ : Span4Mux_v
    port map (
            O => \N__15757\,
            I => \N__15752\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__15752\,
            I => \M_this_state_q_nss_0\
        );

    \I__3312\ : InMux
    port map (
            O => \N__15749\,
            I => \N__15746\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__3310\ : Odrv12
    port map (
            O => \N__15743\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__15740\,
            I => \N__15736\
        );

    \I__3308\ : InMux
    port map (
            O => \N__15739\,
            I => \N__15733\
        );

    \I__3307\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15730\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__15733\,
            I => \this_start_data_delay.N_353_0\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__15730\,
            I => \this_start_data_delay.N_353_0\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__15725\,
            I => \M_this_start_data_delay_out_0_cascade_\
        );

    \I__3303\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15719\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__15719\,
            I => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_11\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__15716\,
            I => \N__15713\
        );

    \I__3300\ : InMux
    port map (
            O => \N__15713\,
            I => \N__15709\
        );

    \I__3299\ : InMux
    port map (
            O => \N__15712\,
            I => \N__15706\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__15709\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__15706\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__15701\,
            I => \N__15698\
        );

    \I__3295\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15694\
        );

    \I__3294\ : InMux
    port map (
            O => \N__15697\,
            I => \N__15691\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__15694\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__15691\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__15686\,
            I => \N__15682\
        );

    \I__3290\ : InMux
    port map (
            O => \N__15685\,
            I => \N__15679\
        );

    \I__3289\ : InMux
    port map (
            O => \N__15682\,
            I => \N__15676\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__15679\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__15676\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__3286\ : InMux
    port map (
            O => \N__15671\,
            I => \N__15667\
        );

    \I__3285\ : InMux
    port map (
            O => \N__15670\,
            I => \N__15664\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__15667\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__15664\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__15659\,
            I => \N__15655\
        );

    \I__3281\ : InMux
    port map (
            O => \N__15658\,
            I => \N__15652\
        );

    \I__3280\ : InMux
    port map (
            O => \N__15655\,
            I => \N__15649\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__15652\,
            I => \N__15646\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__15649\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__3277\ : Odrv4
    port map (
            O => \N__15646\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__3276\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15637\
        );

    \I__3275\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15634\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__15637\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__15634\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3272\ : InMux
    port map (
            O => \N__15629\,
            I => \N__15626\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__15626\,
            I => \this_start_data_delay.M_this_state_q_srsts_i_a2_1_9Z0Z_1\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__15623\,
            I => \this_start_data_delay.M_this_state_q_srsts_i_a2_1_6Z0Z_1_cascade_\
        );

    \I__3269\ : InMux
    port map (
            O => \N__15620\,
            I => \N__15617\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__15617\,
            I => \N__15612\
        );

    \I__3267\ : InMux
    port map (
            O => \N__15616\,
            I => \N__15607\
        );

    \I__3266\ : InMux
    port map (
            O => \N__15615\,
            I => \N__15607\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__15612\,
            I => \this_start_data_delay.N_413\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__15607\,
            I => \this_start_data_delay.N_413\
        );

    \I__3263\ : InMux
    port map (
            O => \N__15602\,
            I => \N__15598\
        );

    \I__3262\ : InMux
    port map (
            O => \N__15601\,
            I => \N__15595\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__15598\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__15595\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__15590\,
            I => \N__15587\
        );

    \I__3258\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15583\
        );

    \I__3257\ : InMux
    port map (
            O => \N__15586\,
            I => \N__15580\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__15583\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__15580\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__15575\,
            I => \N__15571\
        );

    \I__3253\ : CascadeMux
    port map (
            O => \N__15574\,
            I => \N__15568\
        );

    \I__3252\ : InMux
    port map (
            O => \N__15571\,
            I => \N__15565\
        );

    \I__3251\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15562\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__15565\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__15562\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__3248\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15553\
        );

    \I__3247\ : InMux
    port map (
            O => \N__15556\,
            I => \N__15550\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__15553\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__15550\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__3244\ : InMux
    port map (
            O => \N__15545\,
            I => \N__15542\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__15542\,
            I => \this_start_data_delay.M_this_state_q_srsts_i_a2_1_8Z0Z_1\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15535\
        );

    \I__3241\ : InMux
    port map (
            O => \N__15538\,
            I => \N__15532\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__15535\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__15532\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__3238\ : InMux
    port map (
            O => \N__15527\,
            I => \N__15523\
        );

    \I__3237\ : InMux
    port map (
            O => \N__15526\,
            I => \N__15520\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__15523\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__15520\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__3234\ : CascadeMux
    port map (
            O => \N__15515\,
            I => \N__15511\
        );

    \I__3233\ : InMux
    port map (
            O => \N__15514\,
            I => \N__15508\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15505\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__15508\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__15505\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15496\
        );

    \I__3228\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15493\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__15496\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__15493\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__3225\ : InMux
    port map (
            O => \N__15488\,
            I => \N__15485\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15485\,
            I => \this_start_data_delay.M_this_state_q_srsts_i_a2_1_7Z0Z_1\
        );

    \I__3223\ : SRMux
    port map (
            O => \N__15482\,
            I => \N__15479\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__15479\,
            I => \N__15475\
        );

    \I__3221\ : SRMux
    port map (
            O => \N__15478\,
            I => \N__15472\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__15475\,
            I => \N__15467\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__15472\,
            I => \N__15467\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__15467\,
            I => \M_this_state_q_RNI20CEZ0Z_0\
        );

    \I__3217\ : InMux
    port map (
            O => \N__15464\,
            I => \N__15461\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__15461\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__3215\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15453\
        );

    \I__3214\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15448\
        );

    \I__3213\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15448\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__15453\,
            I => \N__15442\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__15448\,
            I => \N__15439\
        );

    \I__3210\ : InMux
    port map (
            O => \N__15447\,
            I => \N__15436\
        );

    \I__3209\ : InMux
    port map (
            O => \N__15446\,
            I => \N__15432\
        );

    \I__3208\ : InMux
    port map (
            O => \N__15445\,
            I => \N__15429\
        );

    \I__3207\ : Span4Mux_v
    port map (
            O => \N__15442\,
            I => \N__15422\
        );

    \I__3206\ : Span4Mux_v
    port map (
            O => \N__15439\,
            I => \N__15422\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__15436\,
            I => \N__15422\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15435\,
            I => \N__15419\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__15432\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__15429\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__15422\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__15419\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3199\ : InMux
    port map (
            O => \N__15410\,
            I => \N__15406\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__15409\,
            I => \N__15403\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__15406\,
            I => \N__15400\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15397\
        );

    \I__3195\ : Odrv4
    port map (
            O => \N__15400\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_1\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__15397\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_1\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__15392\,
            I => \N__15388\
        );

    \I__3192\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15385\
        );

    \I__3191\ : InMux
    port map (
            O => \N__15388\,
            I => \N__15378\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__15385\,
            I => \N__15375\
        );

    \I__3189\ : InMux
    port map (
            O => \N__15384\,
            I => \N__15368\
        );

    \I__3188\ : InMux
    port map (
            O => \N__15383\,
            I => \N__15368\
        );

    \I__3187\ : InMux
    port map (
            O => \N__15382\,
            I => \N__15368\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__15381\,
            I => \N__15365\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__15378\,
            I => \N__15362\
        );

    \I__3184\ : Span4Mux_h
    port map (
            O => \N__15375\,
            I => \N__15359\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__15368\,
            I => \N__15356\
        );

    \I__3182\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15353\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__15362\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__3180\ : Odrv4
    port map (
            O => \N__15359\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__15356\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__15353\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__3177\ : InMux
    port map (
            O => \N__15344\,
            I => \N__15341\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__15341\,
            I => \N__15337\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15340\,
            I => \N__15334\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__15337\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_3\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__15334\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_3\
        );

    \I__3172\ : CEMux
    port map (
            O => \N__15329\,
            I => \N__15324\
        );

    \I__3171\ : CEMux
    port map (
            O => \N__15328\,
            I => \N__15321\
        );

    \I__3170\ : CEMux
    port map (
            O => \N__15327\,
            I => \N__15318\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__15324\,
            I => \N__15313\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__15321\,
            I => \N__15308\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__15318\,
            I => \N__15308\
        );

    \I__3166\ : CEMux
    port map (
            O => \N__15317\,
            I => \N__15303\
        );

    \I__3165\ : CEMux
    port map (
            O => \N__15316\,
            I => \N__15300\
        );

    \I__3164\ : Span4Mux_v
    port map (
            O => \N__15313\,
            I => \N__15296\
        );

    \I__3163\ : Span4Mux_v
    port map (
            O => \N__15308\,
            I => \N__15293\
        );

    \I__3162\ : CEMux
    port map (
            O => \N__15307\,
            I => \N__15289\
        );

    \I__3161\ : CEMux
    port map (
            O => \N__15306\,
            I => \N__15286\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__15303\,
            I => \N__15283\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__15300\,
            I => \N__15280\
        );

    \I__3158\ : CEMux
    port map (
            O => \N__15299\,
            I => \N__15277\
        );

    \I__3157\ : Span4Mux_v
    port map (
            O => \N__15296\,
            I => \N__15272\
        );

    \I__3156\ : Span4Mux_h
    port map (
            O => \N__15293\,
            I => \N__15272\
        );

    \I__3155\ : CEMux
    port map (
            O => \N__15292\,
            I => \N__15269\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__15289\,
            I => \N__15265\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__15286\,
            I => \N__15262\
        );

    \I__3152\ : Span4Mux_v
    port map (
            O => \N__15283\,
            I => \N__15259\
        );

    \I__3151\ : Span4Mux_v
    port map (
            O => \N__15280\,
            I => \N__15256\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__15277\,
            I => \N__15253\
        );

    \I__3149\ : Span4Mux_h
    port map (
            O => \N__15272\,
            I => \N__15248\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__15269\,
            I => \N__15248\
        );

    \I__3147\ : CEMux
    port map (
            O => \N__15268\,
            I => \N__15245\
        );

    \I__3146\ : Span4Mux_h
    port map (
            O => \N__15265\,
            I => \N__15242\
        );

    \I__3145\ : Span4Mux_h
    port map (
            O => \N__15262\,
            I => \N__15239\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__15259\,
            I => \N__15232\
        );

    \I__3143\ : Span4Mux_h
    port map (
            O => \N__15256\,
            I => \N__15232\
        );

    \I__3142\ : Span4Mux_v
    port map (
            O => \N__15253\,
            I => \N__15232\
        );

    \I__3141\ : Span4Mux_v
    port map (
            O => \N__15248\,
            I => \N__15227\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__15245\,
            I => \N__15227\
        );

    \I__3139\ : Odrv4
    port map (
            O => \N__15242\,
            I => \this_vga_signals.N_550_2\
        );

    \I__3138\ : Odrv4
    port map (
            O => \N__15239\,
            I => \this_vga_signals.N_550_2\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__15232\,
            I => \this_vga_signals.N_550_2\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__15227\,
            I => \this_vga_signals.N_550_2\
        );

    \I__3135\ : SRMux
    port map (
            O => \N__15218\,
            I => \N__15212\
        );

    \I__3134\ : SRMux
    port map (
            O => \N__15217\,
            I => \N__15208\
        );

    \I__3133\ : SRMux
    port map (
            O => \N__15216\,
            I => \N__15205\
        );

    \I__3132\ : SRMux
    port map (
            O => \N__15215\,
            I => \N__15201\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__15212\,
            I => \N__15198\
        );

    \I__3130\ : SRMux
    port map (
            O => \N__15211\,
            I => \N__15194\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__15208\,
            I => \N__15190\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__15205\,
            I => \N__15187\
        );

    \I__3127\ : SRMux
    port map (
            O => \N__15204\,
            I => \N__15184\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__15201\,
            I => \N__15180\
        );

    \I__3125\ : Span4Mux_v
    port map (
            O => \N__15198\,
            I => \N__15176\
        );

    \I__3124\ : SRMux
    port map (
            O => \N__15197\,
            I => \N__15173\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__15194\,
            I => \N__15170\
        );

    \I__3122\ : SRMux
    port map (
            O => \N__15193\,
            I => \N__15167\
        );

    \I__3121\ : Span4Mux_v
    port map (
            O => \N__15190\,
            I => \N__15162\
        );

    \I__3120\ : Span4Mux_v
    port map (
            O => \N__15187\,
            I => \N__15162\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__15184\,
            I => \N__15159\
        );

    \I__3118\ : SRMux
    port map (
            O => \N__15183\,
            I => \N__15156\
        );

    \I__3117\ : Span4Mux_h
    port map (
            O => \N__15180\,
            I => \N__15153\
        );

    \I__3116\ : SRMux
    port map (
            O => \N__15179\,
            I => \N__15150\
        );

    \I__3115\ : Span4Mux_h
    port map (
            O => \N__15176\,
            I => \N__15147\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__15173\,
            I => \N__15144\
        );

    \I__3113\ : Span4Mux_h
    port map (
            O => \N__15170\,
            I => \N__15139\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__15167\,
            I => \N__15139\
        );

    \I__3111\ : Span4Mux_v
    port map (
            O => \N__15162\,
            I => \N__15132\
        );

    \I__3110\ : Span4Mux_v
    port map (
            O => \N__15159\,
            I => \N__15132\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15156\,
            I => \N__15132\
        );

    \I__3108\ : Span4Mux_h
    port map (
            O => \N__15153\,
            I => \N__15127\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__15150\,
            I => \N__15127\
        );

    \I__3106\ : Span4Mux_h
    port map (
            O => \N__15147\,
            I => \N__15123\
        );

    \I__3105\ : Span4Mux_v
    port map (
            O => \N__15144\,
            I => \N__15120\
        );

    \I__3104\ : Span4Mux_h
    port map (
            O => \N__15139\,
            I => \N__15115\
        );

    \I__3103\ : Span4Mux_h
    port map (
            O => \N__15132\,
            I => \N__15115\
        );

    \I__3102\ : Sp12to4
    port map (
            O => \N__15127\,
            I => \N__15112\
        );

    \I__3101\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15109\
        );

    \I__3100\ : Odrv4
    port map (
            O => \N__15123\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9\
        );

    \I__3099\ : Odrv4
    port map (
            O => \N__15120\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__15115\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9\
        );

    \I__3097\ : Odrv12
    port map (
            O => \N__15112\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__15109\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9\
        );

    \I__3095\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15094\
        );

    \I__3094\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15091\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__15094\,
            I => \N__15088\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__15091\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__15088\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__3090\ : CascadeMux
    port map (
            O => \N__15083\,
            I => \N__15079\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15074\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15074\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__15074\,
            I => \N__15064\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15061\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15072\,
            I => \N__15052\
        );

    \I__3084\ : InMux
    port map (
            O => \N__15071\,
            I => \N__15052\
        );

    \I__3083\ : InMux
    port map (
            O => \N__15070\,
            I => \N__15052\
        );

    \I__3082\ : InMux
    port map (
            O => \N__15069\,
            I => \N__15052\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__15068\,
            I => \N__15047\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15044\
        );

    \I__3079\ : Span4Mux_v
    port map (
            O => \N__15064\,
            I => \N__15037\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__15061\,
            I => \N__15037\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__15052\,
            I => \N__15037\
        );

    \I__3076\ : CascadeMux
    port map (
            O => \N__15051\,
            I => \N__15034\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15029\
        );

    \I__3074\ : InMux
    port map (
            O => \N__15047\,
            I => \N__15029\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__15044\,
            I => \N__15024\
        );

    \I__3072\ : Span4Mux_v
    port map (
            O => \N__15037\,
            I => \N__15024\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15034\,
            I => \N__15021\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__15029\,
            I => \N__15018\
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__15024\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__15021\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3067\ : Odrv12
    port map (
            O => \N__15018\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__3066\ : CEMux
    port map (
            O => \N__15011\,
            I => \N__15008\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__15008\,
            I => \N__15004\
        );

    \I__3064\ : CEMux
    port map (
            O => \N__15007\,
            I => \N__15000\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__15004\,
            I => \N__14997\
        );

    \I__3062\ : CEMux
    port map (
            O => \N__15003\,
            I => \N__14994\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__15000\,
            I => \N__14991\
        );

    \I__3060\ : Span4Mux_h
    port map (
            O => \N__14997\,
            I => \N__14985\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__14994\,
            I => \N__14985\
        );

    \I__3058\ : Span4Mux_h
    port map (
            O => \N__14991\,
            I => \N__14982\
        );

    \I__3057\ : CEMux
    port map (
            O => \N__14990\,
            I => \N__14979\
        );

    \I__3056\ : Span4Mux_h
    port map (
            O => \N__14985\,
            I => \N__14976\
        );

    \I__3055\ : Sp12to4
    port map (
            O => \N__14982\,
            I => \N__14971\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__14979\,
            I => \N__14971\
        );

    \I__3053\ : Odrv4
    port map (
            O => \N__14976\,
            I => \this_vga_signals.N_550_0\
        );

    \I__3052\ : Odrv12
    port map (
            O => \N__14971\,
            I => \this_vga_signals.N_550_0\
        );

    \I__3051\ : SRMux
    port map (
            O => \N__14966\,
            I => \N__14962\
        );

    \I__3050\ : SRMux
    port map (
            O => \N__14965\,
            I => \N__14959\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__14962\,
            I => \N__14954\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__14959\,
            I => \N__14951\
        );

    \I__3047\ : SRMux
    port map (
            O => \N__14958\,
            I => \N__14948\
        );

    \I__3046\ : SRMux
    port map (
            O => \N__14957\,
            I => \N__14945\
        );

    \I__3045\ : Span4Mux_v
    port map (
            O => \N__14954\,
            I => \N__14942\
        );

    \I__3044\ : Span4Mux_v
    port map (
            O => \N__14951\,
            I => \N__14937\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__14948\,
            I => \N__14937\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__14945\,
            I => \N__14933\
        );

    \I__3041\ : Span4Mux_h
    port map (
            O => \N__14942\,
            I => \N__14928\
        );

    \I__3040\ : Span4Mux_h
    port map (
            O => \N__14937\,
            I => \N__14925\
        );

    \I__3039\ : SRMux
    port map (
            O => \N__14936\,
            I => \N__14922\
        );

    \I__3038\ : Span4Mux_h
    port map (
            O => \N__14933\,
            I => \N__14919\
        );

    \I__3037\ : SRMux
    port map (
            O => \N__14932\,
            I => \N__14916\
        );

    \I__3036\ : InMux
    port map (
            O => \N__14931\,
            I => \N__14913\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__14928\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__14925\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__14922\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9\
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__14919\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__14916\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__14913\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9\
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__14900\,
            I => \this_start_data_delay.M_this_state_q_srsts_i_1_2_cascade_\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__14897\,
            I => \N__14894\
        );

    \I__3027\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14891\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__14891\,
            I => \this_start_data_delay.N_389_1\
        );

    \I__3025\ : IoInMux
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__14885\,
            I => \N__14882\
        );

    \I__3023\ : Span4Mux_s0_h
    port map (
            O => \N__14882\,
            I => \N__14879\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__14879\,
            I => \N__14875\
        );

    \I__3021\ : InMux
    port map (
            O => \N__14878\,
            I => \N__14871\
        );

    \I__3020\ : Sp12to4
    port map (
            O => \N__14875\,
            I => \N__14868\
        );

    \I__3019\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14865\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__14871\,
            I => \N__14862\
        );

    \I__3017\ : Span12Mux_v
    port map (
            O => \N__14868\,
            I => \N__14858\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__14865\,
            I => \N__14855\
        );

    \I__3015\ : Span12Mux_v
    port map (
            O => \N__14862\,
            I => \N__14852\
        );

    \I__3014\ : InMux
    port map (
            O => \N__14861\,
            I => \N__14849\
        );

    \I__3013\ : Span12Mux_h
    port map (
            O => \N__14858\,
            I => \N__14846\
        );

    \I__3012\ : Span12Mux_s7_h
    port map (
            O => \N__14855\,
            I => \N__14843\
        );

    \I__3011\ : Span12Mux_h
    port map (
            O => \N__14852\,
            I => \N__14840\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__14849\,
            I => \N__14837\
        );

    \I__3009\ : Odrv12
    port map (
            O => \N__14846\,
            I => port_dmab_c
        );

    \I__3008\ : Odrv12
    port map (
            O => \N__14843\,
            I => port_dmab_c
        );

    \I__3007\ : Odrv12
    port map (
            O => \N__14840\,
            I => port_dmab_c
        );

    \I__3006\ : Odrv4
    port map (
            O => \N__14837\,
            I => port_dmab_c
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__14828\,
            I => \port_dmab_c_cascade_\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__14825\,
            I => \this_start_data_delay.N_385_cascade_\
        );

    \I__3003\ : InMux
    port map (
            O => \N__14822\,
            I => \bfn_16_25_0_\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__14819\,
            I => \this_vga_signals.mult1_un54_sum_1_c2_1_cascade_\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__14816\,
            I => \N__14809\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__14815\,
            I => \N__14806\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__14814\,
            I => \N__14803\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__14813\,
            I => \N__14795\
        );

    \I__2997\ : InMux
    port map (
            O => \N__14812\,
            I => \N__14792\
        );

    \I__2996\ : InMux
    port map (
            O => \N__14809\,
            I => \N__14786\
        );

    \I__2995\ : InMux
    port map (
            O => \N__14806\,
            I => \N__14783\
        );

    \I__2994\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14780\
        );

    \I__2993\ : InMux
    port map (
            O => \N__14802\,
            I => \N__14777\
        );

    \I__2992\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14774\
        );

    \I__2991\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14771\
        );

    \I__2990\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14767\
        );

    \I__2989\ : InMux
    port map (
            O => \N__14798\,
            I => \N__14762\
        );

    \I__2988\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14762\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__14792\,
            I => \N__14759\
        );

    \I__2986\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14755\
        );

    \I__2985\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14747\
        );

    \I__2984\ : InMux
    port map (
            O => \N__14789\,
            I => \N__14742\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__14786\,
            I => \N__14735\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__14783\,
            I => \N__14735\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__14780\,
            I => \N__14726\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__14777\,
            I => \N__14726\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__14774\,
            I => \N__14726\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__14771\,
            I => \N__14726\
        );

    \I__2977\ : InMux
    port map (
            O => \N__14770\,
            I => \N__14723\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__14767\,
            I => \N__14718\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__14762\,
            I => \N__14718\
        );

    \I__2974\ : Span4Mux_v
    port map (
            O => \N__14759\,
            I => \N__14714\
        );

    \I__2973\ : InMux
    port map (
            O => \N__14758\,
            I => \N__14711\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__14755\,
            I => \N__14708\
        );

    \I__2971\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14705\
        );

    \I__2970\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14700\
        );

    \I__2969\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14700\
        );

    \I__2968\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14695\
        );

    \I__2967\ : InMux
    port map (
            O => \N__14750\,
            I => \N__14695\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__14747\,
            I => \N__14692\
        );

    \I__2965\ : InMux
    port map (
            O => \N__14746\,
            I => \N__14689\
        );

    \I__2964\ : InMux
    port map (
            O => \N__14745\,
            I => \N__14686\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__14742\,
            I => \N__14683\
        );

    \I__2962\ : InMux
    port map (
            O => \N__14741\,
            I => \N__14680\
        );

    \I__2961\ : InMux
    port map (
            O => \N__14740\,
            I => \N__14677\
        );

    \I__2960\ : Span4Mux_v
    port map (
            O => \N__14735\,
            I => \N__14672\
        );

    \I__2959\ : Span4Mux_v
    port map (
            O => \N__14726\,
            I => \N__14672\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__14723\,
            I => \N__14667\
        );

    \I__2957\ : Span4Mux_h
    port map (
            O => \N__14718\,
            I => \N__14667\
        );

    \I__2956\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14664\
        );

    \I__2955\ : Span4Mux_h
    port map (
            O => \N__14714\,
            I => \N__14653\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__14711\,
            I => \N__14653\
        );

    \I__2953\ : Span4Mux_v
    port map (
            O => \N__14708\,
            I => \N__14653\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__14705\,
            I => \N__14653\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__14700\,
            I => \N__14653\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__14695\,
            I => \N__14644\
        );

    \I__2949\ : Span4Mux_h
    port map (
            O => \N__14692\,
            I => \N__14644\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__14689\,
            I => \N__14644\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__14686\,
            I => \N__14644\
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__14683\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__14680\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__14677\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__14672\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__14667\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__14664\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2940\ : Odrv4
    port map (
            O => \N__14653\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2939\ : Odrv4
    port map (
            O => \N__14644\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2938\ : InMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__14624\,
            I => \N__14621\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__14621\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2Z0Z_9\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__14618\,
            I => \this_vga_signals.mult1_un54_sum_1_c2_cascade_\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__14615\,
            I => \N__14612\
        );

    \I__2933\ : InMux
    port map (
            O => \N__14612\,
            I => \N__14603\
        );

    \I__2932\ : InMux
    port map (
            O => \N__14611\,
            I => \N__14595\
        );

    \I__2931\ : InMux
    port map (
            O => \N__14610\,
            I => \N__14595\
        );

    \I__2930\ : InMux
    port map (
            O => \N__14609\,
            I => \N__14595\
        );

    \I__2929\ : InMux
    port map (
            O => \N__14608\,
            I => \N__14592\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__14607\,
            I => \N__14588\
        );

    \I__2927\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14585\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__14603\,
            I => \N__14582\
        );

    \I__2925\ : InMux
    port map (
            O => \N__14602\,
            I => \N__14579\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__14595\,
            I => \N__14572\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__14592\,
            I => \N__14572\
        );

    \I__2922\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14569\
        );

    \I__2921\ : InMux
    port map (
            O => \N__14588\,
            I => \N__14566\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__14585\,
            I => \N__14561\
        );

    \I__2919\ : Span4Mux_v
    port map (
            O => \N__14582\,
            I => \N__14556\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__14579\,
            I => \N__14556\
        );

    \I__2917\ : InMux
    port map (
            O => \N__14578\,
            I => \N__14553\
        );

    \I__2916\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14550\
        );

    \I__2915\ : Span4Mux_h
    port map (
            O => \N__14572\,
            I => \N__14547\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__14569\,
            I => \N__14542\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__14566\,
            I => \N__14542\
        );

    \I__2912\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14539\
        );

    \I__2911\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14536\
        );

    \I__2910\ : Span4Mux_h
    port map (
            O => \N__14561\,
            I => \N__14525\
        );

    \I__2909\ : Span4Mux_h
    port map (
            O => \N__14556\,
            I => \N__14525\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__14553\,
            I => \N__14520\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14550\,
            I => \N__14520\
        );

    \I__2906\ : Span4Mux_h
    port map (
            O => \N__14547\,
            I => \N__14511\
        );

    \I__2905\ : Span4Mux_h
    port map (
            O => \N__14542\,
            I => \N__14511\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__14539\,
            I => \N__14511\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__14536\,
            I => \N__14511\
        );

    \I__2902\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14506\
        );

    \I__2901\ : InMux
    port map (
            O => \N__14534\,
            I => \N__14506\
        );

    \I__2900\ : InMux
    port map (
            O => \N__14533\,
            I => \N__14501\
        );

    \I__2899\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14501\
        );

    \I__2898\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14496\
        );

    \I__2897\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14496\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__14525\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2895\ : Odrv12
    port map (
            O => \N__14520\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__14511\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__14506\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__14501\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__14496\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__14483\,
            I => \N__14473\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__14482\,
            I => \N__14467\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__14481\,
            I => \N__14464\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__14480\,
            I => \N__14459\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__14479\,
            I => \N__14456\
        );

    \I__2885\ : InMux
    port map (
            O => \N__14478\,
            I => \N__14453\
        );

    \I__2884\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14450\
        );

    \I__2883\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14444\
        );

    \I__2882\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14444\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__14472\,
            I => \N__14441\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__14471\,
            I => \N__14438\
        );

    \I__2879\ : InMux
    port map (
            O => \N__14470\,
            I => \N__14434\
        );

    \I__2878\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14431\
        );

    \I__2877\ : InMux
    port map (
            O => \N__14464\,
            I => \N__14428\
        );

    \I__2876\ : InMux
    port map (
            O => \N__14463\,
            I => \N__14423\
        );

    \I__2875\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14423\
        );

    \I__2874\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14418\
        );

    \I__2873\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14418\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__14453\,
            I => \N__14415\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__14450\,
            I => \N__14412\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__14449\,
            I => \N__14409\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__14444\,
            I => \N__14405\
        );

    \I__2868\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14402\
        );

    \I__2867\ : InMux
    port map (
            O => \N__14438\,
            I => \N__14399\
        );

    \I__2866\ : InMux
    port map (
            O => \N__14437\,
            I => \N__14394\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__14434\,
            I => \N__14391\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__14431\,
            I => \N__14388\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__14428\,
            I => \N__14385\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__14423\,
            I => \N__14380\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__14418\,
            I => \N__14380\
        );

    \I__2860\ : Span4Mux_v
    port map (
            O => \N__14415\,
            I => \N__14377\
        );

    \I__2859\ : Span4Mux_v
    port map (
            O => \N__14412\,
            I => \N__14374\
        );

    \I__2858\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14371\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14408\,
            I => \N__14368\
        );

    \I__2856\ : Span4Mux_v
    port map (
            O => \N__14405\,
            I => \N__14365\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__14402\,
            I => \N__14362\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__14399\,
            I => \N__14359\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__14398\,
            I => \N__14356\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__14397\,
            I => \N__14353\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__14394\,
            I => \N__14348\
        );

    \I__2850\ : Span4Mux_v
    port map (
            O => \N__14391\,
            I => \N__14348\
        );

    \I__2849\ : Span4Mux_h
    port map (
            O => \N__14388\,
            I => \N__14341\
        );

    \I__2848\ : Span4Mux_h
    port map (
            O => \N__14385\,
            I => \N__14341\
        );

    \I__2847\ : Span4Mux_v
    port map (
            O => \N__14380\,
            I => \N__14341\
        );

    \I__2846\ : Span4Mux_v
    port map (
            O => \N__14377\,
            I => \N__14336\
        );

    \I__2845\ : Span4Mux_h
    port map (
            O => \N__14374\,
            I => \N__14336\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__14371\,
            I => \N__14331\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__14368\,
            I => \N__14331\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__14365\,
            I => \N__14324\
        );

    \I__2841\ : Span4Mux_v
    port map (
            O => \N__14362\,
            I => \N__14324\
        );

    \I__2840\ : Span4Mux_v
    port map (
            O => \N__14359\,
            I => \N__14324\
        );

    \I__2839\ : InMux
    port map (
            O => \N__14356\,
            I => \N__14319\
        );

    \I__2838\ : InMux
    port map (
            O => \N__14353\,
            I => \N__14319\
        );

    \I__2837\ : Span4Mux_v
    port map (
            O => \N__14348\,
            I => \N__14314\
        );

    \I__2836\ : Span4Mux_h
    port map (
            O => \N__14341\,
            I => \N__14314\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__14336\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2834\ : Odrv12
    port map (
            O => \N__14331\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__14324\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__14319\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__14314\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__14303\,
            I => \N__14299\
        );

    \I__2829\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14293\
        );

    \I__2828\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14287\
        );

    \I__2827\ : InMux
    port map (
            O => \N__14298\,
            I => \N__14287\
        );

    \I__2826\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14284\
        );

    \I__2825\ : InMux
    port map (
            O => \N__14296\,
            I => \N__14280\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__14293\,
            I => \N__14275\
        );

    \I__2823\ : InMux
    port map (
            O => \N__14292\,
            I => \N__14272\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__14287\,
            I => \N__14268\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__14284\,
            I => \N__14260\
        );

    \I__2820\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14255\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__14280\,
            I => \N__14252\
        );

    \I__2818\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14249\
        );

    \I__2817\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14246\
        );

    \I__2816\ : Span4Mux_v
    port map (
            O => \N__14275\,
            I => \N__14243\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__14272\,
            I => \N__14240\
        );

    \I__2814\ : InMux
    port map (
            O => \N__14271\,
            I => \N__14237\
        );

    \I__2813\ : Span4Mux_v
    port map (
            O => \N__14268\,
            I => \N__14234\
        );

    \I__2812\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14231\
        );

    \I__2811\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14228\
        );

    \I__2810\ : InMux
    port map (
            O => \N__14265\,
            I => \N__14225\
        );

    \I__2809\ : InMux
    port map (
            O => \N__14264\,
            I => \N__14220\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14263\,
            I => \N__14220\
        );

    \I__2807\ : Span4Mux_v
    port map (
            O => \N__14260\,
            I => \N__14216\
        );

    \I__2806\ : InMux
    port map (
            O => \N__14259\,
            I => \N__14213\
        );

    \I__2805\ : InMux
    port map (
            O => \N__14258\,
            I => \N__14210\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__14255\,
            I => \N__14205\
        );

    \I__2803\ : Span4Mux_v
    port map (
            O => \N__14252\,
            I => \N__14205\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__14249\,
            I => \N__14200\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__14246\,
            I => \N__14200\
        );

    \I__2800\ : Span4Mux_h
    port map (
            O => \N__14243\,
            I => \N__14191\
        );

    \I__2799\ : Span4Mux_h
    port map (
            O => \N__14240\,
            I => \N__14191\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__14237\,
            I => \N__14191\
        );

    \I__2797\ : Span4Mux_h
    port map (
            O => \N__14234\,
            I => \N__14182\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__14231\,
            I => \N__14182\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__14228\,
            I => \N__14182\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__14225\,
            I => \N__14182\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__14220\,
            I => \N__14179\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__14219\,
            I => \N__14174\
        );

    \I__2791\ : Sp12to4
    port map (
            O => \N__14216\,
            I => \N__14167\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__14213\,
            I => \N__14167\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__14210\,
            I => \N__14167\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__14205\,
            I => \N__14162\
        );

    \I__2787\ : Span4Mux_v
    port map (
            O => \N__14200\,
            I => \N__14162\
        );

    \I__2786\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14157\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14198\,
            I => \N__14157\
        );

    \I__2784\ : Span4Mux_v
    port map (
            O => \N__14191\,
            I => \N__14150\
        );

    \I__2783\ : Span4Mux_v
    port map (
            O => \N__14182\,
            I => \N__14150\
        );

    \I__2782\ : Span4Mux_h
    port map (
            O => \N__14179\,
            I => \N__14150\
        );

    \I__2781\ : InMux
    port map (
            O => \N__14178\,
            I => \N__14147\
        );

    \I__2780\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14144\
        );

    \I__2779\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14141\
        );

    \I__2778\ : Odrv12
    port map (
            O => \N__14167\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__14162\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__14157\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__14150\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__14147\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__14144\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__14141\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__14126\,
            I => \N__14123\
        );

    \I__2770\ : InMux
    port map (
            O => \N__14123\,
            I => \N__14120\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__14120\,
            I => \N__14108\
        );

    \I__2768\ : InMux
    port map (
            O => \N__14119\,
            I => \N__14103\
        );

    \I__2767\ : InMux
    port map (
            O => \N__14118\,
            I => \N__14103\
        );

    \I__2766\ : InMux
    port map (
            O => \N__14117\,
            I => \N__14099\
        );

    \I__2765\ : InMux
    port map (
            O => \N__14116\,
            I => \N__14094\
        );

    \I__2764\ : InMux
    port map (
            O => \N__14115\,
            I => \N__14087\
        );

    \I__2763\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14087\
        );

    \I__2762\ : InMux
    port map (
            O => \N__14113\,
            I => \N__14084\
        );

    \I__2761\ : InMux
    port map (
            O => \N__14112\,
            I => \N__14081\
        );

    \I__2760\ : InMux
    port map (
            O => \N__14111\,
            I => \N__14078\
        );

    \I__2759\ : Span4Mux_v
    port map (
            O => \N__14108\,
            I => \N__14071\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__14103\,
            I => \N__14071\
        );

    \I__2757\ : InMux
    port map (
            O => \N__14102\,
            I => \N__14068\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__14099\,
            I => \N__14065\
        );

    \I__2755\ : InMux
    port map (
            O => \N__14098\,
            I => \N__14062\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14097\,
            I => \N__14059\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__14094\,
            I => \N__14056\
        );

    \I__2752\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14053\
        );

    \I__2751\ : InMux
    port map (
            O => \N__14092\,
            I => \N__14050\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__14087\,
            I => \N__14045\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__14084\,
            I => \N__14045\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__14081\,
            I => \N__14040\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__14078\,
            I => \N__14040\
        );

    \I__2746\ : InMux
    port map (
            O => \N__14077\,
            I => \N__14035\
        );

    \I__2745\ : InMux
    port map (
            O => \N__14076\,
            I => \N__14032\
        );

    \I__2744\ : Span4Mux_h
    port map (
            O => \N__14071\,
            I => \N__14027\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__14068\,
            I => \N__14027\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__14065\,
            I => \N__14020\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__14062\,
            I => \N__14020\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__14059\,
            I => \N__14020\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__14056\,
            I => \N__14015\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__14053\,
            I => \N__14015\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__14050\,
            I => \N__14012\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__14045\,
            I => \N__14007\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__14040\,
            I => \N__14007\
        );

    \I__2734\ : InMux
    port map (
            O => \N__14039\,
            I => \N__14002\
        );

    \I__2733\ : InMux
    port map (
            O => \N__14038\,
            I => \N__14002\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__14035\,
            I => \N__13994\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__14032\,
            I => \N__13994\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__14027\,
            I => \N__13985\
        );

    \I__2729\ : Span4Mux_v
    port map (
            O => \N__14020\,
            I => \N__13985\
        );

    \I__2728\ : Span4Mux_v
    port map (
            O => \N__14015\,
            I => \N__13985\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__14012\,
            I => \N__13985\
        );

    \I__2726\ : Span4Mux_h
    port map (
            O => \N__14007\,
            I => \N__13980\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__14002\,
            I => \N__13980\
        );

    \I__2724\ : InMux
    port map (
            O => \N__14001\,
            I => \N__13975\
        );

    \I__2723\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13975\
        );

    \I__2722\ : InMux
    port map (
            O => \N__13999\,
            I => \N__13972\
        );

    \I__2721\ : Odrv12
    port map (
            O => \N__13994\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__13985\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__13980\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__13975\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__13972\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2716\ : InMux
    port map (
            O => \N__13961\,
            I => \N__13958\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__13958\,
            I => \this_vga_signals.mult1_un54_sum1_i_1_3\
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__13955\,
            I => \N__13952\
        );

    \I__2713\ : CascadeBuf
    port map (
            O => \N__13952\,
            I => \N__13949\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__13949\,
            I => \N__13946\
        );

    \I__2711\ : CascadeBuf
    port map (
            O => \N__13946\,
            I => \N__13943\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__13943\,
            I => \N__13940\
        );

    \I__2709\ : CascadeBuf
    port map (
            O => \N__13940\,
            I => \N__13937\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__13937\,
            I => \N__13934\
        );

    \I__2707\ : CascadeBuf
    port map (
            O => \N__13934\,
            I => \N__13931\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__13931\,
            I => \N__13928\
        );

    \I__2705\ : CascadeBuf
    port map (
            O => \N__13928\,
            I => \N__13925\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__13925\,
            I => \N__13922\
        );

    \I__2703\ : CascadeBuf
    port map (
            O => \N__13922\,
            I => \N__13919\
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__13919\,
            I => \N__13916\
        );

    \I__2701\ : CascadeBuf
    port map (
            O => \N__13916\,
            I => \N__13913\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__13913\,
            I => \N__13910\
        );

    \I__2699\ : CascadeBuf
    port map (
            O => \N__13910\,
            I => \N__13907\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__13907\,
            I => \N__13904\
        );

    \I__2697\ : CascadeBuf
    port map (
            O => \N__13904\,
            I => \N__13901\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__13901\,
            I => \N__13898\
        );

    \I__2695\ : CascadeBuf
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__2693\ : CascadeBuf
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__13889\,
            I => \N__13886\
        );

    \I__2691\ : CascadeBuf
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__13883\,
            I => \N__13880\
        );

    \I__2689\ : CascadeBuf
    port map (
            O => \N__13880\,
            I => \N__13877\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__2687\ : CascadeBuf
    port map (
            O => \N__13874\,
            I => \N__13871\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__13871\,
            I => \N__13868\
        );

    \I__2685\ : CascadeBuf
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__13865\,
            I => \N__13862\
        );

    \I__2683\ : InMux
    port map (
            O => \N__13862\,
            I => \N__13859\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__2681\ : Span12Mux_h
    port map (
            O => \N__13856\,
            I => \N__13853\
        );

    \I__2680\ : Span12Mux_v
    port map (
            O => \N__13853\,
            I => \N__13850\
        );

    \I__2679\ : Odrv12
    port map (
            O => \N__13850\,
            I => \M_this_vga_signals_address_5\
        );

    \I__2678\ : InMux
    port map (
            O => \N__13847\,
            I => \un1_M_this_data_count_q_cry_2\
        );

    \I__2677\ : InMux
    port map (
            O => \N__13844\,
            I => \un1_M_this_data_count_q_cry_3\
        );

    \I__2676\ : InMux
    port map (
            O => \N__13841\,
            I => \un1_M_this_data_count_q_cry_4\
        );

    \I__2675\ : InMux
    port map (
            O => \N__13838\,
            I => \un1_M_this_data_count_q_cry_5\
        );

    \I__2674\ : InMux
    port map (
            O => \N__13835\,
            I => \un1_M_this_data_count_q_cry_6\
        );

    \I__2673\ : InMux
    port map (
            O => \N__13832\,
            I => \bfn_16_24_0_\
        );

    \I__2672\ : InMux
    port map (
            O => \N__13829\,
            I => \un1_M_this_data_count_q_cry_8\
        );

    \I__2671\ : InMux
    port map (
            O => \N__13826\,
            I => \un1_M_this_data_count_q_cry_9\
        );

    \I__2670\ : InMux
    port map (
            O => \N__13823\,
            I => \un1_M_this_data_count_q_cry_10\
        );

    \I__2669\ : InMux
    port map (
            O => \N__13820\,
            I => \un1_M_this_data_count_q_cry_11\
        );

    \I__2668\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13814\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__13814\,
            I => \N__13811\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__13811\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__13808\,
            I => \N__13800\
        );

    \I__2664\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13791\
        );

    \I__2663\ : InMux
    port map (
            O => \N__13806\,
            I => \N__13785\
        );

    \I__2662\ : InMux
    port map (
            O => \N__13805\,
            I => \N__13785\
        );

    \I__2661\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13776\
        );

    \I__2660\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13776\
        );

    \I__2659\ : InMux
    port map (
            O => \N__13800\,
            I => \N__13776\
        );

    \I__2658\ : InMux
    port map (
            O => \N__13799\,
            I => \N__13776\
        );

    \I__2657\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13773\
        );

    \I__2656\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13768\
        );

    \I__2655\ : InMux
    port map (
            O => \N__13796\,
            I => \N__13768\
        );

    \I__2654\ : InMux
    port map (
            O => \N__13795\,
            I => \N__13763\
        );

    \I__2653\ : InMux
    port map (
            O => \N__13794\,
            I => \N__13763\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__13791\,
            I => \N__13760\
        );

    \I__2651\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13757\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__13785\,
            I => \N__13752\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__13776\,
            I => \N__13752\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__13773\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__13768\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__13763\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__13760\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__13757\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__13752\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2642\ : InMux
    port map (
            O => \N__13739\,
            I => \N__13735\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__13738\,
            I => \N__13732\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__13735\,
            I => \N__13729\
        );

    \I__2639\ : InMux
    port map (
            O => \N__13732\,
            I => \N__13724\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__13729\,
            I => \N__13712\
        );

    \I__2637\ : InMux
    port map (
            O => \N__13728\,
            I => \N__13709\
        );

    \I__2636\ : InMux
    port map (
            O => \N__13727\,
            I => \N__13706\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__13724\,
            I => \N__13703\
        );

    \I__2634\ : InMux
    port map (
            O => \N__13723\,
            I => \N__13696\
        );

    \I__2633\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13696\
        );

    \I__2632\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13696\
        );

    \I__2631\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13693\
        );

    \I__2630\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13684\
        );

    \I__2629\ : InMux
    port map (
            O => \N__13718\,
            I => \N__13684\
        );

    \I__2628\ : InMux
    port map (
            O => \N__13717\,
            I => \N__13684\
        );

    \I__2627\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13684\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13715\,
            I => \N__13681\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__13712\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__13709\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__13706\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__13703\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__13696\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__13693\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__13684\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__13681\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2617\ : InMux
    port map (
            O => \N__13664\,
            I => \N__13661\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__13661\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x1\
        );

    \I__2615\ : IoInMux
    port map (
            O => \N__13658\,
            I => \N__13655\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__13655\,
            I => \N__13651\
        );

    \I__2613\ : IoInMux
    port map (
            O => \N__13654\,
            I => \N__13648\
        );

    \I__2612\ : IoSpan4Mux
    port map (
            O => \N__13651\,
            I => \N__13642\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__13648\,
            I => \N__13642\
        );

    \I__2610\ : IoInMux
    port map (
            O => \N__13647\,
            I => \N__13637\
        );

    \I__2609\ : IoSpan4Mux
    port map (
            O => \N__13642\,
            I => \N__13632\
        );

    \I__2608\ : IoInMux
    port map (
            O => \N__13641\,
            I => \N__13629\
        );

    \I__2607\ : IoInMux
    port map (
            O => \N__13640\,
            I => \N__13626\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__13637\,
            I => \N__13620\
        );

    \I__2605\ : IoInMux
    port map (
            O => \N__13636\,
            I => \N__13617\
        );

    \I__2604\ : IoInMux
    port map (
            O => \N__13635\,
            I => \N__13612\
        );

    \I__2603\ : IoSpan4Mux
    port map (
            O => \N__13632\,
            I => \N__13607\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__13629\,
            I => \N__13607\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__13626\,
            I => \N__13604\
        );

    \I__2600\ : IoInMux
    port map (
            O => \N__13625\,
            I => \N__13601\
        );

    \I__2599\ : IoInMux
    port map (
            O => \N__13624\,
            I => \N__13598\
        );

    \I__2598\ : IoInMux
    port map (
            O => \N__13623\,
            I => \N__13595\
        );

    \I__2597\ : IoSpan4Mux
    port map (
            O => \N__13620\,
            I => \N__13587\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__13617\,
            I => \N__13587\
        );

    \I__2595\ : IoInMux
    port map (
            O => \N__13616\,
            I => \N__13584\
        );

    \I__2594\ : IoInMux
    port map (
            O => \N__13615\,
            I => \N__13581\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__13612\,
            I => \N__13577\
        );

    \I__2592\ : IoSpan4Mux
    port map (
            O => \N__13607\,
            I => \N__13574\
        );

    \I__2591\ : IoSpan4Mux
    port map (
            O => \N__13604\,
            I => \N__13567\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__13601\,
            I => \N__13567\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__13598\,
            I => \N__13567\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__13595\,
            I => \N__13564\
        );

    \I__2587\ : IoInMux
    port map (
            O => \N__13594\,
            I => \N__13561\
        );

    \I__2586\ : IoInMux
    port map (
            O => \N__13593\,
            I => \N__13558\
        );

    \I__2585\ : IoInMux
    port map (
            O => \N__13592\,
            I => \N__13555\
        );

    \I__2584\ : IoSpan4Mux
    port map (
            O => \N__13587\,
            I => \N__13550\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__13584\,
            I => \N__13550\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__13581\,
            I => \N__13547\
        );

    \I__2581\ : IoInMux
    port map (
            O => \N__13580\,
            I => \N__13544\
        );

    \I__2580\ : Span4Mux_s3_v
    port map (
            O => \N__13577\,
            I => \N__13541\
        );

    \I__2579\ : IoSpan4Mux
    port map (
            O => \N__13574\,
            I => \N__13536\
        );

    \I__2578\ : IoSpan4Mux
    port map (
            O => \N__13567\,
            I => \N__13536\
        );

    \I__2577\ : Span4Mux_s3_h
    port map (
            O => \N__13564\,
            I => \N__13533\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__13561\,
            I => \N__13530\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__13558\,
            I => \N__13527\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__13555\,
            I => \N__13524\
        );

    \I__2573\ : IoSpan4Mux
    port map (
            O => \N__13550\,
            I => \N__13517\
        );

    \I__2572\ : IoSpan4Mux
    port map (
            O => \N__13547\,
            I => \N__13517\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__13544\,
            I => \N__13517\
        );

    \I__2570\ : Span4Mux_v
    port map (
            O => \N__13541\,
            I => \N__13514\
        );

    \I__2569\ : Span4Mux_s3_h
    port map (
            O => \N__13536\,
            I => \N__13511\
        );

    \I__2568\ : Span4Mux_v
    port map (
            O => \N__13533\,
            I => \N__13504\
        );

    \I__2567\ : Span4Mux_s3_h
    port map (
            O => \N__13530\,
            I => \N__13504\
        );

    \I__2566\ : Span4Mux_s3_h
    port map (
            O => \N__13527\,
            I => \N__13504\
        );

    \I__2565\ : Span4Mux_s3_h
    port map (
            O => \N__13524\,
            I => \N__13501\
        );

    \I__2564\ : IoSpan4Mux
    port map (
            O => \N__13517\,
            I => \N__13498\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__13514\,
            I => \N__13490\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__13511\,
            I => \N__13490\
        );

    \I__2561\ : Span4Mux_h
    port map (
            O => \N__13504\,
            I => \N__13490\
        );

    \I__2560\ : Span4Mux_h
    port map (
            O => \N__13501\,
            I => \N__13487\
        );

    \I__2559\ : Span4Mux_s0_v
    port map (
            O => \N__13498\,
            I => \N__13484\
        );

    \I__2558\ : IoInMux
    port map (
            O => \N__13497\,
            I => \N__13481\
        );

    \I__2557\ : Span4Mux_h
    port map (
            O => \N__13490\,
            I => \N__13478\
        );

    \I__2556\ : Span4Mux_h
    port map (
            O => \N__13487\,
            I => \N__13475\
        );

    \I__2555\ : Sp12to4
    port map (
            O => \N__13484\,
            I => \N__13470\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__13481\,
            I => \N__13470\
        );

    \I__2553\ : Span4Mux_h
    port map (
            O => \N__13478\,
            I => \N__13467\
        );

    \I__2552\ : Span4Mux_h
    port map (
            O => \N__13475\,
            I => \N__13464\
        );

    \I__2551\ : Span12Mux_s6_v
    port map (
            O => \N__13470\,
            I => \N__13461\
        );

    \I__2550\ : Odrv4
    port map (
            O => \N__13467\,
            I => port_dmab_c_i
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__13464\,
            I => port_dmab_c_i
        );

    \I__2548\ : Odrv12
    port map (
            O => \N__13461\,
            I => port_dmab_c_i
        );

    \I__2547\ : InMux
    port map (
            O => \N__13454\,
            I => \N__13449\
        );

    \I__2546\ : InMux
    port map (
            O => \N__13453\,
            I => \N__13446\
        );

    \I__2545\ : InMux
    port map (
            O => \N__13452\,
            I => \N__13442\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__13449\,
            I => \N__13439\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__13446\,
            I => \N__13435\
        );

    \I__2542\ : InMux
    port map (
            O => \N__13445\,
            I => \N__13432\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__13442\,
            I => \N__13429\
        );

    \I__2540\ : Span4Mux_v
    port map (
            O => \N__13439\,
            I => \N__13419\
        );

    \I__2539\ : InMux
    port map (
            O => \N__13438\,
            I => \N__13416\
        );

    \I__2538\ : Span4Mux_h
    port map (
            O => \N__13435\,
            I => \N__13413\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__13432\,
            I => \N__13410\
        );

    \I__2536\ : Span4Mux_h
    port map (
            O => \N__13429\,
            I => \N__13407\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13428\,
            I => \N__13402\
        );

    \I__2534\ : InMux
    port map (
            O => \N__13427\,
            I => \N__13402\
        );

    \I__2533\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13397\
        );

    \I__2532\ : InMux
    port map (
            O => \N__13425\,
            I => \N__13397\
        );

    \I__2531\ : InMux
    port map (
            O => \N__13424\,
            I => \N__13392\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13423\,
            I => \N__13392\
        );

    \I__2529\ : InMux
    port map (
            O => \N__13422\,
            I => \N__13389\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__13419\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__13416\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__13413\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__13410\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2524\ : Odrv4
    port map (
            O => \N__13407\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__13402\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__13397\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__13392\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__13389\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2519\ : InMux
    port map (
            O => \N__13370\,
            I => \N__13367\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__13367\,
            I => \N__13363\
        );

    \I__2517\ : InMux
    port map (
            O => \N__13366\,
            I => \N__13360\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__13363\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__13360\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2514\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13349\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13354\,
            I => \N__13349\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__13349\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13346\,
            I => \un1_M_this_data_count_q_cry_0\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13343\,
            I => \un1_M_this_data_count_q_cry_1\
        );

    \I__2509\ : InMux
    port map (
            O => \N__13340\,
            I => \bfn_15_22_0_\
        );

    \I__2508\ : InMux
    port map (
            O => \N__13337\,
            I => \N__13326\
        );

    \I__2507\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13321\
        );

    \I__2506\ : InMux
    port map (
            O => \N__13335\,
            I => \N__13321\
        );

    \I__2505\ : InMux
    port map (
            O => \N__13334\,
            I => \N__13314\
        );

    \I__2504\ : InMux
    port map (
            O => \N__13333\,
            I => \N__13314\
        );

    \I__2503\ : InMux
    port map (
            O => \N__13332\,
            I => \N__13314\
        );

    \I__2502\ : InMux
    port map (
            O => \N__13331\,
            I => \N__13311\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13330\,
            I => \N__13306\
        );

    \I__2500\ : InMux
    port map (
            O => \N__13329\,
            I => \N__13306\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__13326\,
            I => \N__13301\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__13321\,
            I => \N__13301\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__13314\,
            I => \N__13298\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__13311\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__13306\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__13301\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2493\ : Odrv12
    port map (
            O => \N__13298\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__13289\,
            I => \N__13286\
        );

    \I__2491\ : InMux
    port map (
            O => \N__13286\,
            I => \N__13283\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__13283\,
            I => \N__13278\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13282\,
            I => \N__13275\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13272\
        );

    \I__2487\ : Span4Mux_v
    port map (
            O => \N__13278\,
            I => \N__13269\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__13275\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__13272\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__13269\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__2483\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13259\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__13259\,
            I => \N__13255\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13252\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__13255\,
            I => \N__13249\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__13252\,
            I => \N__13246\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__13249\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__13246\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__13241\,
            I => \N__13238\
        );

    \I__2475\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13235\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__13235\,
            I => \N__13232\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__13232\,
            I => \this_vga_signals.mult1_un54_sum_c2\
        );

    \I__2472\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__13226\,
            I => \N__13223\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__13223\,
            I => \N__13217\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13222\,
            I => \N__13214\
        );

    \I__2468\ : InMux
    port map (
            O => \N__13221\,
            I => \N__13209\
        );

    \I__2467\ : InMux
    port map (
            O => \N__13220\,
            I => \N__13209\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__13217\,
            I => \this_vga_signals.mult1_un47_sum_i_3\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__13214\,
            I => \this_vga_signals.mult1_un47_sum_i_3\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__13209\,
            I => \this_vga_signals.mult1_un47_sum_i_3\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13202\,
            I => \N__13185\
        );

    \I__2462\ : InMux
    port map (
            O => \N__13201\,
            I => \N__13185\
        );

    \I__2461\ : InMux
    port map (
            O => \N__13200\,
            I => \N__13185\
        );

    \I__2460\ : InMux
    port map (
            O => \N__13199\,
            I => \N__13182\
        );

    \I__2459\ : InMux
    port map (
            O => \N__13198\,
            I => \N__13178\
        );

    \I__2458\ : InMux
    port map (
            O => \N__13197\,
            I => \N__13173\
        );

    \I__2457\ : InMux
    port map (
            O => \N__13196\,
            I => \N__13173\
        );

    \I__2456\ : InMux
    port map (
            O => \N__13195\,
            I => \N__13168\
        );

    \I__2455\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13168\
        );

    \I__2454\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13165\
        );

    \I__2453\ : InMux
    port map (
            O => \N__13192\,
            I => \N__13162\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__13185\,
            I => \N__13157\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__13182\,
            I => \N__13157\
        );

    \I__2450\ : InMux
    port map (
            O => \N__13181\,
            I => \N__13154\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13178\,
            I => \N__13151\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__13173\,
            I => \N__13148\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__13168\,
            I => \N__13145\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__13165\,
            I => \N__13138\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__13162\,
            I => \N__13138\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__13157\,
            I => \N__13138\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__13154\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2442\ : Odrv12
    port map (
            O => \N__13151\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__13148\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__13145\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2439\ : Odrv4
    port map (
            O => \N__13138\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2438\ : InMux
    port map (
            O => \N__13127\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__13124\,
            I => \N__13117\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__13123\,
            I => \N__13110\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__13122\,
            I => \N__13107\
        );

    \I__2434\ : InMux
    port map (
            O => \N__13121\,
            I => \N__13104\
        );

    \I__2433\ : InMux
    port map (
            O => \N__13120\,
            I => \N__13101\
        );

    \I__2432\ : InMux
    port map (
            O => \N__13117\,
            I => \N__13098\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13093\
        );

    \I__2430\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13093\
        );

    \I__2429\ : InMux
    port map (
            O => \N__13114\,
            I => \N__13090\
        );

    \I__2428\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13087\
        );

    \I__2427\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13081\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13107\,
            I => \N__13081\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__13104\,
            I => \N__13077\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__13101\,
            I => \N__13068\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__13098\,
            I => \N__13068\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__13093\,
            I => \N__13068\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__13090\,
            I => \N__13068\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__13087\,
            I => \N__13065\
        );

    \I__2419\ : InMux
    port map (
            O => \N__13086\,
            I => \N__13062\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__13081\,
            I => \N__13059\
        );

    \I__2417\ : InMux
    port map (
            O => \N__13080\,
            I => \N__13056\
        );

    \I__2416\ : Span4Mux_h
    port map (
            O => \N__13077\,
            I => \N__13051\
        );

    \I__2415\ : Span4Mux_v
    port map (
            O => \N__13068\,
            I => \N__13051\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__13065\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__13062\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2412\ : Odrv4
    port map (
            O => \N__13059\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__13056\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__13051\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2409\ : InMux
    port map (
            O => \N__13040\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__13037\,
            I => \N__13029\
        );

    \I__2407\ : InMux
    port map (
            O => \N__13036\,
            I => \N__13022\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__13035\,
            I => \N__13014\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__13034\,
            I => \N__13011\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13033\,
            I => \N__13007\
        );

    \I__2403\ : InMux
    port map (
            O => \N__13032\,
            I => \N__12996\
        );

    \I__2402\ : InMux
    port map (
            O => \N__13029\,
            I => \N__12996\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13028\,
            I => \N__12996\
        );

    \I__2400\ : InMux
    port map (
            O => \N__13027\,
            I => \N__12996\
        );

    \I__2399\ : InMux
    port map (
            O => \N__13026\,
            I => \N__12996\
        );

    \I__2398\ : InMux
    port map (
            O => \N__13025\,
            I => \N__12993\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__13022\,
            I => \N__12990\
        );

    \I__2396\ : InMux
    port map (
            O => \N__13021\,
            I => \N__12987\
        );

    \I__2395\ : InMux
    port map (
            O => \N__13020\,
            I => \N__12984\
        );

    \I__2394\ : InMux
    port map (
            O => \N__13019\,
            I => \N__12981\
        );

    \I__2393\ : InMux
    port map (
            O => \N__13018\,
            I => \N__12976\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13017\,
            I => \N__12976\
        );

    \I__2391\ : InMux
    port map (
            O => \N__13014\,
            I => \N__12971\
        );

    \I__2390\ : InMux
    port map (
            O => \N__13011\,
            I => \N__12971\
        );

    \I__2389\ : InMux
    port map (
            O => \N__13010\,
            I => \N__12968\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__13007\,
            I => \N__12963\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__12996\,
            I => \N__12963\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__12993\,
            I => \N__12956\
        );

    \I__2385\ : Span4Mux_h
    port map (
            O => \N__12990\,
            I => \N__12956\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__12987\,
            I => \N__12956\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__12984\,
            I => \N__12947\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__12981\,
            I => \N__12947\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__12976\,
            I => \N__12947\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__12971\,
            I => \N__12947\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__12968\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2378\ : Odrv12
    port map (
            O => \N__12963\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__12956\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__12947\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2375\ : InMux
    port map (
            O => \N__12938\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__2374\ : InMux
    port map (
            O => \N__12935\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__2373\ : InMux
    port map (
            O => \N__12932\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__2372\ : InMux
    port map (
            O => \N__12929\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__2371\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12907\
        );

    \I__2370\ : InMux
    port map (
            O => \N__12925\,
            I => \N__12907\
        );

    \I__2369\ : InMux
    port map (
            O => \N__12924\,
            I => \N__12907\
        );

    \I__2368\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12907\
        );

    \I__2367\ : InMux
    port map (
            O => \N__12922\,
            I => \N__12902\
        );

    \I__2366\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12902\
        );

    \I__2365\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12897\
        );

    \I__2364\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12897\
        );

    \I__2363\ : InMux
    port map (
            O => \N__12918\,
            I => \N__12892\
        );

    \I__2362\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12889\
        );

    \I__2361\ : InMux
    port map (
            O => \N__12916\,
            I => \N__12886\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__12907\,
            I => \N__12876\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__12902\,
            I => \N__12876\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__12897\,
            I => \N__12876\
        );

    \I__2357\ : InMux
    port map (
            O => \N__12896\,
            I => \N__12873\
        );

    \I__2356\ : InMux
    port map (
            O => \N__12895\,
            I => \N__12870\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__12892\,
            I => \N__12865\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__12889\,
            I => \N__12865\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__12886\,
            I => \N__12862\
        );

    \I__2352\ : InMux
    port map (
            O => \N__12885\,
            I => \N__12857\
        );

    \I__2351\ : InMux
    port map (
            O => \N__12884\,
            I => \N__12857\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__12883\,
            I => \N__12854\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__12876\,
            I => \N__12850\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__12873\,
            I => \N__12847\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__12870\,
            I => \N__12844\
        );

    \I__2346\ : Span4Mux_h
    port map (
            O => \N__12865\,
            I => \N__12837\
        );

    \I__2345\ : Span4Mux_v
    port map (
            O => \N__12862\,
            I => \N__12837\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__12857\,
            I => \N__12837\
        );

    \I__2343\ : InMux
    port map (
            O => \N__12854\,
            I => \N__12832\
        );

    \I__2342\ : InMux
    port map (
            O => \N__12853\,
            I => \N__12832\
        );

    \I__2341\ : Span4Mux_h
    port map (
            O => \N__12850\,
            I => \N__12829\
        );

    \I__2340\ : Span12Mux_v
    port map (
            O => \N__12847\,
            I => \N__12826\
        );

    \I__2339\ : Span4Mux_v
    port map (
            O => \N__12844\,
            I => \N__12821\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__12837\,
            I => \N__12821\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__12832\,
            I => \this_vga_signals.GZ0Z_296\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__12829\,
            I => \this_vga_signals.GZ0Z_296\
        );

    \I__2335\ : Odrv12
    port map (
            O => \N__12826\,
            I => \this_vga_signals.GZ0Z_296\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__12821\,
            I => \this_vga_signals.GZ0Z_296\
        );

    \I__2333\ : InMux
    port map (
            O => \N__12812\,
            I => \bfn_15_21_0_\
        );

    \I__2332\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12802\
        );

    \I__2331\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12802\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__12807\,
            I => \N__12799\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__12802\,
            I => \N__12796\
        );

    \I__2328\ : InMux
    port map (
            O => \N__12799\,
            I => \N__12793\
        );

    \I__2327\ : Span4Mux_h
    port map (
            O => \N__12796\,
            I => \N__12788\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__12793\,
            I => \N__12788\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__12788\,
            I => \this_vga_signals.mult1_un40_sum_c3\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__12785\,
            I => \this_vga_signals.mult1_un40_sum_c3_cascade_\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__12782\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x0_cascade_\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__12779\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_ns_cascade_\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__12776\,
            I => \N__12773\
        );

    \I__2320\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12770\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__12770\,
            I => \this_vga_signals.mult1_un47_sum_axb2_0_3_1_1\
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__12767\,
            I => \N__12762\
        );

    \I__2317\ : InMux
    port map (
            O => \N__12766\,
            I => \N__12759\
        );

    \I__2316\ : InMux
    port map (
            O => \N__12765\,
            I => \N__12756\
        );

    \I__2315\ : InMux
    port map (
            O => \N__12762\,
            I => \N__12753\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__12759\,
            I => \N__12746\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__12756\,
            I => \N__12746\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__12753\,
            I => \N__12746\
        );

    \I__2311\ : Odrv12
    port map (
            O => \N__12746\,
            I => \this_vga_signals.M_hcounter_d6_0\
        );

    \I__2310\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12739\
        );

    \I__2309\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12735\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__12739\,
            I => \N__12732\
        );

    \I__2307\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12729\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__12735\,
            I => \N__12726\
        );

    \I__2305\ : Odrv12
    port map (
            O => \N__12732\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__12729\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__12726\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__12719\,
            I => \N__12714\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__12718\,
            I => \N__12709\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__12717\,
            I => \N__12706\
        );

    \I__2299\ : InMux
    port map (
            O => \N__12714\,
            I => \N__12703\
        );

    \I__2298\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12700\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__12712\,
            I => \N__12697\
        );

    \I__2296\ : InMux
    port map (
            O => \N__12709\,
            I => \N__12694\
        );

    \I__2295\ : InMux
    port map (
            O => \N__12706\,
            I => \N__12691\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__12703\,
            I => \N__12685\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__12700\,
            I => \N__12685\
        );

    \I__2292\ : InMux
    port map (
            O => \N__12697\,
            I => \N__12682\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__12694\,
            I => \N__12679\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__12691\,
            I => \N__12676\
        );

    \I__2289\ : InMux
    port map (
            O => \N__12690\,
            I => \N__12673\
        );

    \I__2288\ : Span4Mux_v
    port map (
            O => \N__12685\,
            I => \N__12668\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__12682\,
            I => \N__12668\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__12679\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__12676\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__12673\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__12668\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2282\ : InMux
    port map (
            O => \N__12659\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__2281\ : InMux
    port map (
            O => \N__12656\,
            I => \N__12653\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__12653\,
            I => \this_vga_signals.mult1_un75_sum_c2\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__12650\,
            I => \this_vga_signals.mult1_un82_sum_c3_cascade_\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__12647\,
            I => \N__12644\
        );

    \I__2277\ : CascadeBuf
    port map (
            O => \N__12644\,
            I => \N__12641\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__12641\,
            I => \N__12638\
        );

    \I__2275\ : CascadeBuf
    port map (
            O => \N__12638\,
            I => \N__12635\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__12635\,
            I => \N__12632\
        );

    \I__2273\ : CascadeBuf
    port map (
            O => \N__12632\,
            I => \N__12629\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__12629\,
            I => \N__12626\
        );

    \I__2271\ : CascadeBuf
    port map (
            O => \N__12626\,
            I => \N__12623\
        );

    \I__2270\ : CascadeMux
    port map (
            O => \N__12623\,
            I => \N__12620\
        );

    \I__2269\ : CascadeBuf
    port map (
            O => \N__12620\,
            I => \N__12617\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__12617\,
            I => \N__12614\
        );

    \I__2267\ : CascadeBuf
    port map (
            O => \N__12614\,
            I => \N__12611\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__12611\,
            I => \N__12608\
        );

    \I__2265\ : CascadeBuf
    port map (
            O => \N__12608\,
            I => \N__12605\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__12605\,
            I => \N__12602\
        );

    \I__2263\ : CascadeBuf
    port map (
            O => \N__12602\,
            I => \N__12599\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__12599\,
            I => \N__12596\
        );

    \I__2261\ : CascadeBuf
    port map (
            O => \N__12596\,
            I => \N__12593\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__12593\,
            I => \N__12590\
        );

    \I__2259\ : CascadeBuf
    port map (
            O => \N__12590\,
            I => \N__12587\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__12587\,
            I => \N__12584\
        );

    \I__2257\ : CascadeBuf
    port map (
            O => \N__12584\,
            I => \N__12581\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__12581\,
            I => \N__12578\
        );

    \I__2255\ : CascadeBuf
    port map (
            O => \N__12578\,
            I => \N__12575\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__12575\,
            I => \N__12572\
        );

    \I__2253\ : CascadeBuf
    port map (
            O => \N__12572\,
            I => \N__12569\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__12569\,
            I => \N__12566\
        );

    \I__2251\ : CascadeBuf
    port map (
            O => \N__12566\,
            I => \N__12563\
        );

    \I__2250\ : CascadeMux
    port map (
            O => \N__12563\,
            I => \N__12560\
        );

    \I__2249\ : CascadeBuf
    port map (
            O => \N__12560\,
            I => \N__12557\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__12557\,
            I => \N__12554\
        );

    \I__2247\ : InMux
    port map (
            O => \N__12554\,
            I => \N__12551\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__12551\,
            I => \N__12548\
        );

    \I__2245\ : Span4Mux_v
    port map (
            O => \N__12548\,
            I => \N__12545\
        );

    \I__2244\ : Sp12to4
    port map (
            O => \N__12545\,
            I => \N__12542\
        );

    \I__2243\ : Span12Mux_h
    port map (
            O => \N__12542\,
            I => \N__12539\
        );

    \I__2242\ : Odrv12
    port map (
            O => \N__12539\,
            I => \M_this_vga_signals_address_7\
        );

    \I__2241\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12533\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__12533\,
            I => \this_vga_signals.mult1_un68_sum_axbxc1\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__12530\,
            I => \this_vga_signals.mult1_un75_sum_c3_0_cascade_\
        );

    \I__2238\ : InMux
    port map (
            O => \N__12527\,
            I => \N__12524\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__12524\,
            I => \this_vga_signals.mult1_un82_sum_i_1_3\
        );

    \I__2236\ : InMux
    port map (
            O => \N__12521\,
            I => \N__12517\
        );

    \I__2235\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12514\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__12517\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__12514\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__12509\,
            I => \N__12506\
        );

    \I__2231\ : InMux
    port map (
            O => \N__12506\,
            I => \N__12503\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__12503\,
            I => \N__12499\
        );

    \I__2229\ : InMux
    port map (
            O => \N__12502\,
            I => \N__12496\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__12499\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0_0\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__12496\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0_0\
        );

    \I__2226\ : InMux
    port map (
            O => \N__12491\,
            I => \N__12484\
        );

    \I__2225\ : InMux
    port map (
            O => \N__12490\,
            I => \N__12481\
        );

    \I__2224\ : InMux
    port map (
            O => \N__12489\,
            I => \N__12474\
        );

    \I__2223\ : InMux
    port map (
            O => \N__12488\,
            I => \N__12474\
        );

    \I__2222\ : InMux
    port map (
            O => \N__12487\,
            I => \N__12474\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__12484\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__12481\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__12474\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__12467\,
            I => \N__12464\
        );

    \I__2217\ : CascadeBuf
    port map (
            O => \N__12464\,
            I => \N__12461\
        );

    \I__2216\ : CascadeMux
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__2215\ : CascadeBuf
    port map (
            O => \N__12458\,
            I => \N__12455\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__12455\,
            I => \N__12452\
        );

    \I__2213\ : CascadeBuf
    port map (
            O => \N__12452\,
            I => \N__12449\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__12449\,
            I => \N__12446\
        );

    \I__2211\ : CascadeBuf
    port map (
            O => \N__12446\,
            I => \N__12443\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__12443\,
            I => \N__12440\
        );

    \I__2209\ : CascadeBuf
    port map (
            O => \N__12440\,
            I => \N__12437\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__12437\,
            I => \N__12434\
        );

    \I__2207\ : CascadeBuf
    port map (
            O => \N__12434\,
            I => \N__12431\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__12431\,
            I => \N__12428\
        );

    \I__2205\ : CascadeBuf
    port map (
            O => \N__12428\,
            I => \N__12425\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__12425\,
            I => \N__12422\
        );

    \I__2203\ : CascadeBuf
    port map (
            O => \N__12422\,
            I => \N__12419\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__12419\,
            I => \N__12416\
        );

    \I__2201\ : CascadeBuf
    port map (
            O => \N__12416\,
            I => \N__12413\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__12413\,
            I => \N__12410\
        );

    \I__2199\ : CascadeBuf
    port map (
            O => \N__12410\,
            I => \N__12407\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__12407\,
            I => \N__12404\
        );

    \I__2197\ : CascadeBuf
    port map (
            O => \N__12404\,
            I => \N__12401\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__12401\,
            I => \N__12398\
        );

    \I__2195\ : CascadeBuf
    port map (
            O => \N__12398\,
            I => \N__12395\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__12395\,
            I => \N__12392\
        );

    \I__2193\ : CascadeBuf
    port map (
            O => \N__12392\,
            I => \N__12389\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__12389\,
            I => \N__12386\
        );

    \I__2191\ : CascadeBuf
    port map (
            O => \N__12386\,
            I => \N__12383\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__12383\,
            I => \N__12380\
        );

    \I__2189\ : CascadeBuf
    port map (
            O => \N__12380\,
            I => \N__12377\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__12377\,
            I => \N__12374\
        );

    \I__2187\ : InMux
    port map (
            O => \N__12374\,
            I => \N__12371\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__12371\,
            I => \N__12368\
        );

    \I__2185\ : Span4Mux_s2_v
    port map (
            O => \N__12368\,
            I => \N__12365\
        );

    \I__2184\ : Span4Mux_v
    port map (
            O => \N__12365\,
            I => \N__12362\
        );

    \I__2183\ : Sp12to4
    port map (
            O => \N__12362\,
            I => \N__12359\
        );

    \I__2182\ : Span12Mux_h
    port map (
            O => \N__12359\,
            I => \N__12356\
        );

    \I__2181\ : Odrv12
    port map (
            O => \N__12356\,
            I => \M_this_vga_signals_address_10\
        );

    \I__2180\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12350\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__12350\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_bm\
        );

    \I__2178\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12343\
        );

    \I__2177\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12340\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__12343\,
            I => \this_vga_signals.mult1_un61_sum_axb2\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__12340\,
            I => \this_vga_signals.mult1_un61_sum_axb2\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__12335\,
            I => \N__12332\
        );

    \I__2173\ : InMux
    port map (
            O => \N__12332\,
            I => \N__12325\
        );

    \I__2172\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12325\
        );

    \I__2171\ : InMux
    port map (
            O => \N__12330\,
            I => \N__12322\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12325\,
            I => \this_vga_signals.mult1_un61_sum_c2\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__12322\,
            I => \this_vga_signals.mult1_un61_sum_c2\
        );

    \I__2168\ : InMux
    port map (
            O => \N__12317\,
            I => \N__12314\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__12314\,
            I => \this_vga_signals.if_N_10\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__12311\,
            I => \N__12308\
        );

    \I__2165\ : CascadeBuf
    port map (
            O => \N__12308\,
            I => \N__12305\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__12305\,
            I => \N__12302\
        );

    \I__2163\ : CascadeBuf
    port map (
            O => \N__12302\,
            I => \N__12299\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__12299\,
            I => \N__12296\
        );

    \I__2161\ : CascadeBuf
    port map (
            O => \N__12296\,
            I => \N__12293\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__12293\,
            I => \N__12290\
        );

    \I__2159\ : CascadeBuf
    port map (
            O => \N__12290\,
            I => \N__12287\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__12287\,
            I => \N__12284\
        );

    \I__2157\ : CascadeBuf
    port map (
            O => \N__12284\,
            I => \N__12281\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__12281\,
            I => \N__12278\
        );

    \I__2155\ : CascadeBuf
    port map (
            O => \N__12278\,
            I => \N__12275\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__12275\,
            I => \N__12272\
        );

    \I__2153\ : CascadeBuf
    port map (
            O => \N__12272\,
            I => \N__12269\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__12269\,
            I => \N__12266\
        );

    \I__2151\ : CascadeBuf
    port map (
            O => \N__12266\,
            I => \N__12263\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__12263\,
            I => \N__12260\
        );

    \I__2149\ : CascadeBuf
    port map (
            O => \N__12260\,
            I => \N__12257\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__12257\,
            I => \N__12254\
        );

    \I__2147\ : CascadeBuf
    port map (
            O => \N__12254\,
            I => \N__12251\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__12251\,
            I => \N__12248\
        );

    \I__2145\ : CascadeBuf
    port map (
            O => \N__12248\,
            I => \N__12245\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__12245\,
            I => \N__12242\
        );

    \I__2143\ : CascadeBuf
    port map (
            O => \N__12242\,
            I => \N__12239\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__12239\,
            I => \N__12236\
        );

    \I__2141\ : CascadeBuf
    port map (
            O => \N__12236\,
            I => \N__12233\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__12233\,
            I => \N__12230\
        );

    \I__2139\ : CascadeBuf
    port map (
            O => \N__12230\,
            I => \N__12227\
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__12227\,
            I => \N__12224\
        );

    \I__2137\ : CascadeBuf
    port map (
            O => \N__12224\,
            I => \N__12221\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__12221\,
            I => \N__12218\
        );

    \I__2135\ : InMux
    port map (
            O => \N__12218\,
            I => \N__12215\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__12215\,
            I => \N__12212\
        );

    \I__2133\ : Span4Mux_s3_v
    port map (
            O => \N__12212\,
            I => \N__12209\
        );

    \I__2132\ : Sp12to4
    port map (
            O => \N__12209\,
            I => \N__12206\
        );

    \I__2131\ : Span12Mux_h
    port map (
            O => \N__12206\,
            I => \N__12203\
        );

    \I__2130\ : Odrv12
    port map (
            O => \N__12203\,
            I => \M_this_vga_signals_address_9\
        );

    \I__2129\ : InMux
    port map (
            O => \N__12200\,
            I => \N__12194\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12194\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__12194\,
            I => \this_vga_signals.mult1_un68_sum_axbxc2_0\
        );

    \I__2126\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12183\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12176\
        );

    \I__2124\ : InMux
    port map (
            O => \N__12189\,
            I => \N__12176\
        );

    \I__2123\ : InMux
    port map (
            O => \N__12188\,
            I => \N__12176\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12187\,
            I => \N__12171\
        );

    \I__2121\ : InMux
    port map (
            O => \N__12186\,
            I => \N__12171\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__12183\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__12176\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__12171\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0\
        );

    \I__2117\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12161\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__12161\,
            I => \this_vga_signals.mult1_un68_sum_axbxc2\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12158\,
            I => \N__12155\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__12155\,
            I => \this_vga_signals.mult1_un75_sum_c3_0\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__12152\,
            I => \this_vga_signals.mult1_un68_sum_axbxc2_cascade_\
        );

    \I__2112\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12144\
        );

    \I__2111\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12141\
        );

    \I__2110\ : InMux
    port map (
            O => \N__12147\,
            I => \N__12138\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__12144\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_0\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__12141\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_0\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__12138\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_0\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__12131\,
            I => \N__12128\
        );

    \I__2105\ : CascadeBuf
    port map (
            O => \N__12128\,
            I => \N__12125\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__12125\,
            I => \N__12122\
        );

    \I__2103\ : CascadeBuf
    port map (
            O => \N__12122\,
            I => \N__12119\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__12119\,
            I => \N__12116\
        );

    \I__2101\ : CascadeBuf
    port map (
            O => \N__12116\,
            I => \N__12113\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__12113\,
            I => \N__12110\
        );

    \I__2099\ : CascadeBuf
    port map (
            O => \N__12110\,
            I => \N__12107\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__12107\,
            I => \N__12104\
        );

    \I__2097\ : CascadeBuf
    port map (
            O => \N__12104\,
            I => \N__12101\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__12101\,
            I => \N__12098\
        );

    \I__2095\ : CascadeBuf
    port map (
            O => \N__12098\,
            I => \N__12095\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__2093\ : CascadeBuf
    port map (
            O => \N__12092\,
            I => \N__12089\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__12089\,
            I => \N__12086\
        );

    \I__2091\ : CascadeBuf
    port map (
            O => \N__12086\,
            I => \N__12083\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__12083\,
            I => \N__12080\
        );

    \I__2089\ : CascadeBuf
    port map (
            O => \N__12080\,
            I => \N__12077\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__12077\,
            I => \N__12074\
        );

    \I__2087\ : CascadeBuf
    port map (
            O => \N__12074\,
            I => \N__12071\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__12071\,
            I => \N__12068\
        );

    \I__2085\ : CascadeBuf
    port map (
            O => \N__12068\,
            I => \N__12065\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__12065\,
            I => \N__12062\
        );

    \I__2083\ : CascadeBuf
    port map (
            O => \N__12062\,
            I => \N__12059\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__12059\,
            I => \N__12056\
        );

    \I__2081\ : CascadeBuf
    port map (
            O => \N__12056\,
            I => \N__12053\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__12053\,
            I => \N__12050\
        );

    \I__2079\ : CascadeBuf
    port map (
            O => \N__12050\,
            I => \N__12047\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__12047\,
            I => \N__12044\
        );

    \I__2077\ : CascadeBuf
    port map (
            O => \N__12044\,
            I => \N__12041\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__12041\,
            I => \N__12038\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12038\,
            I => \N__12035\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__12035\,
            I => \N__12032\
        );

    \I__2073\ : Span4Mux_h
    port map (
            O => \N__12032\,
            I => \N__12029\
        );

    \I__2072\ : Span4Mux_h
    port map (
            O => \N__12029\,
            I => \N__12026\
        );

    \I__2071\ : Sp12to4
    port map (
            O => \N__12026\,
            I => \N__12023\
        );

    \I__2070\ : Span12Mux_v
    port map (
            O => \N__12023\,
            I => \N__12020\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__12020\,
            I => \M_this_vga_signals_address_8\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__12017\,
            I => \this_vga_signals.M_vcounter_d7lt9_cascade_\
        );

    \I__2067\ : InMux
    port map (
            O => \N__12014\,
            I => \N__12011\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__12011\,
            I => \this_vga_signals.M_vcounter_d7lto8_1\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__12008\,
            I => \this_vga_signals.un6_vvisibilitylt9_0_cascade_\
        );

    \I__2064\ : InMux
    port map (
            O => \N__12005\,
            I => \N__12001\
        );

    \I__2063\ : InMux
    port map (
            O => \N__12004\,
            I => \N__11998\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__12001\,
            I => \this_vga_signals.vaddress_c5_i\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__11998\,
            I => \this_vga_signals.vaddress_c5_i\
        );

    \I__2060\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11990\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__11990\,
            I => \N__11985\
        );

    \I__2058\ : InMux
    port map (
            O => \N__11989\,
            I => \N__11982\
        );

    \I__2057\ : InMux
    port map (
            O => \N__11988\,
            I => \N__11979\
        );

    \I__2056\ : Span4Mux_h
    port map (
            O => \N__11985\,
            I => \N__11976\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__11982\,
            I => \N__11973\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__11979\,
            I => \N__11969\
        );

    \I__2053\ : Span4Mux_v
    port map (
            O => \N__11976\,
            I => \N__11964\
        );

    \I__2052\ : Span4Mux_v
    port map (
            O => \N__11973\,
            I => \N__11964\
        );

    \I__2051\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11961\
        );

    \I__2050\ : Span12Mux_h
    port map (
            O => \N__11969\,
            I => \N__11958\
        );

    \I__2049\ : Span4Mux_h
    port map (
            O => \N__11964\,
            I => \N__11953\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__11961\,
            I => \N__11953\
        );

    \I__2047\ : Odrv12
    port map (
            O => \N__11958\,
            I => \this_vga_signals.vvisibility\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__11953\,
            I => \this_vga_signals.vvisibility\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__11948\,
            I => \this_vga_signals.vsync_1_0_cascade_\
        );

    \I__2044\ : InMux
    port map (
            O => \N__11945\,
            I => \N__11942\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__11942\,
            I => \this_vga_signals.vsync_1_4\
        );

    \I__2042\ : InMux
    port map (
            O => \N__11939\,
            I => \N__11936\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__11936\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_ns_1\
        );

    \I__2040\ : InMux
    port map (
            O => \N__11933\,
            I => \N__11924\
        );

    \I__2039\ : InMux
    port map (
            O => \N__11932\,
            I => \N__11924\
        );

    \I__2038\ : InMux
    port map (
            O => \N__11931\,
            I => \N__11924\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__11924\,
            I => \N__11921\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__11921\,
            I => \this_vga_signals.SUM_2\
        );

    \I__2035\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11915\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__11915\,
            I => \this_vga_signals.mult1_un47_sum_c2\
        );

    \I__2033\ : InMux
    port map (
            O => \N__11912\,
            I => \N__11908\
        );

    \I__2032\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11905\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__11908\,
            I => \this_vga_signals.mult1_un47_sum_axb2_0_3\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__11905\,
            I => \this_vga_signals.mult1_un47_sum_axb2_0_3\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__11900\,
            I => \this_vga_signals.mult1_un47_sum_c2_cascade_\
        );

    \I__2028\ : InMux
    port map (
            O => \N__11897\,
            I => \N__11891\
        );

    \I__2027\ : InMux
    port map (
            O => \N__11896\,
            I => \N__11891\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__11891\,
            I => \N__11888\
        );

    \I__2025\ : Odrv4
    port map (
            O => \N__11888\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2024\ : InMux
    port map (
            O => \N__11885\,
            I => \N__11882\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__11882\,
            I => \this_vga_signals.mult1_un47_sum_axb2_3_tz\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__11879\,
            I => \N__11875\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__11878\,
            I => \N__11872\
        );

    \I__2020\ : InMux
    port map (
            O => \N__11875\,
            I => \N__11863\
        );

    \I__2019\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11863\
        );

    \I__2018\ : InMux
    port map (
            O => \N__11871\,
            I => \N__11863\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__11870\,
            I => \N__11860\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__11863\,
            I => \N__11857\
        );

    \I__2015\ : InMux
    port map (
            O => \N__11860\,
            I => \N__11854\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__11857\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__11854\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__11849\,
            I => \this_vga_signals.M_vcounter_d7lt8_0_cascade_\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__11846\,
            I => \this_vga_signals.mult1_un54_sum_c2_cascade_\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__11843\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__11840\,
            I => \this_vga_signals.mult1_un61_sum_c2_cascade_\
        );

    \I__2008\ : InMux
    port map (
            O => \N__11837\,
            I => \N__11832\
        );

    \I__2007\ : InMux
    port map (
            O => \N__11836\,
            I => \N__11827\
        );

    \I__2006\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11827\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__11832\,
            I => \this_vga_signals.mult1_un54_sum_axb1_i\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__11827\,
            I => \this_vga_signals.mult1_un54_sum_axb1_i\
        );

    \I__2003\ : InMux
    port map (
            O => \N__11822\,
            I => \N__11818\
        );

    \I__2002\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11815\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__11818\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1_2\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__11815\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1_2\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__11810\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1_2_cascade_\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__11807\,
            I => \N__11804\
        );

    \I__1997\ : InMux
    port map (
            O => \N__11804\,
            I => \N__11799\
        );

    \I__1996\ : InMux
    port map (
            O => \N__11803\,
            I => \N__11794\
        );

    \I__1995\ : InMux
    port map (
            O => \N__11802\,
            I => \N__11794\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__11799\,
            I => \this_vga_signals.mult1_un40_sum_c2\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__11794\,
            I => \this_vga_signals.mult1_un40_sum_c2\
        );

    \I__1992\ : InMux
    port map (
            O => \N__11789\,
            I => \N__11785\
        );

    \I__1991\ : InMux
    port map (
            O => \N__11788\,
            I => \N__11782\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__11785\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__11782\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__11777\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0_cascade_\
        );

    \I__1987\ : InMux
    port map (
            O => \N__11774\,
            I => \N__11769\
        );

    \I__1986\ : InMux
    port map (
            O => \N__11773\,
            I => \N__11764\
        );

    \I__1985\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11764\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__11769\,
            I => \this_vga_signals.mult1_un47_sum_ac0_4\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__11764\,
            I => \this_vga_signals.mult1_un47_sum_ac0_4\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__11759\,
            I => \N__11756\
        );

    \I__1981\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11753\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__11753\,
            I => \this_vga_signals.un2_vsynclt8\
        );

    \I__1979\ : IoInMux
    port map (
            O => \N__11750\,
            I => \N__11747\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__11747\,
            I => \N__11744\
        );

    \I__1977\ : Span4Mux_s0_v
    port map (
            O => \N__11744\,
            I => \N__11741\
        );

    \I__1976\ : Sp12to4
    port map (
            O => \N__11741\,
            I => \N__11738\
        );

    \I__1975\ : Span12Mux_h
    port map (
            O => \N__11738\,
            I => \N__11735\
        );

    \I__1974\ : Odrv12
    port map (
            O => \N__11735\,
            I => this_vga_signals_vsync_1_i
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__11732\,
            I => \N__11729\
        );

    \I__1972\ : CascadeBuf
    port map (
            O => \N__11729\,
            I => \N__11726\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__11726\,
            I => \N__11723\
        );

    \I__1970\ : CascadeBuf
    port map (
            O => \N__11723\,
            I => \N__11720\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__11720\,
            I => \N__11717\
        );

    \I__1968\ : CascadeBuf
    port map (
            O => \N__11717\,
            I => \N__11714\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__11714\,
            I => \N__11711\
        );

    \I__1966\ : CascadeBuf
    port map (
            O => \N__11711\,
            I => \N__11708\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__11708\,
            I => \N__11705\
        );

    \I__1964\ : CascadeBuf
    port map (
            O => \N__11705\,
            I => \N__11702\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__11702\,
            I => \N__11699\
        );

    \I__1962\ : CascadeBuf
    port map (
            O => \N__11699\,
            I => \N__11696\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__11696\,
            I => \N__11693\
        );

    \I__1960\ : CascadeBuf
    port map (
            O => \N__11693\,
            I => \N__11690\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__11690\,
            I => \N__11687\
        );

    \I__1958\ : CascadeBuf
    port map (
            O => \N__11687\,
            I => \N__11684\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__11684\,
            I => \N__11681\
        );

    \I__1956\ : CascadeBuf
    port map (
            O => \N__11681\,
            I => \N__11678\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__11678\,
            I => \N__11675\
        );

    \I__1954\ : CascadeBuf
    port map (
            O => \N__11675\,
            I => \N__11672\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__11672\,
            I => \N__11669\
        );

    \I__1952\ : CascadeBuf
    port map (
            O => \N__11669\,
            I => \N__11666\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__11666\,
            I => \N__11663\
        );

    \I__1950\ : CascadeBuf
    port map (
            O => \N__11663\,
            I => \N__11660\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__11660\,
            I => \N__11657\
        );

    \I__1948\ : CascadeBuf
    port map (
            O => \N__11657\,
            I => \N__11654\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__11654\,
            I => \N__11651\
        );

    \I__1946\ : CascadeBuf
    port map (
            O => \N__11651\,
            I => \N__11648\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__11648\,
            I => \N__11645\
        );

    \I__1944\ : CascadeBuf
    port map (
            O => \N__11645\,
            I => \N__11642\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__11642\,
            I => \N__11639\
        );

    \I__1942\ : InMux
    port map (
            O => \N__11639\,
            I => \N__11636\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__11636\,
            I => \N__11633\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__11633\,
            I => \N__11630\
        );

    \I__1939\ : Sp12to4
    port map (
            O => \N__11630\,
            I => \N__11627\
        );

    \I__1938\ : Span12Mux_h
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__1937\ : Odrv12
    port map (
            O => \N__11624\,
            I => \M_this_vga_signals_address_6\
        );

    \I__1936\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11618\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__11618\,
            I => \this_vga_signals.if_N_9\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__11615\,
            I => \this_vga_signals.if_N_10_cascade_\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__11612\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_0_cascade_\
        );

    \I__1932\ : IoInMux
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__11606\,
            I => \N__11603\
        );

    \I__1930\ : IoSpan4Mux
    port map (
            O => \N__11603\,
            I => \N__11598\
        );

    \I__1929\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11595\
        );

    \I__1928\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11592\
        );

    \I__1927\ : Span4Mux_s2_v
    port map (
            O => \N__11598\,
            I => \N__11589\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__11595\,
            I => \N__11586\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__11592\,
            I => \N__11583\
        );

    \I__1924\ : Sp12to4
    port map (
            O => \N__11589\,
            I => \N__11580\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__11586\,
            I => \N__11577\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__11583\,
            I => \N__11574\
        );

    \I__1921\ : Span12Mux_v
    port map (
            O => \N__11580\,
            I => \N__11570\
        );

    \I__1920\ : Span4Mux_h
    port map (
            O => \N__11577\,
            I => \N__11565\
        );

    \I__1919\ : Span4Mux_h
    port map (
            O => \N__11574\,
            I => \N__11565\
        );

    \I__1918\ : InMux
    port map (
            O => \N__11573\,
            I => \N__11562\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__11570\,
            I => debug_c_1
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__11565\,
            I => debug_c_1
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__11562\,
            I => debug_c_1
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__11555\,
            I => \N__11551\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__11554\,
            I => \N__11545\
        );

    \I__1912\ : InMux
    port map (
            O => \N__11551\,
            I => \N__11542\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__11550\,
            I => \N__11538\
        );

    \I__1910\ : InMux
    port map (
            O => \N__11549\,
            I => \N__11535\
        );

    \I__1909\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11532\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11529\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__11542\,
            I => \N__11525\
        );

    \I__1906\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11522\
        );

    \I__1905\ : InMux
    port map (
            O => \N__11538\,
            I => \N__11519\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__11535\,
            I => \N__11514\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__11532\,
            I => \N__11514\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__11529\,
            I => \N__11510\
        );

    \I__1901\ : InMux
    port map (
            O => \N__11528\,
            I => \N__11507\
        );

    \I__1900\ : Span4Mux_v
    port map (
            O => \N__11525\,
            I => \N__11498\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__11522\,
            I => \N__11498\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__11519\,
            I => \N__11498\
        );

    \I__1897\ : Span4Mux_h
    port map (
            O => \N__11514\,
            I => \N__11498\
        );

    \I__1896\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11495\
        );

    \I__1895\ : Span4Mux_h
    port map (
            O => \N__11510\,
            I => \N__11492\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__11507\,
            I => \N__11487\
        );

    \I__1893\ : Span4Mux_h
    port map (
            O => \N__11498\,
            I => \N__11487\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__11495\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__11492\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__11487\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__11480\,
            I => \N__11477\
        );

    \I__1888\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11472\
        );

    \I__1887\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11464\
        );

    \I__1886\ : InMux
    port map (
            O => \N__11475\,
            I => \N__11461\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__11472\,
            I => \N__11458\
        );

    \I__1884\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11455\
        );

    \I__1883\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11452\
        );

    \I__1882\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11447\
        );

    \I__1881\ : InMux
    port map (
            O => \N__11468\,
            I => \N__11447\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__11467\,
            I => \N__11442\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__11464\,
            I => \N__11436\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__11461\,
            I => \N__11436\
        );

    \I__1877\ : Span4Mux_h
    port map (
            O => \N__11458\,
            I => \N__11431\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__11455\,
            I => \N__11431\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__11452\,
            I => \N__11428\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__11447\,
            I => \N__11425\
        );

    \I__1873\ : InMux
    port map (
            O => \N__11446\,
            I => \N__11422\
        );

    \I__1872\ : InMux
    port map (
            O => \N__11445\,
            I => \N__11419\
        );

    \I__1871\ : InMux
    port map (
            O => \N__11442\,
            I => \N__11415\
        );

    \I__1870\ : InMux
    port map (
            O => \N__11441\,
            I => \N__11412\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__11436\,
            I => \N__11409\
        );

    \I__1868\ : Span4Mux_h
    port map (
            O => \N__11431\,
            I => \N__11406\
        );

    \I__1867\ : Span4Mux_h
    port map (
            O => \N__11428\,
            I => \N__11397\
        );

    \I__1866\ : Span4Mux_h
    port map (
            O => \N__11425\,
            I => \N__11397\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__11422\,
            I => \N__11397\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__11419\,
            I => \N__11397\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11418\,
            I => \N__11394\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__11415\,
            I => \N__11391\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__11412\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__11409\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__11406\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__11397\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__11394\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__11391\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1855\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11375\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__11375\,
            I => \this_vga_signals.g0_0_a2_1\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11372\,
            I => \N__11369\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__11369\,
            I => \N__11366\
        );

    \I__1851\ : Span4Mux_v
    port map (
            O => \N__11366\,
            I => \N__11363\
        );

    \I__1850\ : Sp12to4
    port map (
            O => \N__11363\,
            I => \N__11360\
        );

    \I__1849\ : Odrv12
    port map (
            O => \N__11360\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11354\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__11354\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__11351\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0_0_cascade_\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__11348\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_cascade_\
        );

    \I__1844\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11342\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__11342\,
            I => \N__11330\
        );

    \I__1842\ : SRMux
    port map (
            O => \N__11341\,
            I => \N__11309\
        );

    \I__1841\ : SRMux
    port map (
            O => \N__11340\,
            I => \N__11309\
        );

    \I__1840\ : SRMux
    port map (
            O => \N__11339\,
            I => \N__11309\
        );

    \I__1839\ : SRMux
    port map (
            O => \N__11338\,
            I => \N__11309\
        );

    \I__1838\ : SRMux
    port map (
            O => \N__11337\,
            I => \N__11309\
        );

    \I__1837\ : SRMux
    port map (
            O => \N__11336\,
            I => \N__11309\
        );

    \I__1836\ : SRMux
    port map (
            O => \N__11335\,
            I => \N__11309\
        );

    \I__1835\ : SRMux
    port map (
            O => \N__11334\,
            I => \N__11309\
        );

    \I__1834\ : SRMux
    port map (
            O => \N__11333\,
            I => \N__11309\
        );

    \I__1833\ : Glb2LocalMux
    port map (
            O => \N__11330\,
            I => \N__11309\
        );

    \I__1832\ : GlobalMux
    port map (
            O => \N__11309\,
            I => \N__11306\
        );

    \I__1831\ : gio2CtrlBuf
    port map (
            O => \N__11306\,
            I => \this_vga_signals.N_583_g\
        );

    \I__1830\ : InMux
    port map (
            O => \N__11303\,
            I => \N__11298\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11302\,
            I => \N__11295\
        );

    \I__1828\ : InMux
    port map (
            O => \N__11301\,
            I => \N__11292\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__11298\,
            I => \N__11289\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__11295\,
            I => \N__11284\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__11292\,
            I => \N__11284\
        );

    \I__1824\ : Sp12to4
    port map (
            O => \N__11289\,
            I => \N__11281\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__11284\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRDZ0\
        );

    \I__1822\ : Odrv12
    port map (
            O => \N__11281\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRDZ0\
        );

    \I__1821\ : InMux
    port map (
            O => \N__11276\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__1820\ : InMux
    port map (
            O => \N__11273\,
            I => \N__11268\
        );

    \I__1819\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11263\
        );

    \I__1818\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11263\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__11268\,
            I => \N__11260\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11263\,
            I => \N__11257\
        );

    \I__1815\ : Span4Mux_h
    port map (
            O => \N__11260\,
            I => \N__11254\
        );

    \I__1814\ : Span4Mux_h
    port map (
            O => \N__11257\,
            I => \N__11251\
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__11254\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__11251\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0\
        );

    \I__1811\ : InMux
    port map (
            O => \N__11246\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__1810\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11236\
        );

    \I__1809\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11236\
        );

    \I__1808\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11233\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__11236\,
            I => \N__11228\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__11233\,
            I => \N__11228\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__11228\,
            I => \N__11225\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__11225\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0\
        );

    \I__1803\ : InMux
    port map (
            O => \N__11222\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__1802\ : InMux
    port map (
            O => \N__11219\,
            I => \N__11214\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11211\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11217\,
            I => \N__11208\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__11214\,
            I => \N__11205\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__11211\,
            I => \N__11202\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__11208\,
            I => \N__11199\
        );

    \I__1796\ : Span4Mux_h
    port map (
            O => \N__11205\,
            I => \N__11196\
        );

    \I__1795\ : Span4Mux_v
    port map (
            O => \N__11202\,
            I => \N__11191\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__11199\,
            I => \N__11191\
        );

    \I__1793\ : Odrv4
    port map (
            O => \N__11196\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__11191\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11186\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11183\,
            I => \bfn_12_21_0_\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11180\,
            I => \N__11175\
        );

    \I__1788\ : InMux
    port map (
            O => \N__11179\,
            I => \N__11172\
        );

    \I__1787\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11169\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__11175\,
            I => \N__11164\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__11172\,
            I => \N__11164\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__11169\,
            I => \N__11161\
        );

    \I__1783\ : Span4Mux_h
    port map (
            O => \N__11164\,
            I => \N__11158\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__11161\,
            I => \N__11155\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__11158\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__11155\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__11150\,
            I => \N__11145\
        );

    \I__1778\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11139\
        );

    \I__1777\ : InMux
    port map (
            O => \N__11148\,
            I => \N__11136\
        );

    \I__1776\ : InMux
    port map (
            O => \N__11145\,
            I => \N__11133\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__11144\,
            I => \N__11128\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__11143\,
            I => \N__11125\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__11142\,
            I => \N__11119\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__11139\,
            I => \N__11111\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__11136\,
            I => \N__11111\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__11133\,
            I => \N__11107\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11100\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11100\
        );

    \I__1767\ : InMux
    port map (
            O => \N__11128\,
            I => \N__11100\
        );

    \I__1766\ : InMux
    port map (
            O => \N__11125\,
            I => \N__11097\
        );

    \I__1765\ : InMux
    port map (
            O => \N__11124\,
            I => \N__11094\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__11123\,
            I => \N__11089\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11081\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11072\
        );

    \I__1761\ : InMux
    port map (
            O => \N__11118\,
            I => \N__11072\
        );

    \I__1760\ : InMux
    port map (
            O => \N__11117\,
            I => \N__11072\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11072\
        );

    \I__1758\ : Span4Mux_v
    port map (
            O => \N__11111\,
            I => \N__11069\
        );

    \I__1757\ : InMux
    port map (
            O => \N__11110\,
            I => \N__11066\
        );

    \I__1756\ : Span4Mux_h
    port map (
            O => \N__11107\,
            I => \N__11061\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__11100\,
            I => \N__11061\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__11097\,
            I => \N__11058\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__11094\,
            I => \N__11055\
        );

    \I__1752\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11050\
        );

    \I__1751\ : InMux
    port map (
            O => \N__11092\,
            I => \N__11050\
        );

    \I__1750\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11047\
        );

    \I__1749\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11042\
        );

    \I__1748\ : InMux
    port map (
            O => \N__11087\,
            I => \N__11042\
        );

    \I__1747\ : InMux
    port map (
            O => \N__11086\,
            I => \N__11037\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11085\,
            I => \N__11037\
        );

    \I__1745\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11034\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__11081\,
            I => \N__11027\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__11072\,
            I => \N__11027\
        );

    \I__1742\ : Span4Mux_h
    port map (
            O => \N__11069\,
            I => \N__11027\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__11066\,
            I => \N__11022\
        );

    \I__1740\ : Span4Mux_h
    port map (
            O => \N__11061\,
            I => \N__11022\
        );

    \I__1739\ : Span4Mux_v
    port map (
            O => \N__11058\,
            I => \N__11013\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__11055\,
            I => \N__11013\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__11050\,
            I => \N__11013\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11047\,
            I => \N__11013\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__11042\,
            I => \N__11010\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__11037\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__11034\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__11027\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__11022\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1730\ : Odrv4
    port map (
            O => \N__11013\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__11010\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__10997\,
            I => \N__10993\
        );

    \I__1727\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10987\
        );

    \I__1726\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10984\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__10992\,
            I => \N__10976\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__10991\,
            I => \N__10969\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__10990\,
            I => \N__10966\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__10987\,
            I => \N__10958\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__10984\,
            I => \N__10958\
        );

    \I__1720\ : InMux
    port map (
            O => \N__10983\,
            I => \N__10955\
        );

    \I__1719\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10952\
        );

    \I__1718\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10949\
        );

    \I__1717\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10946\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__10979\,
            I => \N__10942\
        );

    \I__1715\ : InMux
    port map (
            O => \N__10976\,
            I => \N__10939\
        );

    \I__1714\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10936\
        );

    \I__1713\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10933\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__10973\,
            I => \N__10928\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__10972\,
            I => \N__10925\
        );

    \I__1710\ : InMux
    port map (
            O => \N__10969\,
            I => \N__10916\
        );

    \I__1709\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10916\
        );

    \I__1708\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10916\
        );

    \I__1707\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10911\
        );

    \I__1706\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10911\
        );

    \I__1705\ : Span4Mux_h
    port map (
            O => \N__10958\,
            I => \N__10899\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__10955\,
            I => \N__10899\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__10952\,
            I => \N__10899\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__10949\,
            I => \N__10894\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__10946\,
            I => \N__10894\
        );

    \I__1700\ : InMux
    port map (
            O => \N__10945\,
            I => \N__10889\
        );

    \I__1699\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10889\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__10939\,
            I => \N__10886\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__10936\,
            I => \N__10883\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__10933\,
            I => \N__10880\
        );

    \I__1695\ : InMux
    port map (
            O => \N__10932\,
            I => \N__10877\
        );

    \I__1694\ : InMux
    port map (
            O => \N__10931\,
            I => \N__10874\
        );

    \I__1693\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10867\
        );

    \I__1692\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10867\
        );

    \I__1691\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10867\
        );

    \I__1690\ : InMux
    port map (
            O => \N__10923\,
            I => \N__10864\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__10916\,
            I => \N__10861\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__10911\,
            I => \N__10858\
        );

    \I__1687\ : InMux
    port map (
            O => \N__10910\,
            I => \N__10855\
        );

    \I__1686\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10852\
        );

    \I__1685\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10847\
        );

    \I__1684\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10847\
        );

    \I__1683\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10844\
        );

    \I__1682\ : Span4Mux_h
    port map (
            O => \N__10899\,
            I => \N__10841\
        );

    \I__1681\ : Span4Mux_v
    port map (
            O => \N__10894\,
            I => \N__10834\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__10889\,
            I => \N__10834\
        );

    \I__1679\ : Span4Mux_h
    port map (
            O => \N__10886\,
            I => \N__10834\
        );

    \I__1678\ : Span4Mux_h
    port map (
            O => \N__10883\,
            I => \N__10831\
        );

    \I__1677\ : Span4Mux_v
    port map (
            O => \N__10880\,
            I => \N__10826\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__10877\,
            I => \N__10826\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__10874\,
            I => \N__10821\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__10867\,
            I => \N__10821\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__10864\,
            I => \N__10814\
        );

    \I__1672\ : Span4Mux_h
    port map (
            O => \N__10861\,
            I => \N__10814\
        );

    \I__1671\ : Span4Mux_h
    port map (
            O => \N__10858\,
            I => \N__10814\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__10855\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__10852\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__10847\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__10844\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__10841\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__10834\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__10831\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__10826\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__10821\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__10814\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__10793\,
            I => \N__10790\
        );

    \I__1659\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10787\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__10787\,
            I => \this_vga_signals.g0_4_0\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__10784\,
            I => \N__10781\
        );

    \I__1656\ : CascadeBuf
    port map (
            O => \N__10781\,
            I => \N__10778\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__1654\ : CascadeBuf
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__10772\,
            I => \N__10769\
        );

    \I__1652\ : CascadeBuf
    port map (
            O => \N__10769\,
            I => \N__10766\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__10766\,
            I => \N__10763\
        );

    \I__1650\ : CascadeBuf
    port map (
            O => \N__10763\,
            I => \N__10760\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__10760\,
            I => \N__10757\
        );

    \I__1648\ : CascadeBuf
    port map (
            O => \N__10757\,
            I => \N__10754\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__10754\,
            I => \N__10751\
        );

    \I__1646\ : CascadeBuf
    port map (
            O => \N__10751\,
            I => \N__10748\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__10748\,
            I => \N__10745\
        );

    \I__1644\ : CascadeBuf
    port map (
            O => \N__10745\,
            I => \N__10742\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__1642\ : CascadeBuf
    port map (
            O => \N__10739\,
            I => \N__10736\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__10736\,
            I => \N__10733\
        );

    \I__1640\ : CascadeBuf
    port map (
            O => \N__10733\,
            I => \N__10730\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__10730\,
            I => \N__10727\
        );

    \I__1638\ : CascadeBuf
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__10724\,
            I => \N__10721\
        );

    \I__1636\ : CascadeBuf
    port map (
            O => \N__10721\,
            I => \N__10718\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__10718\,
            I => \N__10715\
        );

    \I__1634\ : CascadeBuf
    port map (
            O => \N__10715\,
            I => \N__10712\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__10712\,
            I => \N__10709\
        );

    \I__1632\ : CascadeBuf
    port map (
            O => \N__10709\,
            I => \N__10706\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__1630\ : CascadeBuf
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__1628\ : CascadeBuf
    port map (
            O => \N__10697\,
            I => \N__10694\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__10694\,
            I => \N__10691\
        );

    \I__1626\ : InMux
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__10688\,
            I => \N__10685\
        );

    \I__1624\ : Span4Mux_v
    port map (
            O => \N__10685\,
            I => \N__10682\
        );

    \I__1623\ : Sp12to4
    port map (
            O => \N__10682\,
            I => \N__10679\
        );

    \I__1622\ : Span12Mux_h
    port map (
            O => \N__10679\,
            I => \N__10676\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__10676\,
            I => \M_this_vga_signals_address_0\
        );

    \I__1620\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10667\
        );

    \I__1619\ : InMux
    port map (
            O => \N__10672\,
            I => \N__10662\
        );

    \I__1618\ : InMux
    port map (
            O => \N__10671\,
            I => \N__10662\
        );

    \I__1617\ : InMux
    port map (
            O => \N__10670\,
            I => \N__10659\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__10667\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__10662\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__10659\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0\
        );

    \I__1613\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10644\
        );

    \I__1612\ : InMux
    port map (
            O => \N__10651\,
            I => \N__10641\
        );

    \I__1611\ : InMux
    port map (
            O => \N__10650\,
            I => \N__10634\
        );

    \I__1610\ : InMux
    port map (
            O => \N__10649\,
            I => \N__10634\
        );

    \I__1609\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10634\
        );

    \I__1608\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10631\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__10644\,
            I => \this_vga_signals.mult1_un82_sum_axb2_i\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__10641\,
            I => \this_vga_signals.mult1_un82_sum_axb2_i\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__10634\,
            I => \this_vga_signals.mult1_un82_sum_axb2_i\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__10631\,
            I => \this_vga_signals.mult1_un82_sum_axb2_i\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__10622\,
            I => \N__10619\
        );

    \I__1602\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10616\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__10616\,
            I => \N__10613\
        );

    \I__1600\ : Span4Mux_h
    port map (
            O => \N__10613\,
            I => \N__10606\
        );

    \I__1599\ : InMux
    port map (
            O => \N__10612\,
            I => \N__10603\
        );

    \I__1598\ : InMux
    port map (
            O => \N__10611\,
            I => \N__10600\
        );

    \I__1597\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10595\
        );

    \I__1596\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10595\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__10606\,
            I => \this_vga_signals.mult1_un82_sum_ac0_1\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__10603\,
            I => \this_vga_signals.mult1_un82_sum_ac0_1\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__10600\,
            I => \this_vga_signals.mult1_un82_sum_ac0_1\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__10595\,
            I => \this_vga_signals.mult1_un82_sum_ac0_1\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__10586\,
            I => \N__10581\
        );

    \I__1590\ : InMux
    port map (
            O => \N__10585\,
            I => \N__10577\
        );

    \I__1589\ : InMux
    port map (
            O => \N__10584\,
            I => \N__10572\
        );

    \I__1588\ : InMux
    port map (
            O => \N__10581\,
            I => \N__10572\
        );

    \I__1587\ : InMux
    port map (
            O => \N__10580\,
            I => \N__10569\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__10577\,
            I => \this_vga_signals.mult1_un82_sum_ac0_3_0_0\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__10572\,
            I => \this_vga_signals.mult1_un82_sum_ac0_3_0_0\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__10569\,
            I => \this_vga_signals.mult1_un82_sum_ac0_3_0_0\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__10562\,
            I => \N__10559\
        );

    \I__1582\ : CascadeBuf
    port map (
            O => \N__10559\,
            I => \N__10556\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__10556\,
            I => \N__10553\
        );

    \I__1580\ : CascadeBuf
    port map (
            O => \N__10553\,
            I => \N__10550\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__10550\,
            I => \N__10547\
        );

    \I__1578\ : CascadeBuf
    port map (
            O => \N__10547\,
            I => \N__10544\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__1576\ : CascadeBuf
    port map (
            O => \N__10541\,
            I => \N__10538\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__10538\,
            I => \N__10535\
        );

    \I__1574\ : CascadeBuf
    port map (
            O => \N__10535\,
            I => \N__10532\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__10532\,
            I => \N__10529\
        );

    \I__1572\ : CascadeBuf
    port map (
            O => \N__10529\,
            I => \N__10526\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__10526\,
            I => \N__10523\
        );

    \I__1570\ : CascadeBuf
    port map (
            O => \N__10523\,
            I => \N__10520\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__10520\,
            I => \N__10517\
        );

    \I__1568\ : CascadeBuf
    port map (
            O => \N__10517\,
            I => \N__10514\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__10514\,
            I => \N__10511\
        );

    \I__1566\ : CascadeBuf
    port map (
            O => \N__10511\,
            I => \N__10508\
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__10508\,
            I => \N__10505\
        );

    \I__1564\ : CascadeBuf
    port map (
            O => \N__10505\,
            I => \N__10502\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__10502\,
            I => \N__10499\
        );

    \I__1562\ : CascadeBuf
    port map (
            O => \N__10499\,
            I => \N__10496\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__10496\,
            I => \N__10493\
        );

    \I__1560\ : CascadeBuf
    port map (
            O => \N__10493\,
            I => \N__10490\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__10490\,
            I => \N__10487\
        );

    \I__1558\ : CascadeBuf
    port map (
            O => \N__10487\,
            I => \N__10484\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__10484\,
            I => \N__10481\
        );

    \I__1556\ : CascadeBuf
    port map (
            O => \N__10481\,
            I => \N__10478\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__10478\,
            I => \N__10475\
        );

    \I__1554\ : CascadeBuf
    port map (
            O => \N__10475\,
            I => \N__10472\
        );

    \I__1553\ : CascadeMux
    port map (
            O => \N__10472\,
            I => \N__10469\
        );

    \I__1552\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10466\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__10466\,
            I => \N__10463\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__10463\,
            I => \N__10460\
        );

    \I__1549\ : Span4Mux_v
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__1548\ : Sp12to4
    port map (
            O => \N__10457\,
            I => \N__10454\
        );

    \I__1547\ : Span12Mux_h
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__1546\ : Odrv12
    port map (
            O => \N__10451\,
            I => \M_this_vga_signals_address_1\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__10448\,
            I => \N__10441\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10447\,
            I => \N__10436\
        );

    \I__1543\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10433\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10428\
        );

    \I__1541\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10428\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10441\,
            I => \N__10421\
        );

    \I__1539\ : InMux
    port map (
            O => \N__10440\,
            I => \N__10421\
        );

    \I__1538\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10421\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__10436\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_i\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__10433\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_i\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__10428\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_i\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__10421\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_i\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10407\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__10411\,
            I => \N__10404\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__10410\,
            I => \N__10401\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__10407\,
            I => \N__10393\
        );

    \I__1529\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10386\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10401\,
            I => \N__10386\
        );

    \I__1527\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10386\
        );

    \I__1526\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10377\
        );

    \I__1525\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10377\
        );

    \I__1524\ : InMux
    port map (
            O => \N__10397\,
            I => \N__10377\
        );

    \I__1523\ : InMux
    port map (
            O => \N__10396\,
            I => \N__10377\
        );

    \I__1522\ : Odrv4
    port map (
            O => \N__10393\,
            I => \this_vga_signals.mult1_un75_sum_c3\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__10386\,
            I => \this_vga_signals.mult1_un75_sum_c3\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__10377\,
            I => \this_vga_signals.mult1_un75_sum_c3\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__1518\ : CascadeBuf
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__1516\ : CascadeBuf
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__1514\ : CascadeBuf
    port map (
            O => \N__10355\,
            I => \N__10352\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__1512\ : CascadeBuf
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__10346\,
            I => \N__10343\
        );

    \I__1510\ : CascadeBuf
    port map (
            O => \N__10343\,
            I => \N__10340\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__1508\ : CascadeBuf
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__1506\ : CascadeBuf
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__1504\ : CascadeBuf
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__10322\,
            I => \N__10319\
        );

    \I__1502\ : CascadeBuf
    port map (
            O => \N__10319\,
            I => \N__10316\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__10316\,
            I => \N__10313\
        );

    \I__1500\ : CascadeBuf
    port map (
            O => \N__10313\,
            I => \N__10310\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__10310\,
            I => \N__10307\
        );

    \I__1498\ : CascadeBuf
    port map (
            O => \N__10307\,
            I => \N__10304\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__10304\,
            I => \N__10301\
        );

    \I__1496\ : CascadeBuf
    port map (
            O => \N__10301\,
            I => \N__10298\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__10298\,
            I => \N__10295\
        );

    \I__1494\ : CascadeBuf
    port map (
            O => \N__10295\,
            I => \N__10292\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__10292\,
            I => \N__10289\
        );

    \I__1492\ : CascadeBuf
    port map (
            O => \N__10289\,
            I => \N__10286\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__10286\,
            I => \N__10283\
        );

    \I__1490\ : CascadeBuf
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__1488\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10274\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__10274\,
            I => \N__10271\
        );

    \I__1486\ : Span4Mux_h
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__1485\ : Sp12to4
    port map (
            O => \N__10268\,
            I => \N__10265\
        );

    \I__1484\ : Span12Mux_s9_v
    port map (
            O => \N__10265\,
            I => \N__10262\
        );

    \I__1483\ : Odrv12
    port map (
            O => \N__10262\,
            I => \M_this_vga_signals_address_2\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10256\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__10256\,
            I => \N__10252\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__10255\,
            I => \N__10247\
        );

    \I__1479\ : Span4Mux_v
    port map (
            O => \N__10252\,
            I => \N__10243\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10251\,
            I => \N__10240\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10237\
        );

    \I__1476\ : InMux
    port map (
            O => \N__10247\,
            I => \N__10232\
        );

    \I__1475\ : InMux
    port map (
            O => \N__10246\,
            I => \N__10232\
        );

    \I__1474\ : Odrv4
    port map (
            O => \N__10243\,
            I => \this_vga_signals.mult1_un61_sum_ac0_1\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__10240\,
            I => \this_vga_signals.mult1_un61_sum_ac0_1\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10237\,
            I => \this_vga_signals.mult1_un61_sum_ac0_1\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__10232\,
            I => \this_vga_signals.mult1_un61_sum_ac0_1\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10223\,
            I => \N__10216\
        );

    \I__1469\ : InMux
    port map (
            O => \N__10222\,
            I => \N__10212\
        );

    \I__1468\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10209\
        );

    \I__1467\ : InMux
    port map (
            O => \N__10220\,
            I => \N__10203\
        );

    \I__1466\ : InMux
    port map (
            O => \N__10219\,
            I => \N__10203\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10216\,
            I => \N__10196\
        );

    \I__1464\ : InMux
    port map (
            O => \N__10215\,
            I => \N__10193\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__10212\,
            I => \N__10190\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__10209\,
            I => \N__10187\
        );

    \I__1461\ : InMux
    port map (
            O => \N__10208\,
            I => \N__10184\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__10203\,
            I => \N__10181\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10178\
        );

    \I__1458\ : InMux
    port map (
            O => \N__10201\,
            I => \N__10175\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__10200\,
            I => \N__10172\
        );

    \I__1456\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10165\
        );

    \I__1455\ : Span4Mux_v
    port map (
            O => \N__10196\,
            I => \N__10154\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__10193\,
            I => \N__10154\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__10190\,
            I => \N__10141\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__10187\,
            I => \N__10141\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__10184\,
            I => \N__10141\
        );

    \I__1450\ : Span4Mux_h
    port map (
            O => \N__10181\,
            I => \N__10141\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__10178\,
            I => \N__10141\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__10175\,
            I => \N__10141\
        );

    \I__1447\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10136\
        );

    \I__1446\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10136\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10129\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10129\
        );

    \I__1443\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10129\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__10165\,
            I => \N__10126\
        );

    \I__1441\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10123\
        );

    \I__1440\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10120\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10111\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10111\
        );

    \I__1437\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10111\
        );

    \I__1436\ : InMux
    port map (
            O => \N__10159\,
            I => \N__10111\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__10154\,
            I => \this_vga_signals.mult1_un54_sum_i_0_3\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__10141\,
            I => \this_vga_signals.mult1_un54_sum_i_0_3\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__10136\,
            I => \this_vga_signals.mult1_un54_sum_i_0_3\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__10129\,
            I => \this_vga_signals.mult1_un54_sum_i_0_3\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__10126\,
            I => \this_vga_signals.mult1_un54_sum_i_0_3\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__10123\,
            I => \this_vga_signals.mult1_un54_sum_i_0_3\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__10120\,
            I => \this_vga_signals.mult1_un54_sum_i_0_3\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__10111\,
            I => \this_vga_signals.mult1_un54_sum_i_0_3\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__10094\,
            I => \N__10090\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10087\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10090\,
            I => \N__10083\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__10087\,
            I => \N__10080\
        );

    \I__1423\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10077\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__10083\,
            I => \N__10074\
        );

    \I__1421\ : Span4Mux_v
    port map (
            O => \N__10080\,
            I => \N__10071\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10077\,
            I => \N__10068\
        );

    \I__1419\ : Odrv12
    port map (
            O => \N__10074\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c\
        );

    \I__1418\ : Odrv4
    port map (
            O => \N__10071\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c\
        );

    \I__1417\ : Odrv4
    port map (
            O => \N__10068\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10057\
        );

    \I__1415\ : InMux
    port map (
            O => \N__10060\,
            I => \N__10046\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__10057\,
            I => \N__10043\
        );

    \I__1413\ : InMux
    port map (
            O => \N__10056\,
            I => \N__10034\
        );

    \I__1412\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10034\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10054\,
            I => \N__10034\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10053\,
            I => \N__10034\
        );

    \I__1409\ : InMux
    port map (
            O => \N__10052\,
            I => \N__10029\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__10051\,
            I => \N__10023\
        );

    \I__1407\ : InMux
    port map (
            O => \N__10050\,
            I => \N__10020\
        );

    \I__1406\ : InMux
    port map (
            O => \N__10049\,
            I => \N__10017\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__10046\,
            I => \N__10014\
        );

    \I__1404\ : Span4Mux_v
    port map (
            O => \N__10043\,
            I => \N__10009\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__10034\,
            I => \N__10009\
        );

    \I__1402\ : InMux
    port map (
            O => \N__10033\,
            I => \N__10004\
        );

    \I__1401\ : InMux
    port map (
            O => \N__10032\,
            I => \N__10004\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__10029\,
            I => \N__10001\
        );

    \I__1399\ : InMux
    port map (
            O => \N__10028\,
            I => \N__9996\
        );

    \I__1398\ : InMux
    port map (
            O => \N__10027\,
            I => \N__9996\
        );

    \I__1397\ : InMux
    port map (
            O => \N__10026\,
            I => \N__9991\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10023\,
            I => \N__9991\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__10020\,
            I => \this_vga_signals.mult1_un54_sum_m_ns_1\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__10017\,
            I => \this_vga_signals.mult1_un54_sum_m_ns_1\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__10014\,
            I => \this_vga_signals.mult1_un54_sum_m_ns_1\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__10009\,
            I => \this_vga_signals.mult1_un54_sum_m_ns_1\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__10004\,
            I => \this_vga_signals.mult1_un54_sum_m_ns_1\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__10001\,
            I => \this_vga_signals.mult1_un54_sum_m_ns_1\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__9996\,
            I => \this_vga_signals.mult1_un54_sum_m_ns_1\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__9991\,
            I => \this_vga_signals.mult1_un54_sum_m_ns_1\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__1386\ : CascadeBuf
    port map (
            O => \N__9971\,
            I => \N__9968\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__9968\,
            I => \N__9965\
        );

    \I__1384\ : CascadeBuf
    port map (
            O => \N__9965\,
            I => \N__9962\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__9962\,
            I => \N__9959\
        );

    \I__1382\ : CascadeBuf
    port map (
            O => \N__9959\,
            I => \N__9956\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__1380\ : CascadeBuf
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__9950\,
            I => \N__9947\
        );

    \I__1378\ : CascadeBuf
    port map (
            O => \N__9947\,
            I => \N__9944\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__1376\ : CascadeBuf
    port map (
            O => \N__9941\,
            I => \N__9938\
        );

    \I__1375\ : CascadeMux
    port map (
            O => \N__9938\,
            I => \N__9935\
        );

    \I__1374\ : CascadeBuf
    port map (
            O => \N__9935\,
            I => \N__9932\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__9932\,
            I => \N__9929\
        );

    \I__1372\ : CascadeBuf
    port map (
            O => \N__9929\,
            I => \N__9926\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__9926\,
            I => \N__9923\
        );

    \I__1370\ : CascadeBuf
    port map (
            O => \N__9923\,
            I => \N__9920\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__1368\ : CascadeBuf
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__9914\,
            I => \N__9911\
        );

    \I__1366\ : CascadeBuf
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__1364\ : CascadeBuf
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__1362\ : CascadeBuf
    port map (
            O => \N__9899\,
            I => \N__9896\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__9896\,
            I => \N__9893\
        );

    \I__1360\ : CascadeBuf
    port map (
            O => \N__9893\,
            I => \N__9890\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__9890\,
            I => \N__9887\
        );

    \I__1358\ : CascadeBuf
    port map (
            O => \N__9887\,
            I => \N__9884\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__9884\,
            I => \N__9881\
        );

    \I__1356\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9878\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__9878\,
            I => \N__9875\
        );

    \I__1354\ : Span4Mux_v
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__1353\ : Span4Mux_h
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__1352\ : Sp12to4
    port map (
            O => \N__9869\,
            I => \N__9866\
        );

    \I__1351\ : Span12Mux_h
    port map (
            O => \N__9866\,
            I => \N__9863\
        );

    \I__1350\ : Odrv12
    port map (
            O => \N__9863\,
            I => \M_this_vga_signals_address_4\
        );

    \I__1349\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9855\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__9859\,
            I => \N__9851\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__9858\,
            I => \N__9847\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__9855\,
            I => \N__9844\
        );

    \I__1345\ : InMux
    port map (
            O => \N__9854\,
            I => \N__9841\
        );

    \I__1344\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9834\
        );

    \I__1343\ : InMux
    port map (
            O => \N__9850\,
            I => \N__9834\
        );

    \I__1342\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9831\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__9844\,
            I => \N__9826\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__9841\,
            I => \N__9826\
        );

    \I__1339\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9821\
        );

    \I__1338\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9821\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__9834\,
            I => \N__9816\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__9831\,
            I => \N__9816\
        );

    \I__1335\ : Span4Mux_h
    port map (
            O => \N__9826\,
            I => \N__9813\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__9821\,
            I => \this_vga_signals.new_pixel_1\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__9816\,
            I => \this_vga_signals.new_pixel_1\
        );

    \I__1332\ : Odrv4
    port map (
            O => \N__9813\,
            I => \this_vga_signals.new_pixel_1\
        );

    \I__1331\ : InMux
    port map (
            O => \N__9806\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__1330\ : InMux
    port map (
            O => \N__9803\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__1329\ : InMux
    port map (
            O => \N__9800\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__9797\,
            I => \N__9787\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__9796\,
            I => \N__9782\
        );

    \I__1326\ : InMux
    port map (
            O => \N__9795\,
            I => \N__9774\
        );

    \I__1325\ : InMux
    port map (
            O => \N__9794\,
            I => \N__9774\
        );

    \I__1324\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9769\
        );

    \I__1323\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9769\
        );

    \I__1322\ : InMux
    port map (
            O => \N__9791\,
            I => \N__9764\
        );

    \I__1321\ : InMux
    port map (
            O => \N__9790\,
            I => \N__9764\
        );

    \I__1320\ : InMux
    port map (
            O => \N__9787\,
            I => \N__9757\
        );

    \I__1319\ : InMux
    port map (
            O => \N__9786\,
            I => \N__9757\
        );

    \I__1318\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9757\
        );

    \I__1317\ : InMux
    port map (
            O => \N__9782\,
            I => \N__9752\
        );

    \I__1316\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9752\
        );

    \I__1315\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9749\
        );

    \I__1314\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9746\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__9774\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__9769\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__9764\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__9757\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__9752\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__9749\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__9746\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1306\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9725\
        );

    \I__1305\ : InMux
    port map (
            O => \N__9730\,
            I => \N__9725\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__9725\,
            I => \this_vga_signals.N_19\
        );

    \I__1303\ : InMux
    port map (
            O => \N__9722\,
            I => \N__9718\
        );

    \I__1302\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9715\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__9718\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_0_1\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__9715\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_0_1\
        );

    \I__1299\ : CascadeMux
    port map (
            O => \N__9710\,
            I => \this_vga_signals.mult1_un75_sum_axb2_i_0_cascade_\
        );

    \I__1298\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9701\
        );

    \I__1297\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9701\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__9701\,
            I => \this_vga_signals.mult1_un75_sum_ac0_1_0\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__9698\,
            I => \this_vga_signals.g0_i_x2_0_0_a2_3_cascade_\
        );

    \I__1294\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9689\
        );

    \I__1293\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9689\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__9689\,
            I => \this_vga_signals.mult1_un75_sum_c3_0_0\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__9686\,
            I => \this_vga_signals.if_i4_mux_0_cascade_\
        );

    \I__1290\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9680\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__9680\,
            I => \this_vga_signals.g1_0_a2\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__9677\,
            I => \N__9674\
        );

    \I__1287\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9671\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__9671\,
            I => \this_vga_signals.g0_i_x2_0_0_a2_0\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__1284\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9662\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__9662\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0\
        );

    \I__1282\ : InMux
    port map (
            O => \N__9659\,
            I => \N__9656\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__9656\,
            I => \N__9652\
        );

    \I__1280\ : InMux
    port map (
            O => \N__9655\,
            I => \N__9649\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__9652\,
            I => \this_vga_signals.g1_1\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__9649\,
            I => \this_vga_signals.g1_1\
        );

    \I__1277\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__9641\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__9638\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0_cascade_\
        );

    \I__1274\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9628\
        );

    \I__1273\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9628\
        );

    \I__1272\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9625\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__9628\,
            I => \this_vga_signals.mult1_un68_sum_0_3\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__9625\,
            I => \this_vga_signals.mult1_un68_sum_0_3\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__9617\,
            I => \this_vga_signals.g0_0_a2_4\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9614\,
            I => \N__9608\
        );

    \I__1266\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9608\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__9608\,
            I => \N__9604\
        );

    \I__1264\ : InMux
    port map (
            O => \N__9607\,
            I => \N__9601\
        );

    \I__1263\ : Span4Mux_h
    port map (
            O => \N__9604\,
            I => \N__9598\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__9601\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_0\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__9598\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_0\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__9593\,
            I => \N__9590\
        );

    \I__1259\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9583\
        );

    \I__1258\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9583\
        );

    \I__1257\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9578\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__9583\,
            I => \N__9575\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9582\,
            I => \N__9570\
        );

    \I__1254\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9570\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__9578\,
            I => \this_vga_signals.mult1_un89_sum_c3\
        );

    \I__1252\ : Odrv12
    port map (
            O => \N__9575\,
            I => \this_vga_signals.mult1_un89_sum_c3\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__9570\,
            I => \this_vga_signals.mult1_un89_sum_c3\
        );

    \I__1250\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9560\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__9560\,
            I => \N__9555\
        );

    \I__1248\ : InMux
    port map (
            O => \N__9559\,
            I => \N__9550\
        );

    \I__1247\ : InMux
    port map (
            O => \N__9558\,
            I => \N__9550\
        );

    \I__1246\ : Span4Mux_v
    port map (
            O => \N__9555\,
            I => \N__9544\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__9550\,
            I => \N__9544\
        );

    \I__1244\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9541\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__9544\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__9541\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9533\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__9533\,
            I => \N__9530\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__9530\,
            I => \N__9527\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__9527\,
            I => \this_vga_signals.mult1_un75_sum_ac0_1_1\
        );

    \I__1237\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9521\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__9521\,
            I => \this_vga_signals.g0_13_N_4L5\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__9518\,
            I => \this_vga_signals.mult1_un75_sum_ac0_1_1_cascade_\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9515\,
            I => \N__9512\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__9512\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_3\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9503\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9500\
        );

    \I__1230\ : InMux
    port map (
            O => \N__9507\,
            I => \N__9495\
        );

    \I__1229\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9495\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__9503\,
            I => \this_vga_signals.mult1_un68_sum_1_3\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__9500\,
            I => \this_vga_signals.mult1_un68_sum_1_3\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__9495\,
            I => \this_vga_signals.mult1_un68_sum_1_3\
        );

    \I__1225\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9485\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__9485\,
            I => \this_vga_signals.mult1_un75_sum_axb2_i_1_0_0\
        );

    \I__1223\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9479\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__9479\,
            I => \this_vga_signals.g4\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__9476\,
            I => \this_vga_signals.g0_0_2_cascade_\
        );

    \I__1220\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9470\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__9470\,
            I => \this_vga_signals.g1_1_1_0_0\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__9467\,
            I => \N__9463\
        );

    \I__1217\ : InMux
    port map (
            O => \N__9466\,
            I => \N__9458\
        );

    \I__1216\ : InMux
    port map (
            O => \N__9463\,
            I => \N__9458\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__9455\,
            I => \this_vga_signals.N_4_0_0\
        );

    \I__1213\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__9446\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__9443\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_cascade_\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__9440\,
            I => \this_vga_signals.mult1_un68_sum_0_3_cascade_\
        );

    \I__1208\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__9431\,
            I => \this_vga_signals.g1_0_a2_0\
        );

    \I__1205\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9425\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__9425\,
            I => \N__9421\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__9424\,
            I => \N__9418\
        );

    \I__1202\ : Span4Mux_h
    port map (
            O => \N__9421\,
            I => \N__9415\
        );

    \I__1201\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9412\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__9415\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_6\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__9412\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_6\
        );

    \I__1198\ : InMux
    port map (
            O => \N__9407\,
            I => \N__9404\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__9404\,
            I => \N__9401\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__9401\,
            I => \this_vga_signals.M_hcounter_q_fast_esr_RNI52HLZ0Z_9\
        );

    \I__1195\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9394\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__9397\,
            I => \N__9389\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__9394\,
            I => \N__9386\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9383\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9378\
        );

    \I__1190\ : InMux
    port map (
            O => \N__9389\,
            I => \N__9378\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__9386\,
            I => \this_vga_signals.m8_0_1_0\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__9383\,
            I => \this_vga_signals.m8_0_1_0\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9378\,
            I => \this_vga_signals.m8_0_1_0\
        );

    \I__1186\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9364\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9359\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9369\,
            I => \N__9359\
        );

    \I__1183\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9352\
        );

    \I__1182\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9352\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__9364\,
            I => \N__9347\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__9359\,
            I => \N__9347\
        );

    \I__1179\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9342\
        );

    \I__1178\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9342\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__9352\,
            I => \this_vga_signals.M_hcounter_q_8_repZ0Z1\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__9347\,
            I => \this_vga_signals.M_hcounter_q_8_repZ0Z1\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__9342\,
            I => \this_vga_signals.M_hcounter_q_8_repZ0Z1\
        );

    \I__1174\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9331\
        );

    \I__1173\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9328\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__9331\,
            I => \this_vga_signals.m8_0_3\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__9328\,
            I => \this_vga_signals.m8_0_3\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9320\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__9320\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__9317\,
            I => \N__9314\
        );

    \I__1167\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__9311\,
            I => \this_vga_signals.g1_1_0_0\
        );

    \I__1165\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9305\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__9305\,
            I => \N__9302\
        );

    \I__1163\ : Span4Mux_h
    port map (
            O => \N__9302\,
            I => \N__9299\
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__9299\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_2_0\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__9296\,
            I => \this_vga_signals.g1_0_0_cascade_\
        );

    \I__1160\ : InMux
    port map (
            O => \N__9293\,
            I => \N__9290\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__9290\,
            I => \this_vga_signals.g1_6_0\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__9284\,
            I => \this_vga_signals.g4_1\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__9278\,
            I => \N__9274\
        );

    \I__1154\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9268\
        );

    \I__1153\ : Span4Mux_v
    port map (
            O => \N__9274\,
            I => \N__9265\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9262\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9257\
        );

    \I__1150\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9257\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__9268\,
            I => \N__9254\
        );

    \I__1148\ : Odrv4
    port map (
            O => \N__9265\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__9262\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__9257\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__9254\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__1144\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9241\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9238\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9241\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_9\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__9238\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_9\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__9233\,
            I => \N__9228\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__9232\,
            I => \N__9225\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__9231\,
            I => \N__9219\
        );

    \I__1137\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9216\
        );

    \I__1136\ : InMux
    port map (
            O => \N__9225\,
            I => \N__9213\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9210\
        );

    \I__1134\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9207\
        );

    \I__1133\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9204\
        );

    \I__1132\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9201\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__9216\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_7\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__9213\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_7\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__9210\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_7\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__9207\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_7\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__9204\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_7\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__9201\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_7\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__9188\,
            I => \N__9182\
        );

    \I__1124\ : InMux
    port map (
            O => \N__9187\,
            I => \N__9176\
        );

    \I__1123\ : InMux
    port map (
            O => \N__9186\,
            I => \N__9171\
        );

    \I__1122\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9171\
        );

    \I__1121\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9168\
        );

    \I__1120\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9165\
        );

    \I__1119\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9162\
        );

    \I__1118\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9159\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__9176\,
            I => \this_vga_signals.M_hcounter_q_6_repZ0Z1\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__9171\,
            I => \this_vga_signals.M_hcounter_q_6_repZ0Z1\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__9168\,
            I => \this_vga_signals.M_hcounter_q_6_repZ0Z1\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__9165\,
            I => \this_vga_signals.M_hcounter_q_6_repZ0Z1\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__9162\,
            I => \this_vga_signals.M_hcounter_q_6_repZ0Z1\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__9159\,
            I => \this_vga_signals.M_hcounter_q_6_repZ0Z1\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__9146\,
            I => \N__9139\
        );

    \I__1110\ : InMux
    port map (
            O => \N__9145\,
            I => \N__9136\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9130\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9125\
        );

    \I__1107\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9125\
        );

    \I__1106\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9122\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__9136\,
            I => \N__9119\
        );

    \I__1104\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9114\
        );

    \I__1103\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9114\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9133\,
            I => \N__9111\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__9130\,
            I => \this_vga_signals.M_hcounter_q_9_repZ0Z1\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__9125\,
            I => \this_vga_signals.M_hcounter_q_9_repZ0Z1\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__9122\,
            I => \this_vga_signals.M_hcounter_q_9_repZ0Z1\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__9119\,
            I => \this_vga_signals.M_hcounter_q_9_repZ0Z1\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__9114\,
            I => \this_vga_signals.M_hcounter_q_9_repZ0Z1\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__9111\,
            I => \this_vga_signals.M_hcounter_q_9_repZ0Z1\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__9098\,
            I => \this_vga_signals.M_hcounter_q_fast_esr_RNIHH441Z0Z_5_cascade_\
        );

    \I__1094\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9092\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__9092\,
            I => \this_vga_signals.M_hcounter_q_fast_esr_RNIN6RRZ0Z_7\
        );

    \I__1092\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__9086\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_5\
        );

    \I__1090\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__9080\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_8\
        );

    \I__1088\ : CEMux
    port map (
            O => \N__9077\,
            I => \N__9073\
        );

    \I__1087\ : CEMux
    port map (
            O => \N__9076\,
            I => \N__9070\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__9073\,
            I => \N__9063\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__9070\,
            I => \N__9063\
        );

    \I__1084\ : CEMux
    port map (
            O => \N__9069\,
            I => \N__9059\
        );

    \I__1083\ : CEMux
    port map (
            O => \N__9068\,
            I => \N__9055\
        );

    \I__1082\ : Span4Mux_v
    port map (
            O => \N__9063\,
            I => \N__9051\
        );

    \I__1081\ : CEMux
    port map (
            O => \N__9062\,
            I => \N__9048\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__9059\,
            I => \N__9045\
        );

    \I__1079\ : CEMux
    port map (
            O => \N__9058\,
            I => \N__9042\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__9055\,
            I => \N__9039\
        );

    \I__1077\ : CEMux
    port map (
            O => \N__9054\,
            I => \N__9036\
        );

    \I__1076\ : Span4Mux_h
    port map (
            O => \N__9051\,
            I => \N__9033\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__9048\,
            I => \N__9030\
        );

    \I__1074\ : Span4Mux_v
    port map (
            O => \N__9045\,
            I => \N__9023\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9042\,
            I => \N__9023\
        );

    \I__1072\ : Span4Mux_v
    port map (
            O => \N__9039\,
            I => \N__9023\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__9036\,
            I => \N__9020\
        );

    \I__1070\ : Odrv4
    port map (
            O => \N__9033\,
            I => \this_vga_signals.N_550_1\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__9030\,
            I => \this_vga_signals.N_550_1\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__9023\,
            I => \this_vga_signals.N_550_1\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__9020\,
            I => \this_vga_signals.N_550_1\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9011\,
            I => \N__9007\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9010\,
            I => \N__9002\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__9007\,
            I => \N__8999\
        );

    \I__1063\ : InMux
    port map (
            O => \N__9006\,
            I => \N__8996\
        );

    \I__1062\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8993\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__9002\,
            I => \this_vga_signals.m8_0_2\
        );

    \I__1060\ : Odrv4
    port map (
            O => \N__8999\,
            I => \this_vga_signals.m8_0_2\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__8996\,
            I => \this_vga_signals.m8_0_2\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__8993\,
            I => \this_vga_signals.m8_0_2\
        );

    \I__1057\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__8981\,
            I => \N__8978\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__8978\,
            I => \this_vga_signals.g1_0_1\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__8975\,
            I => \this_vga_signals.g4_1_1_cascade_\
        );

    \I__1053\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8967\
        );

    \I__1052\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8964\
        );

    \I__1051\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8961\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__8967\,
            I => \this_vga_signals.un1_haddress_0\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__8964\,
            I => \this_vga_signals.un1_haddress_0\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__8961\,
            I => \this_vga_signals.un1_haddress_0\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__8954\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_\
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__1045\ : InMux
    port map (
            O => \N__8948\,
            I => \N__8945\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__8945\,
            I => \this_vga_signals.un1_haddress_0_cry_1_c_RNOZ0\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__1042\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8935\
        );

    \I__1041\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8932\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__8935\,
            I => \N__8929\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__8932\,
            I => \this_vga_signals.m8_0_1_tz\
        );

    \I__1038\ : Odrv12
    port map (
            O => \N__8929\,
            I => \this_vga_signals.m8_0_1_tz\
        );

    \I__1037\ : InMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__8921\,
            I => \this_vga_signals.ANC2_4_1\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__8918\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__8915\,
            I => \N__8910\
        );

    \I__1033\ : InMux
    port map (
            O => \N__8914\,
            I => \N__8907\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__8913\,
            I => \N__8904\
        );

    \I__1031\ : InMux
    port map (
            O => \N__8910\,
            I => \N__8901\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__8907\,
            I => \N__8898\
        );

    \I__1029\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8895\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__8901\,
            I => \this_vga_signals.M_hcounter_q_7_repZ0Z1\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__8898\,
            I => \this_vga_signals.M_hcounter_q_7_repZ0Z1\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__8895\,
            I => \this_vga_signals.M_hcounter_q_7_repZ0Z1\
        );

    \I__1025\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8877\
        );

    \I__1024\ : InMux
    port map (
            O => \N__8887\,
            I => \N__8877\
        );

    \I__1023\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8872\
        );

    \I__1022\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8872\
        );

    \I__1021\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8867\
        );

    \I__1020\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8867\
        );

    \I__1019\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8864\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__8877\,
            I => \N__8861\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__8872\,
            I => \this_vga_signals.M_hcounter_q_5_repZ0Z1\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__8867\,
            I => \this_vga_signals.M_hcounter_q_5_repZ0Z1\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__8864\,
            I => \this_vga_signals.M_hcounter_q_5_repZ0Z1\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__8861\,
            I => \this_vga_signals.M_hcounter_q_5_repZ0Z1\
        );

    \I__1013\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8846\
        );

    \I__1012\ : InMux
    port map (
            O => \N__8851\,
            I => \N__8846\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__8846\,
            I => \this_vga_signals.mult1_un75_sum_axb1\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__8843\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_i_cascade_\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__8840\,
            I => \this_vga_signals.mult1_un82_sum_ac0_3_0_0_cascade_\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__8837\,
            I => \this_vga_signals.new_pixel_1_axb_1_N_4L5_xZ0Z1_cascade_\
        );

    \I__1007\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__8831\,
            I => \this_vga_signals.M_hcounter_q_RNIPIQRNRZ0Z_2\
        );

    \I__1005\ : InMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__8825\,
            I => \this_vga_signals.M_hcounter_q_RNI5HOBQCZ0Z_1\
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__8822\,
            I => \this_vga_signals.M_hcounter_q_RNI8TTVN32Z0Z_2_cascade_\
        );

    \I__1002\ : InMux
    port map (
            O => \N__8819\,
            I => \N__8816\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__8816\,
            I => \N__8813\
        );

    \I__1000\ : Span4Mux_h
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__8810\,
            I => \this_vga_signals.new_pixel_1_axb_1\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__8807\,
            I => \this_vga_signals.N_510_cascade_\
        );

    \I__997\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8801\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__8801\,
            I => \N__8797\
        );

    \I__995\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8794\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__8797\,
            I => \this_vga_signals.un1_haddress_0_axb_6\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__8794\,
            I => \this_vga_signals.un1_haddress_0_axb_6\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__8789\,
            I => \this_vga_signals.mult1_un75_sum_axb2_i_cascade_\
        );

    \I__991\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8781\
        );

    \I__990\ : InMux
    port map (
            O => \N__8785\,
            I => \N__8778\
        );

    \I__989\ : InMux
    port map (
            O => \N__8784\,
            I => \N__8771\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__8781\,
            I => \N__8766\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__8778\,
            I => \N__8766\
        );

    \I__986\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8763\
        );

    \I__985\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8758\
        );

    \I__984\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8758\
        );

    \I__983\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8755\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__8771\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__8766\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__8763\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__8758\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__8755\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__977\ : InMux
    port map (
            O => \N__8744\,
            I => \N__8741\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__8741\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_0_1_x1\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__8738\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_0_1_x0_cascade_\
        );

    \I__974\ : InMux
    port map (
            O => \N__8735\,
            I => \N__8729\
        );

    \I__973\ : InMux
    port map (
            O => \N__8734\,
            I => \N__8729\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__8729\,
            I => \this_vga_signals.mult1_un75_sum_ac0_1\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__8726\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_0_1_cascade_\
        );

    \I__970\ : InMux
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__8720\,
            I => \this_vga_signals.mult1_un75_sum_axb2_i\
        );

    \I__968\ : InMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__8714\,
            I => \this_vga_signals.mult1_un75_sum_axbxc2\
        );

    \I__966\ : InMux
    port map (
            O => \N__8711\,
            I => \N__8705\
        );

    \I__965\ : InMux
    port map (
            O => \N__8710\,
            I => \N__8700\
        );

    \I__964\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8700\
        );

    \I__963\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8697\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__8705\,
            I => \this_vga_signals.N_510_i\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__8700\,
            I => \this_vga_signals.N_510_i\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__8697\,
            I => \this_vga_signals.N_510_i\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__958\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8681\
        );

    \I__957\ : InMux
    port map (
            O => \N__8686\,
            I => \N__8681\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__8681\,
            I => \N__8673\
        );

    \I__955\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8670\
        );

    \I__954\ : InMux
    port map (
            O => \N__8679\,
            I => \N__8665\
        );

    \I__953\ : InMux
    port map (
            O => \N__8678\,
            I => \N__8665\
        );

    \I__952\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8659\
        );

    \I__951\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8656\
        );

    \I__950\ : Span4Mux_v
    port map (
            O => \N__8673\,
            I => \N__8649\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__8670\,
            I => \N__8649\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__8665\,
            I => \N__8649\
        );

    \I__947\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8642\
        );

    \I__946\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8642\
        );

    \I__945\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8642\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__8659\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__8656\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__8649\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__8642\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__8633\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_cascade_\
        );

    \I__939\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8627\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__8627\,
            I => \this_vga_signals.mult1_un75_sum_axb2_0_0\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__8624\,
            I => \this_vga_signals.mult1_un75_sum_axb2_0_0_cascade_\
        );

    \I__936\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8615\
        );

    \I__935\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8610\
        );

    \I__934\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8610\
        );

    \I__933\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8607\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__8615\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__8610\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__8607\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__8600\,
            I => \N__8595\
        );

    \I__928\ : InMux
    port map (
            O => \N__8599\,
            I => \N__8588\
        );

    \I__927\ : InMux
    port map (
            O => \N__8598\,
            I => \N__8588\
        );

    \I__926\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8581\
        );

    \I__925\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8581\
        );

    \I__924\ : InMux
    port map (
            O => \N__8593\,
            I => \N__8581\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__8588\,
            I => \this_vga_signals.if_m2_0\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__8581\,
            I => \this_vga_signals.if_m2_0\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__8576\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5_cascade_\
        );

    \I__920\ : InMux
    port map (
            O => \N__8573\,
            I => \N__8570\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__8570\,
            I => \this_vga_signals.g0_10_3_0_a2_0_0\
        );

    \I__918\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__8564\,
            I => \N__8561\
        );

    \I__916\ : Span4Mux_v
    port map (
            O => \N__8561\,
            I => \N__8558\
        );

    \I__915\ : Odrv4
    port map (
            O => \N__8558\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_1\
        );

    \I__914\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8551\
        );

    \I__913\ : InMux
    port map (
            O => \N__8554\,
            I => \N__8548\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__8551\,
            I => \N__8545\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__8548\,
            I => \this_vga_signals.g1_0\
        );

    \I__910\ : Odrv12
    port map (
            O => \N__8545\,
            I => \this_vga_signals.g1_0\
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__8540\,
            I => \this_vga_signals.g0_10_3_0_a2_0_0_cascade_\
        );

    \I__908\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__8534\,
            I => \this_vga_signals.mult1_un75_sum_axb2_x0\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__905\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8525\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__8525\,
            I => \this_vga_signals.mult1_un75_sum_axb2_x1\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__8522\,
            I => \this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOMZ0Z71_cascade_\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__8519\,
            I => \this_vga_signals.m8_0_2_cascade_\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__8516\,
            I => \this_vga_signals.mult1_un61_sum_ac0_1_cascade_\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__8513\,
            I => \this_vga_signals.mult1_un54_sum_i_0_3_cascade_\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__8510\,
            I => \this_vga_signals.g1_6_0_cascade_\
        );

    \I__898\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__8504\,
            I => \N__8500\
        );

    \I__896\ : InMux
    port map (
            O => \N__8503\,
            I => \N__8497\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__8500\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__8497\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3\
        );

    \I__893\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__8489\,
            I => \this_vga_signals.g0_13_N_3L3_ns\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__8486\,
            I => \this_vga_signals.g0_13_N_2L1_cascade_\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__8483\,
            I => \this_vga_signals.N_75_cascade_\
        );

    \I__889\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__8477\,
            I => \this_vga_signals.mult1_un54_sum_m_1_1\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__8474\,
            I => \this_vga_signals.mult1_un54_sum_m_1_1_cascade_\
        );

    \I__886\ : InMux
    port map (
            O => \N__8471\,
            I => \N__8468\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__8468\,
            I => \this_vga_signals.N_75\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__8465\,
            I => \this_vga_signals.mult1_un54_sum_m_x0_1_cascade_\
        );

    \I__883\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8459\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__8459\,
            I => \this_vga_signals.mult1_un54_sum_m_x1_1\
        );

    \I__881\ : InMux
    port map (
            O => \N__8456\,
            I => \this_vga_signals.un1_haddress_0_cry_5\
        );

    \I__880\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8449\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__8452\,
            I => \N__8446\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__8449\,
            I => \N__8443\
        );

    \I__877\ : InMux
    port map (
            O => \N__8446\,
            I => \N__8440\
        );

    \I__876\ : Odrv12
    port map (
            O => \N__8443\,
            I => \this_vga_signals.un1_haddress_0_axb_7\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__8440\,
            I => \this_vga_signals.un1_haddress_0_axb_7\
        );

    \I__874\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8432\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__872\ : Span4Mux_h
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__871\ : Odrv4
    port map (
            O => \N__8426\,
            I => \this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQUZ0\
        );

    \I__870\ : InMux
    port map (
            O => \N__8423\,
            I => \this_vga_signals.un1_haddress_0_cry_6\
        );

    \I__869\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8416\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__8419\,
            I => \N__8413\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__8416\,
            I => \N__8410\
        );

    \I__866\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8407\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__8410\,
            I => \this_vga_signals.un1_haddress_0_cry_7_i\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__8407\,
            I => \this_vga_signals.un1_haddress_0_cry_7_i\
        );

    \I__863\ : InMux
    port map (
            O => \N__8402\,
            I => \this_vga_signals.un1_haddress_0_cry_7\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__861\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8393\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__859\ : Span4Mux_h
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__858\ : Odrv4
    port map (
            O => \N__8387\,
            I => \this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBSZ0Z7\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__8384\,
            I => \this_vga_signals.m8_0_1_tz_cascade_\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__8381\,
            I => \this_vga_signals.g1_cascade_\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__8378\,
            I => \this_vga_signals.g1_1_0_cascade_\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__8375\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9_cascade_\
        );

    \I__853\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8369\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8369\,
            I => \N__8366\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__8366\,
            I => \N__8363\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__8363\,
            I => \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TAZ0Z7\
        );

    \I__849\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8357\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__8357\,
            I => \this_vga_signals.mult1_un75_sum_i_0_3\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__8354\,
            I => \N__8351\
        );

    \I__846\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8348\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__8348\,
            I => \this_vga_signals.un1_haddress_0_axb_2_l_ofxZ0\
        );

    \I__844\ : InMux
    port map (
            O => \N__8345\,
            I => \N__8342\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__842\ : Span4Mux_h
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__841\ : Odrv4
    port map (
            O => \N__8336\,
            I => \this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44VZ0Z02\
        );

    \I__840\ : InMux
    port map (
            O => \N__8333\,
            I => \this_vga_signals.un1_haddress_0_cry_1\
        );

    \I__839\ : InMux
    port map (
            O => \N__8330\,
            I => \N__8327\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__8327\,
            I => \this_vga_signals.un1_haddress_0_axb_3_l_fxZ0\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__8324\,
            I => \N__8321\
        );

    \I__836\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8317\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__8320\,
            I => \N__8314\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__8317\,
            I => \N__8311\
        );

    \I__833\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8308\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__8311\,
            I => \this_vga_signals.mult1_un68_sum_i_3\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8308\,
            I => \this_vga_signals.mult1_un68_sum_i_3\
        );

    \I__830\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8300\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__8300\,
            I => \N__8297\
        );

    \I__828\ : Span4Mux_v
    port map (
            O => \N__8297\,
            I => \N__8294\
        );

    \I__827\ : Odrv4
    port map (
            O => \N__8294\,
            I => \this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9DZ0\
        );

    \I__826\ : InMux
    port map (
            O => \N__8291\,
            I => \this_vga_signals.un1_haddress_0_cry_2\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__8288\,
            I => \N__8285\
        );

    \I__824\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8282\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__8282\,
            I => \N__8279\
        );

    \I__822\ : Odrv12
    port map (
            O => \N__8279\,
            I => \this_vga_signals.un1_haddress_0_axb_4_l_fxZ0\
        );

    \I__821\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8273\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8270\
        );

    \I__819\ : Span4Mux_v
    port map (
            O => \N__8270\,
            I => \N__8267\
        );

    \I__818\ : Odrv4
    port map (
            O => \N__8267\,
            I => \this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4TZ0Z72\
        );

    \I__817\ : InMux
    port map (
            O => \N__8264\,
            I => \this_vga_signals.un1_haddress_0_cry_3\
        );

    \I__816\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8258\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__8258\,
            I => \N__8255\
        );

    \I__814\ : Span4Mux_h
    port map (
            O => \N__8255\,
            I => \N__8252\
        );

    \I__813\ : Odrv4
    port map (
            O => \N__8252\,
            I => \this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJLZ0\
        );

    \I__812\ : InMux
    port map (
            O => \N__8249\,
            I => \this_vga_signals.un1_haddress_0_cry_4\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__8246\,
            I => \N__8243\
        );

    \I__810\ : InMux
    port map (
            O => \N__8243\,
            I => \N__8240\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__8240\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9\
        );

    \I__808\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8231\
        );

    \I__807\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8231\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__8231\,
            I => \this_vga_signals.un1_haddress_0_cry_5_THRU_CO\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__8228\,
            I => \this_vga_signals.mult1_un75_sum_axb2_i_1_cascade_\
        );

    \I__804\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8222\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__8222\,
            I => \N__8219\
        );

    \I__802\ : Odrv12
    port map (
            O => \N__8219\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_1\
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__8216\,
            I => \this_vga_signals.N_4_i_1_cascade_\
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__8213\,
            I => \this_vga_signals.mult1_un82_sum_ac0_1_cascade_\
        );

    \I__799\ : InMux
    port map (
            O => \N__8210\,
            I => \N__8207\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__8207\,
            I => \this_vga_signals.N_4_i\
        );

    \I__797\ : CascadeMux
    port map (
            O => \N__8204\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_cascade_\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__8201\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_cascade_\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__794\ : CascadeBuf
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__8192\,
            I => \N__8189\
        );

    \I__792\ : CascadeBuf
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__8186\,
            I => \N__8183\
        );

    \I__790\ : CascadeBuf
    port map (
            O => \N__8183\,
            I => \N__8180\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__8180\,
            I => \N__8177\
        );

    \I__788\ : CascadeBuf
    port map (
            O => \N__8177\,
            I => \N__8174\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__8174\,
            I => \N__8171\
        );

    \I__786\ : CascadeBuf
    port map (
            O => \N__8171\,
            I => \N__8168\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__8168\,
            I => \N__8165\
        );

    \I__784\ : CascadeBuf
    port map (
            O => \N__8165\,
            I => \N__8162\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__8162\,
            I => \N__8159\
        );

    \I__782\ : CascadeBuf
    port map (
            O => \N__8159\,
            I => \N__8156\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__8156\,
            I => \N__8153\
        );

    \I__780\ : CascadeBuf
    port map (
            O => \N__8153\,
            I => \N__8150\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__8150\,
            I => \N__8147\
        );

    \I__778\ : CascadeBuf
    port map (
            O => \N__8147\,
            I => \N__8144\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__8144\,
            I => \N__8141\
        );

    \I__776\ : CascadeBuf
    port map (
            O => \N__8141\,
            I => \N__8138\
        );

    \I__775\ : CascadeMux
    port map (
            O => \N__8138\,
            I => \N__8135\
        );

    \I__774\ : CascadeBuf
    port map (
            O => \N__8135\,
            I => \N__8132\
        );

    \I__773\ : CascadeMux
    port map (
            O => \N__8132\,
            I => \N__8129\
        );

    \I__772\ : CascadeBuf
    port map (
            O => \N__8129\,
            I => \N__8126\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__8126\,
            I => \N__8123\
        );

    \I__770\ : CascadeBuf
    port map (
            O => \N__8123\,
            I => \N__8120\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__8120\,
            I => \N__8117\
        );

    \I__768\ : CascadeBuf
    port map (
            O => \N__8117\,
            I => \N__8114\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__8114\,
            I => \N__8111\
        );

    \I__766\ : CascadeBuf
    port map (
            O => \N__8111\,
            I => \N__8108\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__8108\,
            I => \N__8105\
        );

    \I__764\ : InMux
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__8102\,
            I => \N__8099\
        );

    \I__762\ : Span12Mux_s10_h
    port map (
            O => \N__8099\,
            I => \N__8096\
        );

    \I__761\ : Span12Mux_v
    port map (
            O => \N__8096\,
            I => \N__8093\
        );

    \I__760\ : Span12Mux_h
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__759\ : Odrv12
    port map (
            O => \N__8090\,
            I => \M_this_vga_signals_address_3\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__8087\,
            I => \this_vga_signals.M_hcounter_d6lt9_cascade_\
        );

    \I__757\ : InMux
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__755\ : Span4Mux_v
    port map (
            O => \N__8078\,
            I => \N__8073\
        );

    \I__754\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8068\
        );

    \I__753\ : InMux
    port map (
            O => \N__8076\,
            I => \N__8068\
        );

    \I__752\ : Span4Mux_h
    port map (
            O => \N__8073\,
            I => \N__8065\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8068\,
            I => \this_pixel_clock_M_counter_q_i_1\
        );

    \I__750\ : Odrv4
    port map (
            O => \N__8065\,
            I => \this_pixel_clock_M_counter_q_i_1\
        );

    \I__749\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8055\
        );

    \I__748\ : InMux
    port map (
            O => \N__8059\,
            I => \N__8049\
        );

    \I__747\ : InMux
    port map (
            O => \N__8058\,
            I => \N__8049\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__8055\,
            I => \N__8046\
        );

    \I__745\ : InMux
    port map (
            O => \N__8054\,
            I => \N__8043\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__8049\,
            I => \N__8040\
        );

    \I__743\ : Span4Mux_h
    port map (
            O => \N__8046\,
            I => \N__8037\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__8043\,
            I => \this_pixel_clock_M_counter_q_0\
        );

    \I__741\ : Odrv4
    port map (
            O => \N__8040\,
            I => \this_pixel_clock_M_counter_q_0\
        );

    \I__740\ : Odrv4
    port map (
            O => \N__8037\,
            I => \this_pixel_clock_M_counter_q_0\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__8030\,
            I => \this_vga_signals.M_hcounter_d6_0_cascade_\
        );

    \I__738\ : IoInMux
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__736\ : IoSpan4Mux
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__735\ : Span4Mux_s2_h
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__734\ : Sp12to4
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__733\ : Span12Mux_s5_h
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__732\ : Span12Mux_h
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__731\ : Odrv12
    port map (
            O => \N__8006\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIUKG82Z0Z_9\
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__8003\,
            I => \this_vga_signals.mult1_un75_sum_ac0_1_sx_cascade_\
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__8000\,
            I => \this_vga_signals.if_m2_0_cascade_\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__7997\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__7994\,
            I => \this_vga_signals.g0_13_N_3L3_x0_cascade_\
        );

    \I__726\ : InMux
    port map (
            O => \N__7991\,
            I => \N__7987\
        );

    \I__725\ : InMux
    port map (
            O => \N__7990\,
            I => \N__7984\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__7987\,
            I => \N__7981\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__7984\,
            I => \N__7978\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__7981\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_2_0_0\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__7978\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_2_0_0\
        );

    \I__720\ : InMux
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__7970\,
            I => \this_vga_signals.g0_13_N_3L3_x1\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__7967\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_\
        );

    \I__717\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7961\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__7961\,
            I => \this_vga_signals.M_hcounter_q_RNIUA42NDZ0Z_1\
        );

    \I__715\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7955\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__7955\,
            I => \this_vga_signals.new_pixel_1_cry_0_c_RNOZ0\
        );

    \I__713\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7949\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__7949\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIG53KZ0Z_9\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__7946\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1_cascade_\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__7943\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_1_cascade_\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__7940\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4_cascade_\
        );

    \I__708\ : IoInMux
    port map (
            O => \N__7937\,
            I => \N__7934\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__706\ : IoSpan4Mux
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__705\ : Span4Mux_s1_v
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__704\ : Span4Mux_v
    port map (
            O => \N__7925\,
            I => \N__7922\
        );

    \I__703\ : Odrv4
    port map (
            O => \N__7922\,
            I => debug_c_i_1
        );

    \I__702\ : CascadeMux
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__701\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__7913\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIG53K_1Z0Z_9\
        );

    \I__699\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__7907\,
            I => \this_vga_signals.un3_hsynclt8_0\
        );

    \I__697\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7901\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__7901\,
            I => \N__7898\
        );

    \I__695\ : Odrv4
    port map (
            O => \N__7898\,
            I => \this_vga_signals.new_pixel_1_i_0\
        );

    \I__694\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7892\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__7892\,
            I => \this_vga_signals.new_pixel_1_5\
        );

    \I__692\ : InMux
    port map (
            O => \N__7889\,
            I => \this_vga_signals.new_pixel_1_cry_4\
        );

    \I__691\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__7883\,
            I => \this_vga_signals.new_pixel_1_6\
        );

    \I__689\ : InMux
    port map (
            O => \N__7880\,
            I => \this_vga_signals.new_pixel_1_cry_5\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__687\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7871\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__7871\,
            I => \this_vga_signals.M_hcounter_q_i_7\
        );

    \I__685\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7865\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__7865\,
            I => \this_vga_signals.new_pixel_1_7\
        );

    \I__683\ : InMux
    port map (
            O => \N__7862\,
            I => \this_vga_signals.new_pixel_1_cry_6\
        );

    \I__682\ : InMux
    port map (
            O => \N__7859\,
            I => \N__7856\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__7856\,
            I => \this_vga_signals.new_pixel_1_8\
        );

    \I__680\ : InMux
    port map (
            O => \N__7853\,
            I => \bfn_6_22_0_\
        );

    \I__679\ : InMux
    port map (
            O => \N__7850\,
            I => \N__7847\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__7847\,
            I => \this_vga_signals.new_pixel_1_9\
        );

    \I__677\ : InMux
    port map (
            O => \N__7844\,
            I => \this_vga_signals.new_pixel_1_cry_8\
        );

    \I__676\ : InMux
    port map (
            O => \N__7841\,
            I => \N__7838\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__7838\,
            I => \this_vga_signals.new_pixel_1_10\
        );

    \I__674\ : InMux
    port map (
            O => \N__7835\,
            I => \this_vga_signals.new_pixel_1_cry_9\
        );

    \I__673\ : InMux
    port map (
            O => \N__7832\,
            I => \this_vga_signals.new_pixel_1_cry_10\
        );

    \I__672\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__7826\,
            I => \this_vga_signals.new_pixel_1_11\
        );

    \I__670\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__7820\,
            I => \N__7817\
        );

    \I__668\ : Odrv12
    port map (
            O => \N__7817\,
            I => \this_vga_signals.un4_hsynclt8_0\
        );

    \I__667\ : IoInMux
    port map (
            O => \N__7814\,
            I => \N__7811\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__7811\,
            I => \N__7808\
        );

    \I__665\ : Span4Mux_s3_v
    port map (
            O => \N__7808\,
            I => \N__7805\
        );

    \I__664\ : Span4Mux_h
    port map (
            O => \N__7805\,
            I => \N__7802\
        );

    \I__663\ : Span4Mux_v
    port map (
            O => \N__7802\,
            I => \N__7799\
        );

    \I__662\ : Odrv4
    port map (
            O => \N__7799\,
            I => this_vga_signals_hsync_1_i
        );

    \I__661\ : CascadeMux
    port map (
            O => \N__7796\,
            I => \N_50_cascade_\
        );

    \I__660\ : IoInMux
    port map (
            O => \N__7793\,
            I => \N__7790\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__7790\,
            I => \N__7787\
        );

    \I__658\ : Span4Mux_s0_v
    port map (
            O => \N__7787\,
            I => \N__7784\
        );

    \I__657\ : Sp12to4
    port map (
            O => \N__7784\,
            I => \N__7781\
        );

    \I__656\ : Span12Mux_h
    port map (
            O => \N__7781\,
            I => \N__7777\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__7780\,
            I => \N__7771\
        );

    \I__654\ : Span12Mux_v
    port map (
            O => \N__7777\,
            I => \N__7767\
        );

    \I__653\ : InMux
    port map (
            O => \N__7776\,
            I => \N__7764\
        );

    \I__652\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7759\
        );

    \I__651\ : InMux
    port map (
            O => \N__7774\,
            I => \N__7759\
        );

    \I__650\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7754\
        );

    \I__649\ : InMux
    port map (
            O => \N__7770\,
            I => \N__7754\
        );

    \I__648\ : Odrv12
    port map (
            O => \N__7767\,
            I => debug_c_0
        );

    \I__647\ : LocalMux
    port map (
            O => \N__7764\,
            I => debug_c_0
        );

    \I__646\ : LocalMux
    port map (
            O => \N__7759\,
            I => debug_c_0
        );

    \I__645\ : LocalMux
    port map (
            O => \N__7754\,
            I => debug_c_0
        );

    \I__644\ : IoInMux
    port map (
            O => \N__7745\,
            I => \N__7742\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__7742\,
            I => \N__7739\
        );

    \I__642\ : IoSpan4Mux
    port map (
            O => \N__7739\,
            I => \N__7735\
        );

    \I__641\ : InMux
    port map (
            O => \N__7738\,
            I => \N__7732\
        );

    \I__640\ : Span4Mux_s3_h
    port map (
            O => \N__7735\,
            I => \N__7727\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__7732\,
            I => \N__7727\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__7727\,
            I => rgb_c_2
        );

    \I__637\ : InMux
    port map (
            O => \N__7724\,
            I => \N__7716\
        );

    \I__636\ : InMux
    port map (
            O => \N__7723\,
            I => \N__7713\
        );

    \I__635\ : InMux
    port map (
            O => \N__7722\,
            I => \N__7708\
        );

    \I__634\ : InMux
    port map (
            O => \N__7721\,
            I => \N__7708\
        );

    \I__633\ : InMux
    port map (
            O => \N__7720\,
            I => \N__7703\
        );

    \I__632\ : InMux
    port map (
            O => \N__7719\,
            I => \N__7703\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__7716\,
            I => \M_hcounter_q_esr_RNIH8GJ4_9\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__7713\,
            I => \M_hcounter_q_esr_RNIH8GJ4_9\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__7708\,
            I => \M_hcounter_q_esr_RNIH8GJ4_9\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__7703\,
            I => \M_hcounter_q_esr_RNIH8GJ4_9\
        );

    \I__627\ : InMux
    port map (
            O => \N__7694\,
            I => \N__7691\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__7691\,
            I => \this_vga_signals.new_pixel_1Z0Z_1\
        );

    \I__625\ : InMux
    port map (
            O => \N__7688\,
            I => \this_vga_signals.new_pixel_1_cry_0\
        );

    \I__624\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7682\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__7682\,
            I => \this_vga_signals.new_pixel_1_2\
        );

    \I__622\ : InMux
    port map (
            O => \N__7679\,
            I => \this_vga_signals.new_pixel_1_cry_1\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__7676\,
            I => \N__7673\
        );

    \I__620\ : InMux
    port map (
            O => \N__7673\,
            I => \N__7670\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__7670\,
            I => \N__7667\
        );

    \I__618\ : Odrv4
    port map (
            O => \N__7667\,
            I => \this_vga_signals.new_pixel_1_3\
        );

    \I__617\ : InMux
    port map (
            O => \N__7664\,
            I => \this_vga_signals.new_pixel_1_cry_2\
        );

    \I__616\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7658\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__7658\,
            I => \this_vga_signals.new_pixel_1_4\
        );

    \I__614\ : InMux
    port map (
            O => \N__7655\,
            I => \this_vga_signals.new_pixel_1_cry_3\
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__7652\,
            I => \this_vga_signals.new_pixel_1_1_cascade_\
        );

    \I__612\ : CascadeMux
    port map (
            O => \N__7649\,
            I => \debug_c_0_cascade_\
        );

    \I__611\ : IoInMux
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__7643\,
            I => \N__7640\
        );

    \I__609\ : Span4Mux_s2_h
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__608\ : Span4Mux_v
    port map (
            O => \N__7637\,
            I => \N__7633\
        );

    \I__607\ : InMux
    port map (
            O => \N__7636\,
            I => \N__7630\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__7633\,
            I => rgb_c_3
        );

    \I__605\ : LocalMux
    port map (
            O => \N__7630\,
            I => rgb_c_3
        );

    \I__604\ : InMux
    port map (
            O => \N__7625\,
            I => \N__7622\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__7622\,
            I => \N__7619\
        );

    \I__602\ : Odrv4
    port map (
            O => \N__7619\,
            I => \N_37\
        );

    \I__601\ : IoInMux
    port map (
            O => \N__7616\,
            I => \N__7613\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__7613\,
            I => \N__7610\
        );

    \I__599\ : IoSpan4Mux
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__598\ : Span4Mux_s3_v
    port map (
            O => \N__7607\,
            I => \N__7604\
        );

    \I__597\ : Span4Mux_v
    port map (
            O => \N__7604\,
            I => \N__7600\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__7603\,
            I => \N__7597\
        );

    \I__595\ : Span4Mux_v
    port map (
            O => \N__7600\,
            I => \N__7594\
        );

    \I__594\ : InMux
    port map (
            O => \N__7597\,
            I => \N__7591\
        );

    \I__593\ : Odrv4
    port map (
            O => \N__7594\,
            I => rgb_c_4
        );

    \I__592\ : LocalMux
    port map (
            O => \N__7591\,
            I => rgb_c_4
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__7586\,
            I => \this_vga_signals.new_pixel_1_3_1_cascade_\
        );

    \I__590\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7580\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__7580\,
            I => \this_vga_signals.new_pixel_sx_0\
        );

    \I__588\ : IoInMux
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__586\ : Odrv12
    port map (
            O => \N__7571\,
            I => this_vga_signals_vvisibility_i
        );

    \I__585\ : InMux
    port map (
            O => \N__7568\,
            I => \N__7565\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__7565\,
            I => \N_60\
        );

    \I__583\ : InMux
    port map (
            O => \N__7562\,
            I => \N__7559\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__7559\,
            I => \N__7556\
        );

    \I__581\ : Odrv4
    port map (
            O => \N__7556\,
            I => i7_mux
        );

    \I__580\ : IoInMux
    port map (
            O => \N__7553\,
            I => \N__7550\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__7550\,
            I => \N__7547\
        );

    \I__578\ : Span12Mux_s3_h
    port map (
            O => \N__7547\,
            I => \N__7544\
        );

    \I__577\ : Odrv12
    port map (
            O => \N__7544\,
            I => port_nmib_0_i
        );

    \I__576\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7538\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__7538\,
            I => \N__7535\
        );

    \I__574\ : Odrv12
    port map (
            O => \N__7535\,
            I => port_clk_c
        );

    \I__573\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7529\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__7529\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__571\ : IoInMux
    port map (
            O => \N__7526\,
            I => \N__7523\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__7523\,
            I => \N__7520\
        );

    \I__569\ : Span4Mux_s0_h
    port map (
            O => \N__7520\,
            I => \N__7517\
        );

    \I__568\ : Span4Mux_h
    port map (
            O => \N__7517\,
            I => \N__7514\
        );

    \I__567\ : Sp12to4
    port map (
            O => \N__7514\,
            I => \N__7511\
        );

    \I__566\ : Span12Mux_v
    port map (
            O => \N__7511\,
            I => \N__7507\
        );

    \I__565\ : InMux
    port map (
            O => \N__7510\,
            I => \N__7504\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__7507\,
            I => rgb_c_0
        );

    \I__563\ : LocalMux
    port map (
            O => \N__7504\,
            I => rgb_c_0
        );

    \I__562\ : InMux
    port map (
            O => \N__7499\,
            I => \N__7496\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__7496\,
            I => i7_mux_0
        );

    \I__560\ : IoInMux
    port map (
            O => \N__7493\,
            I => \N__7490\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__558\ : IoSpan4Mux
    port map (
            O => \N__7487\,
            I => \N__7483\
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__7486\,
            I => \N__7480\
        );

    \I__556\ : Span4Mux_s2_h
    port map (
            O => \N__7483\,
            I => \N__7477\
        );

    \I__555\ : InMux
    port map (
            O => \N__7480\,
            I => \N__7474\
        );

    \I__554\ : Odrv4
    port map (
            O => \N__7477\,
            I => rgb_c_1
        );

    \I__553\ : LocalMux
    port map (
            O => \N__7474\,
            I => rgb_c_1
        );

    \I__552\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7466\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__7466\,
            I => \N__7463\
        );

    \I__550\ : Odrv4
    port map (
            O => \N__7463\,
            I => \N_28_0\
        );

    \I__549\ : IoInMux
    port map (
            O => \N__7460\,
            I => \N__7457\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__547\ : IoSpan4Mux
    port map (
            O => \N__7454\,
            I => \N__7450\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__7453\,
            I => \N__7447\
        );

    \I__545\ : IoSpan4Mux
    port map (
            O => \N__7450\,
            I => \N__7444\
        );

    \I__544\ : InMux
    port map (
            O => \N__7447\,
            I => \N__7441\
        );

    \I__543\ : Span4Mux_s3_h
    port map (
            O => \N__7444\,
            I => \N__7438\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__7441\,
            I => \N__7435\
        );

    \I__541\ : Odrv4
    port map (
            O => \N__7438\,
            I => rgb_c_5
        );

    \I__540\ : Odrv4
    port map (
            O => \N__7435\,
            I => rgb_c_5
        );

    \I__539\ : IoInMux
    port map (
            O => \N__7430\,
            I => \N__7427\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__7427\,
            I => \N_377_i\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_6_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_21_0_\
        );

    \IN_MUX_bfv_6_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.new_pixel_1_cry_7\,
            carryinitout => \bfn_6_22_0_\
        );

    \IN_MUX_bfv_30_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_30_23_0_\
        );

    \IN_MUX_bfv_30_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_external_address_q_cry_7\,
            carryinitout => \bfn_30_24_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_20_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_21_0_\
        );

    \IN_MUX_bfv_20_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_internal_address_q_cry_7\,
            carryinitout => \bfn_20_22_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_data_count_q_cry_7\,
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_16_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO\,
            carryinitout => \bfn_16_25_0_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIUKG82_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8027\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_583_g\
        );

    \this_reset_cond.M_stage_q_RNI6VB7_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__15770\,
            GLOBALBUFFEROUTPUT => \M_this_state_q_nss_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_start_data_delay.N_377_i_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__14874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15907\,
            lcout => \N_377_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILC1D4_9_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__14878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11988\,
            lcout => port_nmib_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7541\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7532\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.m27_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100100101"
        )
    port map (
            in0 => \N__18460\,
            in1 => \N__17926\,
            in2 => \N__18417\,
            in3 => \N__18308\,
            lcout => \N_28_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.m36_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110101110001"
        )
    port map (
            in0 => \N__18459\,
            in1 => \N__17925\,
            in2 => \N__18418\,
            in3 => \N__18309\,
            lcout => \N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.m55_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111101111"
        )
    port map (
            in0 => \N__18310\,
            in1 => \N__18461\,
            in2 => \N__17930\,
            in3 => \N__18412\,
            lcout => i7_mux_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_pixel_data_q_0_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__7510\,
            in1 => \N__7720\,
            in2 => \N__7780\,
            in3 => \N__7568\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_pixel_data_q_1_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__7719\,
            in1 => \N__7499\,
            in2 => \N__7486\,
            in3 => \N__7770\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_pixel_data_q_5_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__7722\,
            in1 => \N__7469\,
            in2 => \N__7453\,
            in3 => \N__7775\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_2_c_RNIIU2M1G_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7661\,
            in1 => \N__7859\,
            in2 => \N__7676\,
            in3 => \N__7850\,
            lcout => OPEN,
            ltout => \this_vga_signals.new_pixel_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_9_c_RNIKG4BDR1_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7583\,
            in1 => \N__7841\,
            in2 => \N__7652\,
            in3 => \N__7829\,
            lcout => debug_c_0,
            ltout => \debug_c_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_pixel_data_q_3_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011100"
        )
    port map (
            in0 => \N__7562\,
            in1 => \N__7636\,
            in2 => \N__7649\,
            in3 => \N__7721\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_pixel_data_q_4_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100110000"
        )
    port map (
            in0 => \N__7625\,
            in1 => \N__7724\,
            in2 => \N__7603\,
            in3 => \N__7774\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_1_c_RNI7QR2DF2_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7694\,
            in1 => \N__7685\,
            in2 => \_gnd_net_\,
            in3 => \N__7895\,
            lcout => OPEN,
            ltout => \this_vga_signals.new_pixel_1_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_5_c_RNIG1FT9B1_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__7904\,
            in1 => \N__7886\,
            in2 => \N__7586\,
            in3 => \N__7868\,
            lcout => \this_vga_signals.new_pixel_sx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIR31O3_0_9_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11993\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => this_vga_signals_vvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.m59_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010000"
        )
    port map (
            in0 => \N__17923\,
            in1 => \_gnd_net_\,
            in2 => \N__18467\,
            in3 => \N__18306\,
            lcout => \N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.m43_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000100110111"
        )
    port map (
            in0 => \N__18307\,
            in1 => \N__17922\,
            in2 => \N__18413\,
            in3 => \N__18462\,
            lcout => i7_mux,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIFBM6_7_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14111\,
            lcout => \this_vga_signals.M_hcounter_q_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIUTFM_6_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__10931\,
            in1 => \N__14789\,
            in2 => \_gnd_net_\,
            in3 => \N__14606\,
            lcout => \this_vga_signals.un4_hsynclt8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.m49_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101100111"
        )
    port map (
            in0 => \N__17924\,
            in1 => \N__18466\,
            in2 => \N__18419\,
            in3 => \N__18317\,
            lcout => OPEN,
            ltout => \N_50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_pixel_data_q_2_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100100010"
        )
    port map (
            in0 => \N__7738\,
            in1 => \N__7723\,
            in2 => \N__7796\,
            in3 => \N__7776\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIH8GJ4_9_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__11601\,
            in1 => \N__21390\,
            in2 => \_gnd_net_\,
            in3 => \N__11989\,
            lcout => \M_hcounter_q_esr_RNIH8GJ4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_0_c_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7958\,
            in2 => \N__9858\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_21_0_\,
            carryout => \this_vga_signals.new_pixel_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_0_c_RNIA47RND_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7964\,
            in2 => \N__11555\,
            in3 => \N__7688\,
            lcout => \this_vga_signals.new_pixel_1Z0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.new_pixel_1_cry_0\,
            carryout => \this_vga_signals.new_pixel_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_1_c_RNIRL8DV02_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8345\,
            in2 => \N__11480\,
            in3 => \N__7679\,
            lcout => \this_vga_signals.new_pixel_1_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.new_pixel_1_cry_1\,
            carryout => \this_vga_signals.new_pixel_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_2_c_RNIFPSJ9D_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8303\,
            in2 => \N__11150\,
            in3 => \N__7664\,
            lcout => \this_vga_signals.new_pixel_1_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.new_pixel_1_cry_2\,
            carryout => \this_vga_signals.new_pixel_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_3_c_RNITQA682_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8276\,
            in2 => \N__10997\,
            in3 => \N__7655\,
            lcout => \this_vga_signals.new_pixel_1_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.new_pixel_1_cry_3\,
            carryout => \this_vga_signals.new_pixel_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_4_c_RNI20CQL_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8261\,
            in2 => \N__14815\,
            in3 => \N__7889\,
            lcout => \this_vga_signals.new_pixel_1_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.new_pixel_1_cry_4\,
            carryout => \this_vga_signals.new_pixel_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_5_c_RNIJ8OH7_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8372\,
            in2 => \N__14607\,
            in3 => \N__7880\,
            lcout => \this_vga_signals.new_pixel_1_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.new_pixel_1_cry_5\,
            carryout => \this_vga_signals.new_pixel_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_6_c_RNI6UM51_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8435\,
            in2 => \N__7877\,
            in3 => \N__7862\,
            lcout => \this_vga_signals.new_pixel_1_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.new_pixel_1_cry_6\,
            carryout => \this_vga_signals.new_pixel_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_7_c_RNI22G7F_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8420\,
            in2 => \N__8399\,
            in3 => \N__7853\,
            lcout => \this_vga_signals.new_pixel_1_8\,
            ltout => OPEN,
            carryin => \bfn_6_22_0_\,
            carryout => \this_vga_signals.new_pixel_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_8_c_RNI48BK_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7952\,
            in2 => \N__20356\,
            in3 => \N__7844\,
            lcout => \this_vga_signals.new_pixel_1_9\,
            ltout => OPEN,
            carryin => \this_vga_signals.new_pixel_1_cry_8\,
            carryout => \this_vga_signals.new_pixel_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_9_c_RNI5ACK_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20312\,
            in2 => \N__7919\,
            in3 => \N__7835\,
            lcout => \this_vga_signals.new_pixel_1_10\,
            ltout => OPEN,
            carryin => \this_vga_signals.new_pixel_1_cry_9\,
            carryout => \this_vga_signals.new_pixel_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_10_c_RNID6631_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111111110"
        )
    port map (
            in0 => \N__14112\,
            in1 => \N__14298\,
            in2 => \N__14483\,
            in3 => \N__7832\,
            lcout => \this_vga_signals.new_pixel_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIC1312_9_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__7823\,
            in1 => \N__7910\,
            in2 => \N__14303\,
            in3 => \N__14476\,
            lcout => this_vga_signals_hsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIG53K_2_9_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => debug_c_i_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clock.M_counter_q_0_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8054\,
            lcout => \this_pixel_clock_M_counter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21632\,
            ce => 'H',
            sr => \N__21349\
        );

    \this_vga_signals.M_hcounter_q_0_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12853\,
            in2 => \_gnd_net_\,
            in3 => \N__9840\,
            lcout => \this_vga_signals.new_pixel_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21634\,
            ce => 'H',
            sr => \N__11341\
        );

    \this_vga_signals.M_hcounter_q_1_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__9839\,
            in1 => \_gnd_net_\,
            in2 => \N__12883\,
            in3 => \N__11513\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21634\,
            ce => 'H',
            sr => \N__11341\
        );

    \this_pixel_clock.M_counter_q_1_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8077\,
            in1 => \N__8059\,
            in2 => \_gnd_net_\,
            in3 => \N__21386\,
            lcout => \this_pixel_clock_M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21638\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIG53K_1_9_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14437\,
            in1 => \N__14283\,
            in2 => \_gnd_net_\,
            in3 => \N__14114\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNIG53K_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.G_296_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8076\,
            in1 => \N__8058\,
            in2 => \_gnd_net_\,
            in3 => \N__21385\,
            lcout => \this_vga_signals.GZ0Z_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNID96T_6_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__14591\,
            in1 => \N__10996\,
            in2 => \N__14816\,
            in3 => \N__14115\,
            lcout => \this_vga_signals.un3_hsynclt8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIG043KR2_0_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9559\,
            in1 => \N__9850\,
            in2 => \N__9593\,
            in3 => \N__9614\,
            lcout => \this_vga_signals.new_pixel_1_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIUA42ND_1_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8819\,
            lcout => \this_vga_signals.M_hcounter_q_RNIUA42NDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_cry_0_c_RNO_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__9613\,
            in1 => \N__9589\,
            in2 => \N__9859\,
            in3 => \N__9558\,
            lcout => \this_vga_signals.new_pixel_1_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIG53K_9_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__14470\,
            in1 => \N__14296\,
            in2 => \_gnd_net_\,
            in3 => \N__14113\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNIG53KZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_6_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11273\,
            lcout => \this_vga_signals.M_hcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21603\,
            ce => \N__9062\,
            sr => \N__11339\
        );

    \this_vga_signals.un4_haddress_g0_6_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111010111"
        )
    port map (
            in0 => \N__14198\,
            in1 => \N__14000\,
            in2 => \N__14397\,
            in3 => \N__14532\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_5_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7946\,
            in3 => \N__14750\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_1\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_2_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010111"
        )
    port map (
            in0 => \N__11124\,
            in1 => \N__10974\,
            in2 => \N__7943\,
            in3 => \N__8554\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11180\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21613\,
            ce => \N__9068\,
            sr => \N__11336\
        );

    \this_vga_signals.un4_haddress_g0_25_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111010111"
        )
    port map (
            in0 => \N__14199\,
            in1 => \N__14001\,
            in2 => \N__14398\,
            in3 => \N__14533\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_23_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7940\,
            in3 => \N__14751\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIHGHF3_9_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__12895\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11345\,
            lcout => \this_vga_signals.N_550_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_30_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100110011111"
        )
    port map (
            in0 => \N__13999\,
            in1 => \N__9144\,
            in2 => \N__14219\,
            in3 => \N__9187\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_28_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7997\,
            in3 => \N__14745\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_13_N_3L3_x0_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110100101"
        )
    port map (
            in0 => \N__7991\,
            in1 => \N__10161\,
            in2 => \N__10991\,
            in3 => \N__10032\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_13_N_3L3_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_13_N_3L3_ns_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7973\,
            in2 => \N__7994\,
            in3 => \N__10246\,
            lcout => \this_vga_signals.g0_13_N_3L3_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_13_N_3L3_x1_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100001"
        )
    port map (
            in0 => \N__10026\,
            in1 => \N__7990\,
            in2 => \N__10990\,
            in3 => \N__10160\,
            lcout => \this_vga_signals.g0_13_N_3L3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110101001011"
        )
    port map (
            in0 => \N__10965\,
            in1 => \N__14746\,
            in2 => \N__10051\,
            in3 => \N__10159\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_0\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_axb_4_l_fx_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8677\,
            in2 => \N__7967\,
            in3 => \N__9794\,
            lcout => \this_vga_signals.un1_haddress_0_axb_4_l_fxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010101"
        )
    port map (
            in0 => \N__10093\,
            in1 => \N__10162\,
            in2 => \N__10255\,
            in3 => \N__10033\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_address_buffer_q_esr_3_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8784\,
            in2 => \N__8201\,
            in3 => \N__9795\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21623\,
            ce => \N__15307\,
            sr => \N__15218\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIAV2K_6_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14741\,
            in1 => \N__14092\,
            in2 => \_gnd_net_\,
            in3 => \N__14564\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hcounter_d6lt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIBPF11_9_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14408\,
            in2 => \N__8087\,
            in3 => \N__14271\,
            lcout => \this_vga_signals.M_hcounter_d6_0\,
            ltout => \this_vga_signals.M_hcounter_d6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIUKG82_9_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__8084\,
            in1 => \N__8060\,
            in2 => \N__8030\,
            in3 => \N__21384\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNIUKG82Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_1_sx_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101101111"
        )
    port map (
            in0 => \N__11092\,
            in1 => \N__8620\,
            in2 => \N__11467\,
            in3 => \N__8598\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_ac0_1_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_1_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001101"
        )
    port map (
            in0 => \N__8599\,
            in1 => \N__11093\,
            in2 => \N__8003\,
            in3 => \N__8676\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_5_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11303\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21628\,
            ce => \N__9069\,
            sr => \N__11340\
        );

    \this_vga_signals.un4_haddress_if_m2_0_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000010010"
        )
    port map (
            in0 => \N__10932\,
            in1 => \N__14717\,
            in2 => \N__11123\,
            in3 => \N__10163\,
            lcout => \this_vga_signals.if_m2_0\,
            ltout => \this_vga_signals.if_m2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_x0_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010101001"
        )
    port map (
            in0 => \N__8630\,
            in1 => \N__8619\,
            in2 => \N__8000\,
            in3 => \N__8774\,
            lcout => \this_vga_signals.mult1_un75_sum_axb2_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_1_9_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110011001010"
        )
    port map (
            in0 => \N__14565\,
            in1 => \N__14267\,
            in2 => \N__14449\,
            in3 => \N__14093\,
            lcout => \this_vga_signals.un1_haddress_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_3_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__8573\,
            in1 => \N__10983\,
            in2 => \N__11143\,
            in3 => \N__9792\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_axb2_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_N_4_i_1_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011000100"
        )
    port map (
            in0 => \N__9536\,
            in1 => \N__9722\,
            in2 => \N__8228\,
            in3 => \N__9509\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_4_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_N_4_i_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14770\,
            in1 => \N__8225\,
            in2 => \N__8216\,
            in3 => \N__10208\,
            lcout => \this_vga_signals.N_4_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_i_3_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8786\,
            in1 => \N__8507\,
            in2 => \_gnd_net_\,
            in3 => \N__9793\,
            lcout => \this_vga_signals.mult1_un68_sum_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_1_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__11470\,
            in1 => \N__10439\,
            in2 => \N__11550\,
            in3 => \N__10396\,
            lcout => \this_vga_signals.mult1_un82_sum_ac0_1\,
            ltout => \this_vga_signals.mult1_un82_sum_ac0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001111011100"
        )
    port map (
            in0 => \N__10647\,
            in1 => \N__10580\,
            in2 => \N__8213\,
            in3 => \N__10670\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_axb_2_l_ofx_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__8210\,
            in1 => \N__10440\,
            in2 => \N__8204\,
            in3 => \N__10397\,
            lcout => \this_vga_signals.un1_haddress_0_axb_2_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_i_3_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__10398\,
            in1 => \_gnd_net_\,
            in2 => \N__10448\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un75_sum_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_axb_3_l_fx_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10446\,
            in1 => \N__9281\,
            in2 => \N__8320\,
            in3 => \N__10399\,
            lcout => \this_vga_signals.un1_haddress_0_axb_3_l_fxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIGF3C6_9_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8800\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8708\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9\,
            ltout => \this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TA7_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__8237\,
            in1 => \_gnd_net_\,
            in2 => \N__8375\,
            in3 => \N__8710\,
            lcout => \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TAZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TA7_0_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111111011111"
        )
    port map (
            in0 => \N__8709\,
            in1 => \N__8804\,
            in2 => \N__8452\,
            in3 => \N__8236\,
            lcout => \this_vga_signals.un1_haddress_0_cry_7_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_1_c_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8970\,
            in2 => \N__8951\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \this_vga_signals.un1_haddress_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44V02_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8360\,
            in2 => \N__8354\,
            in3 => \N__8333\,
            lcout => \this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44VZ0Z02\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_haddress_0_cry_1\,
            carryout => \this_vga_signals.un1_haddress_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9D_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8330\,
            in2 => \N__8324\,
            in3 => \N__8291\,
            lcout => \this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9DZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_haddress_0_cry_2\,
            carryout => \this_vga_signals.un1_haddress_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4T72_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8686\,
            in2 => \N__8288\,
            in3 => \N__8264\,
            lcout => \this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4TZ0Z72\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_haddress_0_cry_3\,
            carryout => \this_vga_signals.un1_haddress_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJL_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10222\,
            in2 => \N__8690\,
            in3 => \N__8249\,
            lcout => \this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJLZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_haddress_0_cry_4\,
            carryout => \this_vga_signals.un1_haddress_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_5_THRU_LUT4_0_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8711\,
            in2 => \N__8246\,
            in3 => \N__8456\,
            lcout => \this_vga_signals.un1_haddress_0_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_haddress_0_cry_5\,
            carryout => \this_vga_signals.un1_haddress_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQU_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8453\,
            in2 => \_gnd_net_\,
            in3 => \N__8423\,
            lcout => \this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQUZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_haddress_0_cry_6\,
            carryout => \this_vga_signals.un1_haddress_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBS7_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14292\,
            in1 => \N__14116\,
            in2 => \N__8419\,
            in3 => \N__8402\,
            lcout => \this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBSZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNI0EQT_6_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111111"
        )
    port map (
            in0 => \N__9245\,
            in1 => \N__8882\,
            in2 => \N__9424\,
            in3 => \N__9224\,
            lcout => \this_vga_signals.m8_0_1_tz\,
            ltout => \this_vga_signals.m8_0_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIGQG41_8_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__14177\,
            in1 => \_gnd_net_\,
            in2 => \N__8384\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__14790\,
            in1 => \N__9011\,
            in2 => \N__8381\,
            in3 => \N__9398\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_0_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010000000"
        )
    port map (
            in0 => \N__10975\,
            in1 => \N__10052\,
            in2 => \N__8378\,
            in3 => \N__10199\,
            lcout => \this_vga_signals.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_7_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11242\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21596\,
            ce => \N__9076\,
            sr => \N__11334\
        );

    \this_vga_signals.M_hcounter_q_esr_8_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11219\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21596\,
            ce => \N__9076\,
            sr => \N__11334\
        );

    \this_vga_signals.M_hcounter_q_9_rep1_esr_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11179\,
            lcout => \this_vga_signals.M_hcounter_q_9_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21596\,
            ce => \N__9076\,
            sr => \N__11334\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNIN6RR_7_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9133\,
            in2 => \N__9231\,
            in3 => \N__9179\,
            lcout => \this_vga_signals.M_hcounter_q_fast_esr_RNIN6RRZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_7_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11243\,
            lcout => \this_vga_signals.M_hcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21596\,
            ce => \N__9076\,
            sr => \N__11334\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNIPO3M_7_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100000000"
        )
    port map (
            in0 => \N__9358\,
            in1 => \_gnd_net_\,
            in2 => \N__9232\,
            in3 => \N__9135\,
            lcout => \this_vga_signals.N_75\,
            ltout => \this_vga_signals.N_75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_x1_1_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111001001"
        )
    port map (
            in0 => \N__14530\,
            in1 => \N__8885\,
            in2 => \N__8483\,
            in3 => \N__8480\,
            lcout => \this_vga_signals.mult1_un54_sum_m_x1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_1_1_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000101011"
        )
    port map (
            in0 => \N__9357\,
            in1 => \N__9134\,
            in2 => \N__8913\,
            in3 => \N__9180\,
            lcout => \this_vga_signals.mult1_un54_sum_m_1_1\,
            ltout => \this_vga_signals.mult1_un54_sum_m_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_x0_1_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001100110"
        )
    port map (
            in0 => \N__14531\,
            in1 => \N__8886\,
            in2 => \N__8474\,
            in3 => \N__8471\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_m_x0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_ns_1_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8924\,
            in2 => \N__8465\,
            in3 => \N__8462\,
            lcout => \this_vga_signals.mult1_un54_sum_m_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_6_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11272\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21605\,
            ce => \N__9054\,
            sr => \N__11337\
        );

    \this_vga_signals.M_hcounter_q_6_rep1_esr_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11271\,
            lcout => \this_vga_signals.M_hcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21605\,
            ce => \N__9054\,
            sr => \N__11337\
        );

    \this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOM71_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100100001001"
        )
    port map (
            in0 => \N__9145\,
            in1 => \N__8914\,
            in2 => \N__9188\,
            in3 => \N__8887\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOMZ0Z71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_8_rep1_esr_RNI1Q1C1_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__20360\,
            in1 => \_gnd_net_\,
            in2 => \N__8522\,
            in3 => \N__9369\,
            lcout => \this_vga_signals.m8_0_2\,
            ltout => \this_vga_signals.m8_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_1_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__10963\,
            in1 => \N__8888\,
            in2 => \N__8519\,
            in3 => \N__9335\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_1\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101100"
        )
    port map (
            in0 => \N__10027\,
            in1 => \N__10086\,
            in2 => \N__8516\,
            in3 => \N__10164\,
            lcout => \this_vga_signals.mult1_un61_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_8_rep1_esr_RNIKFGM4_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__9370\,
            in1 => \N__9393\,
            in2 => \N__8942\,
            in3 => \N__9005\,
            lcout => \this_vga_signals.mult1_un54_sum_i_0_3\,
            ltout => \this_vga_signals.mult1_un54_sum_i_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_31_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111110101"
        )
    port map (
            in0 => \N__14740\,
            in1 => \_gnd_net_\,
            in2 => \N__8513\,
            in3 => \N__10964\,
            lcout => \this_vga_signals.g1_6_0\,
            ltout => \this_vga_signals.g1_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_13_N_2L1_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8510\,
            in3 => \N__10028\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_13_N_2L1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_13_N_4L5_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000100010010"
        )
    port map (
            in0 => \N__8503\,
            in1 => \N__8492\,
            in2 => \N__8486\,
            in3 => \N__9779\,
            lcout => \this_vga_signals.g0_13_N_4L5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011000001001"
        )
    port map (
            in0 => \N__8663\,
            in1 => \N__8621\,
            in2 => \N__8600\,
            in3 => \N__8776\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_x1_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010010101"
        )
    port map (
            in0 => \N__11088\,
            in1 => \N__8777\,
            in2 => \N__10992\,
            in3 => \N__8664\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_3_0_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_0_0_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11087\,
            lcout => \this_vga_signals.mult1_un75_sum_axb2_0_0\,
            ltout => \this_vga_signals.mult1_un75_sum_axb2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_x1_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010100101"
        )
    port map (
            in0 => \N__8775\,
            in1 => \N__8593\,
            in2 => \N__8624\,
            in3 => \N__8618\,
            lcout => \this_vga_signals.mult1_un75_sum_axb2_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI43A65_5_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110100101"
        )
    port map (
            in0 => \N__14752\,
            in1 => \N__9006\,
            in2 => \N__10972\,
            in3 => \N__9334\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5\,
            ltout => \this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_3_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8594\,
            in2 => \N__8576\,
            in3 => \N__8662\,
            lcout => \this_vga_signals.mult1_un68_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_10_3_0_a2_0_0_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010111101"
        )
    port map (
            in0 => \N__14753\,
            in1 => \N__10201\,
            in2 => \N__10973\,
            in3 => \N__10060\,
            lcout => \this_vga_signals.g0_10_3_0_a2_0_0\,
            ltout => \this_vga_signals.g0_10_3_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_1_3_a2_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100011110"
        )
    port map (
            in0 => \N__8567\,
            in1 => \N__8555\,
            in2 => \N__8540\,
            in3 => \N__9780\,
            lcout => \this_vga_signals.mult1_un68_sum_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__11131\,
            in1 => \_gnd_net_\,
            in2 => \N__9796\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un75_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_ns_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8537\,
            in2 => \N__8531\,
            in3 => \N__8678\,
            lcout => \this_vga_signals.mult1_un75_sum_axb2_i\,
            ltout => \this_vga_signals.mult1_un75_sum_axb2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc2_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000101101"
        )
    port map (
            in0 => \N__9271\,
            in1 => \N__11132\,
            in2 => \N__8789\,
            in3 => \N__8734\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_x0_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101100101101"
        )
    port map (
            in0 => \N__10982\,
            in1 => \N__8785\,
            in2 => \N__11144\,
            in3 => \N__8679\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_ac0_3_0_1_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_ns_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8744\,
            in2 => \N__8738\,
            in3 => \N__9781\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_3_0_1\,
            ltout => \this_vga_signals.mult1_un75_sum_ac0_3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111101011"
        )
    port map (
            in0 => \N__8735\,
            in1 => \N__9272\,
            in2 => \N__8726\,
            in3 => \N__8723\,
            lcout => \this_vga_signals.mult1_un75_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10445\,
            in2 => \N__10411\,
            in3 => \N__8717\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_0_9_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101100101000"
        )
    port map (
            in0 => \N__14266\,
            in1 => \N__14077\,
            in2 => \N__14472\,
            in3 => \N__14578\,
            lcout => \this_vga_signals.N_510_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axb2_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8851\,
            in1 => \N__11469\,
            in2 => \N__10410\,
            in3 => \N__10444\,
            lcout => \this_vga_signals.mult1_un82_sum_axb2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_1_0_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__11148\,
            in1 => \N__10980\,
            in2 => \_gnd_net_\,
            in3 => \N__8680\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14801\,
            in1 => \N__9277\,
            in2 => \N__8633\,
            in3 => \N__10202\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_1_i\,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_0_0_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001100100"
        )
    port map (
            in0 => \N__11468\,
            in1 => \N__8852\,
            in2 => \N__8843\,
            in3 => \N__10400\,
            lcout => \this_vga_signals.mult1_un82_sum_ac0_3_0_0\,
            ltout => \this_vga_signals.mult1_un82_sum_ac0_3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_i_3_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011011000011"
        )
    port map (
            in0 => \N__10651\,
            in1 => \N__10671\,
            in2 => \N__8840\,
            in3 => \N__10611\,
            lcout => \this_vga_signals.un1_haddress_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI5HOBQC_1_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10672\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11541\,
            lcout => \this_vga_signals.M_hcounter_q_RNI5HOBQCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIPIQRNR_2_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111110010110"
        )
    port map (
            in0 => \N__11476\,
            in1 => \N__10649\,
            in2 => \N__10586\,
            in3 => \N__10612\,
            lcout => \this_vga_signals.M_hcounter_q_RNIPIQRNRZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.new_pixel_1_axb_1_N_4L5_x1_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110011001"
        )
    port map (
            in0 => \N__10650\,
            in1 => \N__10584\,
            in2 => \_gnd_net_\,
            in3 => \N__10610\,
            lcout => OPEN,
            ltout => \this_vga_signals.new_pixel_1_axb_1_N_4L5_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI8TTVN32_2_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__9466\,
            in1 => \_gnd_net_\,
            in2 => \N__8837\,
            in3 => \N__8834\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hcounter_q_RNI8TTVN32Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIU31PMD_1_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8828\,
            in1 => \N__8971\,
            in2 => \N__8822\,
            in3 => \N__9582\,
            lcout => \this_vga_signals.new_pixel_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_9_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010011010111"
        )
    port map (
            in0 => \N__14265\,
            in1 => \N__14076\,
            in2 => \N__14471\,
            in3 => \N__14577\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIIV9H5_9_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8807\,
            in3 => \N__10221\,
            lcout => \this_vga_signals.un1_haddress_0_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_4_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101101010100"
        )
    port map (
            in0 => \N__10609\,
            in1 => \N__11475\,
            in2 => \N__9467\,
            in3 => \N__10648\,
            lcout => \this_vga_signals.mult1_un89_sum_axbxc3_0\,
            ltout => \this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_haddress_0_cry_1_c_RNO_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__8972\,
            in1 => \N__9581\,
            in2 => \N__8954\,
            in3 => \N__9549\,
            lcout => \this_vga_signals.un1_haddress_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIGQG41_0_8_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8938\,
            in2 => \_gnd_net_\,
            in3 => \N__14178\,
            lcout => \this_vga_signals.g1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNI58601_7_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100100000"
        )
    port map (
            in0 => \N__9367\,
            in1 => \N__9142\,
            in2 => \N__9233\,
            in3 => \N__9185\,
            lcout => \this_vga_signals.ANC2_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_8_rep1_esr_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11218\,
            lcout => \this_vga_signals.M_hcounter_q_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21590\,
            ce => \N__9077\,
            sr => \N__11333\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_2_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111010111"
        )
    port map (
            in0 => \N__9368\,
            in1 => \N__9143\,
            in2 => \N__8915\,
            in3 => \N__9186\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__8884\,
            in1 => \_gnd_net_\,
            in2 => \N__8918\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_7_rep1_esr_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11241\,
            lcout => \this_vga_signals.M_hcounter_q_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21590\,
            ce => \N__9077\,
            sr => \N__11333\
        );

    \this_vga_signals.M_hcounter_q_5_rep1_esr_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11302\,
            lcout => \this_vga_signals.M_hcounter_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21590\,
            ce => \N__9077\,
            sr => \N__11333\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNI52HL_9_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__9244\,
            in1 => \N__8883\,
            in2 => \_gnd_net_\,
            in3 => \N__9222\,
            lcout => \this_vga_signals.M_hcounter_q_fast_esr_RNI52HLZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_9_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11178\,
            lcout => \this_vga_signals.M_hcounter_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21590\,
            ce => \N__9077\,
            sr => \N__11333\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNIHH441_5_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101001011"
        )
    port map (
            in0 => \N__9223\,
            in1 => \N__9181\,
            in2 => \N__9146\,
            in3 => \N__9089\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hcounter_q_fast_esr_RNIHH441Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNI56982_8_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9083\,
            in2 => \N__9098\,
            in3 => \N__9095\,
            lcout => \this_vga_signals.m8_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_5_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11301\,
            lcout => \this_vga_signals.M_hcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21597\,
            ce => \N__9058\,
            sr => \N__11335\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_8_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11217\,
            lcout => \this_vga_signals.M_hcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21597\,
            ce => \N__9058\,
            sr => \N__11335\
        );

    \this_vga_signals.un4_haddress_g0_17_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__9392\,
            in1 => \N__9010\,
            in2 => \N__14813\,
            in3 => \N__8984\,
            lcout => \this_vga_signals.g1_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g4_1_1_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__10049\,
            in1 => \N__10171\,
            in2 => \_gnd_net_\,
            in3 => \N__10251\,
            lcout => OPEN,
            ltout => \this_vga_signals.g4_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g4_1_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000011111"
        )
    port map (
            in0 => \N__14798\,
            in1 => \N__9323\,
            in2 => \N__8975\,
            in3 => \N__10907\,
            lcout => \this_vga_signals.g4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_8_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111010111"
        )
    port map (
            in0 => \N__14263\,
            in1 => \N__14038\,
            in2 => \N__14479\,
            in3 => \N__14534\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_0_a2_0_0_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101001011001"
        )
    port map (
            in0 => \N__10050\,
            in1 => \N__10908\,
            in2 => \N__10200\,
            in3 => \N__14799\,
            lcout => \this_vga_signals.g1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNIJLEA3_6_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__9428\,
            in1 => \N__9407\,
            in2 => \N__9397\,
            in3 => \N__9371\,
            lcout => \this_vga_signals.m8_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_16_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111010111"
        )
    port map (
            in0 => \N__14264\,
            in1 => \N__14039\,
            in2 => \N__14480\,
            in3 => \N__14535\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_14_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010000000"
        )
    port map (
            in0 => \N__10170\,
            in1 => \N__10909\,
            in2 => \N__9317\,
            in3 => \N__10055\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_21_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100110111"
        )
    port map (
            in0 => \N__9308\,
            in1 => \N__11116\,
            in2 => \N__9296\,
            in3 => \N__10945\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_0_a2_0_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010011011011"
        )
    port map (
            in0 => \N__10168\,
            in1 => \N__14754\,
            in2 => \N__10979\,
            in3 => \N__10054\,
            lcout => \this_vga_signals.N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_29_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10056\,
            in1 => \N__9293\,
            in2 => \N__10793\,
            in3 => \N__9791\,
            lcout => \this_vga_signals.mult1_un75_sum_axb2_i_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g4_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010010"
        )
    port map (
            in0 => \N__9287\,
            in1 => \N__9273\,
            in2 => \N__11142\,
            in3 => \N__9507\,
            lcout => \this_vga_signals.g4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_9_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__11418\,
            in1 => \N__11117\,
            in2 => \_gnd_net_\,
            in3 => \N__9790\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_1_1\,
            ltout => \this_vga_signals.mult1_un75_sum_ac0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_13_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__11118\,
            in1 => \N__9524\,
            in2 => \N__9518\,
            in3 => \N__9506\,
            lcout => \this_vga_signals.g1_1_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_1_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__10053\,
            in1 => \N__10250\,
            in2 => \_gnd_net_\,
            in3 => \N__10169\,
            lcout => \this_vga_signals.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_0_2_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9515\,
            in1 => \N__10215\,
            in2 => \N__14814\,
            in3 => \N__9508\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_12_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110101111000"
        )
    port map (
            in0 => \N__9488\,
            in1 => \N__9482\,
            in2 => \N__9476\,
            in3 => \N__9473\,
            lcout => \this_vga_signals.N_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_7_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9452\,
            in2 => \_gnd_net_\,
            in3 => \N__14800\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_2_0_a2_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101010110"
        )
    port map (
            in0 => \N__9730\,
            in1 => \N__9655\,
            in2 => \N__9443\,
            in3 => \N__9786\,
            lcout => \this_vga_signals.mult1_un68_sum_0_3\,
            ltout => \this_vga_signals.mult1_un68_sum_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_0_a2_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101001000101"
        )
    port map (
            in0 => \N__9707\,
            in1 => \N__11110\,
            in2 => \N__9440\,
            in3 => \N__9437\,
            lcout => \this_vga_signals.g1_0_a2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_11_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__11471\,
            in1 => \N__11085\,
            in2 => \_gnd_net_\,
            in3 => \N__9785\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_12_0_a2_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11086\,
            in1 => \N__10981\,
            in2 => \N__9797\,
            in3 => \N__9731\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_axb2_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_1_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100011001"
        )
    port map (
            in0 => \N__9721\,
            in1 => \N__9633\,
            in2 => \N__9710\,
            in3 => \N__9706\,
            lcout => \this_vga_signals.mult1_un75_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_x2_0_0_a2_3_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9644\,
            in1 => \N__10220\,
            in2 => \N__9677\,
            in3 => \N__9635\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_i_x2_0_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000110"
        )
    port map (
            in0 => \N__11549\,
            in1 => \N__9854\,
            in2 => \N__9698\,
            in3 => \N__9694\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_i4_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011011110110"
        )
    port map (
            in0 => \N__9695\,
            in1 => \N__9620\,
            in2 => \N__9686\,
            in3 => \N__9683\,
            lcout => \this_vga_signals.mult1_un89_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_x2_0_0_a2_0_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11445\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14802\,
            lcout => \this_vga_signals.g0_i_x2_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_10_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010111"
        )
    port map (
            in0 => \N__11149\,
            in1 => \N__10923\,
            in2 => \N__9668\,
            in3 => \N__9659\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0\,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_0_a2_4_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11378\,
            in1 => \N__10219\,
            in2 => \N__9638\,
            in3 => \N__9634\,
            lcout => \this_vga_signals.g0_0_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_address_buffer_q_esr_0_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__9607\,
            in1 => \N__9588\,
            in2 => \_gnd_net_\,
            in3 => \N__9563\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21629\,
            ce => \N__15292\,
            sr => \N__15204\
        );

    \this_vga_signals.M_address_buffer_q_esr_1_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100101"
        )
    port map (
            in0 => \N__10673\,
            in1 => \N__10652\,
            in2 => \N__10622\,
            in3 => \N__10585\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21629\,
            ce => \N__15292\,
            sr => \N__15204\
        );

    \this_vga_signals.M_address_buffer_q_esr_2_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10447\,
            in2 => \_gnd_net_\,
            in3 => \N__10412\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21629\,
            ce => \N__15292\,
            sr => \N__15204\
        );

    \this_vga_signals.M_address_buffer_q_esr_4_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111000"
        )
    port map (
            in0 => \N__10259\,
            in1 => \N__10223\,
            in2 => \N__10094\,
            in3 => \N__10061\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21633\,
            ce => \N__15306\,
            sr => \N__15197\
        );

    \this_vga_signals.M_address_buffer_q_esr_12_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__11789\,
            in1 => \N__11822\,
            in2 => \N__11807\,
            in3 => \N__11774\,
            lcout => \M_this_vga_signals_address_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21598\,
            ce => \N__15268\,
            sr => \N__15179\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9860\,
            in2 => \N__11554\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12921\,
            in1 => \N__11441\,
            in2 => \_gnd_net_\,
            in3 => \N__9806\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__21606\,
            ce => 'H',
            sr => \N__11338\
        );

    \this_vga_signals.M_hcounter_q_3_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12896\,
            in1 => \N__11122\,
            in2 => \_gnd_net_\,
            in3 => \N__9803\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__21606\,
            ce => 'H',
            sr => \N__11338\
        );

    \this_vga_signals.M_hcounter_q_4_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12922\,
            in1 => \N__10910\,
            in2 => \_gnd_net_\,
            in3 => \N__9800\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__21606\,
            ce => 'H',
            sr => \N__11338\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRD_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14758\,
            in2 => \_gnd_net_\,
            in3 => \N__11276\,
            lcout => \this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRDZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSD_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14602\,
            in2 => \_gnd_net_\,
            in3 => \N__11246\,
            lcout => \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTD_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14098\,
            in2 => \_gnd_net_\,
            in3 => \N__11222\,
            lcout => \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUD_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14279\,
            in2 => \_gnd_net_\,
            in3 => \N__11186\,
            lcout => \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVD_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14463\,
            in2 => \_gnd_net_\,
            in3 => \N__11183\,
            lcout => \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU45J5_9_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__11573\,
            in1 => \N__12884\,
            in2 => \_gnd_net_\,
            in3 => \N__11972\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIH06Q6_9_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12885\,
            in2 => \_gnd_net_\,
            in3 => \N__15126\,
            lcout => \this_vga_signals.N_550_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_4_0_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11084\,
            in2 => \_gnd_net_\,
            in3 => \N__10906\,
            lcout => \this_vga_signals.g0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIG53K_0_9_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__14462\,
            in1 => \N__14278\,
            in2 => \_gnd_net_\,
            in3 => \N__14097\,
            lcout => debug_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_0_a2_1_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11548\,
            in1 => \N__11446\,
            in2 => \_gnd_net_\,
            in3 => \N__14791\,
            lcout => \this_vga_signals.g0_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11357\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11372\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21617\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000101101"
        )
    port map (
            in0 => \N__13036\,
            in1 => \N__13453\,
            in2 => \N__13289\,
            in3 => \N__13222\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_0_0\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m7_0_o4_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011101000"
        )
    port map (
            in0 => \N__13114\,
            in1 => \N__13199\,
            in2 => \N__11351\,
            in3 => \N__11837\,
            lcout => \this_vga_signals.if_N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__11896\,
            in1 => \N__11871\,
            in2 => \_gnd_net_\,
            in3 => \N__11931\,
            lcout => \this_vga_signals.mult1_un40_sum_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_4_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100010000100"
        )
    port map (
            in0 => \N__11932\,
            in1 => \N__12809\,
            in2 => \N__11878\,
            in3 => \N__11897\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11911\,
            in2 => \_gnd_net_\,
            in3 => \N__11918\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3\,
            ltout => \this_vga_signals.mult1_un47_sum_ac0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__11802\,
            in1 => \N__11821\,
            in2 => \N__11348\,
            in3 => \N__11772\,
            lcout => \this_vga_signals.mult1_un47_sum_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_2_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__11933\,
            in1 => \_gnd_net_\,
            in2 => \N__11879\,
            in3 => \N__12808\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_1_2\,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc3_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_0_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__13021\,
            in1 => \_gnd_net_\,
            in2 => \N__11810\,
            in3 => \N__13452\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__11803\,
            in1 => \N__11788\,
            in2 => \N__11777\,
            in3 => \N__11773\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010101"
        )
    port map (
            in0 => \N__13025\,
            in1 => \N__13198\,
            in2 => \N__12718\,
            in3 => \N__13121\,
            lcout => \this_vga_signals.un2_vsynclt8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI6CLG4_5_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__13454\,
            in1 => \N__11945\,
            in2 => \N__11759\,
            in3 => \N__13739\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_address_buffer_q_esr_6_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010110111000"
        )
    port map (
            in0 => \N__14302\,
            in1 => \N__14117\,
            in2 => \N__14615\,
            in3 => \N__14478\,
            lcout => \M_this_vga_signals_address_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21615\,
            ce => \N__15299\,
            sr => \N__15183\
        );

    \this_vga_signals.un5_vaddress_if_m7_0_m2_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000011111001"
        )
    port map (
            in0 => \N__13033\,
            in1 => \N__12490\,
            in2 => \N__13124\,
            in3 => \N__11621\,
            lcout => \this_vga_signals.if_N_10\,
            ltout => \this_vga_signals.if_N_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12330\,
            in1 => \N__12346\,
            in2 => \N__11615\,
            in3 => \N__12186\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_0_0\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_c2_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101010000"
        )
    port map (
            in0 => \N__13202\,
            in1 => \_gnd_net_\,
            in2 => \N__11612\,
            in3 => \N__12713\,
            lcout => \this_vga_signals.mult1_un75_sum_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__13120\,
            in1 => \N__13200\,
            in2 => \_gnd_net_\,
            in3 => \N__12187\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_ns_1_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13201\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12147\,
            lcout => \this_vga_signals.mult1_un82_sum_c3_0_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__11836\,
            in1 => \_gnd_net_\,
            in2 => \N__13037\,
            in3 => \N__12487\,
            lcout => \this_vga_signals.mult1_un61_sum_axb2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__13026\,
            in1 => \N__13445\,
            in2 => \_gnd_net_\,
            in3 => \N__13220\,
            lcout => \this_vga_signals.mult1_un54_sum_c2\,
            ltout => \this_vga_signals.mult1_un54_sum_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110101000010"
        )
    port map (
            in0 => \N__13221\,
            in1 => \N__13281\,
            in2 => \N__11846\,
            in3 => \N__13258\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__13028\,
            in1 => \_gnd_net_\,
            in2 => \N__11843\,
            in3 => \N__13115\,
            lcout => \this_vga_signals.mult1_un61_sum_c2\,
            ltout => \this_vga_signals.mult1_un61_sum_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001001"
        )
    port map (
            in0 => \N__12488\,
            in1 => \N__12502\,
            in2 => \N__11840\,
            in3 => \N__12520\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_0_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13032\,
            in1 => \N__13116\,
            in2 => \_gnd_net_\,
            in3 => \N__12489\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13027\,
            in2 => \_gnd_net_\,
            in3 => \N__11835\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI48605_9_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111110011101"
        )
    port map (
            in0 => \N__13335\,
            in1 => \N__13817\,
            in2 => \N__11870\,
            in3 => \N__12004\,
            lcout => \this_vga_signals.SUM_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_0_3_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110011111"
        )
    port map (
            in0 => \N__15070\,
            in1 => \N__15456\,
            in2 => \N__12776\,
            in3 => \N__13805\,
            lcout => \this_vga_signals.mult1_un47_sum_axb2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011100001110"
        )
    port map (
            in0 => \N__13018\,
            in1 => \N__13428\,
            in2 => \N__12807\,
            in3 => \N__15071\,
            lcout => \this_vga_signals.mult1_un47_sum_c2\,
            ltout => \this_vga_signals.mult1_un47_sum_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_0_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100000111100"
        )
    port map (
            in0 => \N__11885\,
            in1 => \N__11912\,
            in2 => \N__11900\,
            in3 => \N__15457\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI87V41_6_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__13017\,
            in1 => \N__15069\,
            in2 => \_gnd_net_\,
            in3 => \N__13427\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_4_tz_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111110111"
        )
    port map (
            in0 => \N__15072\,
            in1 => \N__13806\,
            in2 => \N__13738\,
            in3 => \N__13336\,
            lcout => \this_vga_signals.mult1_un47_sum_axb2_3_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNI94581_6_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000010011"
        )
    port map (
            in0 => \N__13425\,
            in1 => \N__15391\,
            in2 => \N__13034\,
            in3 => \N__13722\,
            lcout => \this_vga_signals.vaddress_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_1_6_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13721\,
            in1 => \N__15447\,
            in2 => \N__15068\,
            in3 => \N__13794\,
            lcout => \this_vga_signals.vaddress_c5_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__12742\,
            in1 => \N__13080\,
            in2 => \N__12712\,
            in3 => \N__13192\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_d7lt8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIBJQP3_6_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__15050\,
            in1 => \N__12014\,
            in2 => \N__11849\,
            in3 => \N__13795\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_d7lt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI8MOD6_9_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__12916\,
            in1 => \N__13337\,
            in2 => \N__12017\,
            in3 => \N__12765\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI0IM71_5_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__13426\,
            in1 => \_gnd_net_\,
            in2 => \N__13035\,
            in3 => \N__13723\,
            lcout => \this_vga_signals.M_vcounter_d7lto8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_0_6_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__15458\,
            in1 => \N__13796\,
            in2 => \N__15083\,
            in3 => \N__13727\,
            lcout => OPEN,
            ltout => \this_vga_signals.un6_vvisibilitylt9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIR31O3_9_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13329\,
            in2 => \N__12008\,
            in3 => \N__12005\,
            lcout => \this_vga_signals.vvisibility\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_a5_1_0_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__13330\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13797\,
            lcout => OPEN,
            ltout => \this_vga_signals.vsync_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIP8HU1_6_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__13181\,
            in1 => \N__15082\,
            in2 => \N__11948\,
            in3 => \N__13010\,
            lcout => \this_vga_signals.vsync_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIRHPK7_9_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__14931\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12917\,
            lcout => \this_vga_signals.N_550_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13370\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21607\,
            ce => \N__14990\,
            sr => \N__14957\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_ns_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100000001111"
        )
    port map (
            in0 => \N__12743\,
            in1 => \N__12353\,
            in2 => \N__12719\,
            in3 => \N__11939\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_address_buffer_q_esr_7_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12656\,
            in1 => \N__12527\,
            in2 => \N__12650\,
            in3 => \N__12191\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21579\,
            ce => \N__15329\,
            sr => \N__15216\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_ac0_3_0_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011011100"
        )
    port map (
            in0 => \N__13196\,
            in1 => \N__12536\,
            in2 => \N__12717\,
            in3 => \N__12148\,
            lcout => \this_vga_signals.mult1_un75_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un75_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_i_1_3_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13113\,
            in1 => \N__13197\,
            in2 => \N__12530\,
            in3 => \N__12164\,
            lcout => \this_vga_signals.mult1_un82_sum_i_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_address_buffer_q_esr_10_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000011100011110"
        )
    port map (
            in0 => \N__12521\,
            in1 => \N__12331\,
            in2 => \N__12509\,
            in3 => \N__12491\,
            lcout => \M_this_vga_signals_address_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21582\,
            ce => \N__15327\,
            sr => \N__15193\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_bm_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001001"
        )
    port map (
            in0 => \N__13194\,
            in1 => \N__12199\,
            in2 => \N__13122\,
            in3 => \N__12188\,
            lcout => \this_vga_signals.mult1_un82_sum_c3_0_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_address_buffer_q_esr_9_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12190\,
            in1 => \N__12347\,
            in2 => \N__12335\,
            in3 => \N__12317\,
            lcout => \M_this_vga_signals_address_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21582\,
            ce => \N__15327\,
            sr => \N__15193\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001100111001"
        )
    port map (
            in0 => \N__13195\,
            in1 => \N__12200\,
            in2 => \N__13123\,
            in3 => \N__12189\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc2\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_address_buffer_q_esr_8_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12158\,
            in2 => \N__12152\,
            in3 => \N__12149\,
            lcout => \M_this_vga_signals_address_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21582\,
            ce => \N__15327\,
            sr => \N__15193\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011000"
        )
    port map (
            in0 => \N__15445\,
            in1 => \N__15384\,
            in2 => \N__15409\,
            in3 => \N__15340\,
            lcout => \this_vga_signals.mult1_un40_sum_c3\,
            ltout => \this_vga_signals.mult1_un40_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__15073\,
            in1 => \N__13019\,
            in2 => \N__12785\,
            in3 => \N__13424\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__13717\,
            in1 => \N__13332\,
            in2 => \N__13808\,
            in3 => \N__15383\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_x0_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__15382\,
            in1 => \N__13799\,
            in2 => \_gnd_net_\,
            in3 => \N__13716\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_ns_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__13423\,
            in1 => \_gnd_net_\,
            in2 => \N__12782\,
            in3 => \N__13664\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_3_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110100"
        )
    port map (
            in0 => \N__13333\,
            in1 => \N__13803\,
            in2 => \N__12779\,
            in3 => \N__13718\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_0_3_1_1_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010011001"
        )
    port map (
            in0 => \N__13334\,
            in1 => \N__13804\,
            in2 => \_gnd_net_\,
            in3 => \N__13719\,
            lcout => \this_vga_signals.mult1_un47_sum_axb2_0_3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12919\,
            in1 => \N__12738\,
            in2 => \N__12767\,
            in3 => \N__12766\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__21588\,
            ce => 'H',
            sr => \N__14932\
        );

    \this_vga_signals.M_vcounter_q_1_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12923\,
            in1 => \N__12690\,
            in2 => \_gnd_net_\,
            in3 => \N__12659\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__21588\,
            ce => 'H',
            sr => \N__14932\
        );

    \this_vga_signals.M_vcounter_q_2_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12920\,
            in1 => \N__13193\,
            in2 => \_gnd_net_\,
            in3 => \N__13127\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__21588\,
            ce => 'H',
            sr => \N__14932\
        );

    \this_vga_signals.M_vcounter_q_3_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12924\,
            in1 => \N__13086\,
            in2 => \_gnd_net_\,
            in3 => \N__13040\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__21588\,
            ce => 'H',
            sr => \N__14932\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13020\,
            in2 => \_gnd_net_\,
            in3 => \N__12938\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12925\,
            in1 => \N__13438\,
            in2 => \_gnd_net_\,
            in3 => \N__12935\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \N__21588\,
            ce => 'H',
            sr => \N__14932\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15067\,
            in2 => \_gnd_net_\,
            in3 => \N__12932\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12926\,
            in1 => \N__13728\,
            in2 => \_gnd_net_\,
            in3 => \N__12929\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \N__21588\,
            ce => 'H',
            sr => \N__14932\
        );

    \this_vga_signals.M_vcounter_q_8_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12918\,
            in1 => \N__13798\,
            in2 => \_gnd_net_\,
            in3 => \N__12812\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \N__21591\,
            ce => 'H',
            sr => \N__14936\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_0_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20255\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_1_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__20316\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_0_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_2_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20259\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_1_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_3_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__20317\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_2_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_4_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20263\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_3_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_5_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__20318\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_4_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_6_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20267\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_5_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13331\,
            in2 => \_gnd_net_\,
            in3 => \N__13340\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21599\,
            ce => \N__15003\,
            sr => \N__14965\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2_9_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101101111000"
        )
    port map (
            in0 => \N__14258\,
            in1 => \N__14102\,
            in2 => \N__14481\,
            in3 => \N__14608\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_address_buffer_q_esr_11_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011010010011"
        )
    port map (
            in0 => \N__13282\,
            in1 => \N__13262\,
            in2 => \N__13241\,
            in3 => \N__13229\,
            lcout => \M_this_vga_signals_address_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21578\,
            ce => \N__15328\,
            sr => \N__15217\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_6_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001001"
        )
    port map (
            in0 => \N__15435\,
            in1 => \N__13807\,
            in2 => \N__15051\,
            in3 => \N__13720\,
            lcout => \this_vga_signals.vaddress_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_x1_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__13354\,
            in1 => \N__13790\,
            in2 => \N__15381\,
            in3 => \N__13715\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_dmab_c_sbtinv_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14861\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => port_dmab_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIP3JE_4_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13422\,
            lcout => \this_vga_signals.vaddress_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15097\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21587\,
            ce => \N__15007\,
            sr => \N__14966\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13366\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21587\,
            ce => \N__15007\,
            sr => \N__14966\
        );

    \M_this_data_count_q_0_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15641\,
            in2 => \N__20047\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => \un1_M_this_data_count_q_cry_0\,
            clk => \N__21595\,
            ce => 'H',
            sr => \N__15482\
        );

    \M_this_data_count_q_1_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20011\,
            in2 => \N__15701\,
            in3 => \N__13346\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_0\,
            carryout => \un1_M_this_data_count_q_cry_1\,
            clk => \N__21595\,
            ce => 'H',
            sr => \N__15482\
        );

    \M_this_data_count_q_2_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15671\,
            in2 => \N__20048\,
            in3 => \N__13343\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_1\,
            carryout => \un1_M_this_data_count_q_cry_2\,
            clk => \N__21595\,
            ce => 'H',
            sr => \N__15482\
        );

    \M_this_data_count_q_3_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20015\,
            in2 => \N__15716\,
            in3 => \N__13847\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_2\,
            carryout => \un1_M_this_data_count_q_cry_3\,
            clk => \N__21595\,
            ce => 'H',
            sr => \N__15482\
        );

    \M_this_data_count_q_4_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15557\,
            in2 => \N__20049\,
            in3 => \N__13844\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_3\,
            carryout => \un1_M_this_data_count_q_cry_4\,
            clk => \N__21595\,
            ce => 'H',
            sr => \N__15482\
        );

    \M_this_data_count_q_5_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20019\,
            in2 => \N__15590\,
            in3 => \N__13841\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_4\,
            carryout => \un1_M_this_data_count_q_cry_5\,
            clk => \N__21595\,
            ce => 'H',
            sr => \N__15482\
        );

    \M_this_data_count_q_6_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15602\,
            in2 => \N__20050\,
            in3 => \N__13838\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_5\,
            carryout => \un1_M_this_data_count_q_cry_6\,
            clk => \N__21595\,
            ce => 'H',
            sr => \N__15482\
        );

    \M_this_data_count_q_7_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20023\,
            in2 => \N__15575\,
            in3 => \N__13835\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_6\,
            carryout => \un1_M_this_data_count_q_cry_7\,
            clk => \N__21595\,
            ce => 'H',
            sr => \N__15482\
        );

    \M_this_data_count_q_8_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15527\,
            in2 => \N__20051\,
            in3 => \N__13832\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_24_0_\,
            carryout => \un1_M_this_data_count_q_cry_8\,
            clk => \N__21604\,
            ce => 'H',
            sr => \N__15478\
        );

    \M_this_data_count_q_9_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15500\,
            in2 => \N__20054\,
            in3 => \N__13829\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_8\,
            carryout => \un1_M_this_data_count_q_cry_9\,
            clk => \N__21604\,
            ce => 'H',
            sr => \N__15478\
        );

    \M_this_data_count_q_10_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15539\,
            in2 => \N__20052\,
            in3 => \N__13826\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_9\,
            carryout => \un1_M_this_data_count_q_cry_10\,
            clk => \N__21604\,
            ce => 'H',
            sr => \N__15478\
        );

    \M_this_data_count_q_11_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15514\,
            in2 => \N__20055\,
            in3 => \N__13823\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_10\,
            carryout => \un1_M_this_data_count_q_cry_11\,
            clk => \N__21604\,
            ce => 'H',
            sr => \N__15478\
        );

    \M_this_data_count_q_12_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15685\,
            in2 => \N__20053\,
            in3 => \N__13820\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_11\,
            carryout => \un1_M_this_data_count_q_cry_12\,
            clk => \N__21604\,
            ce => 'H',
            sr => \N__15478\
        );

    \un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20131\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_12\,
            carryout => \un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__20181\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO\,
            carryout => \un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20135\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO\,
            carryout => \un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21761\,
            in1 => \N__20040\,
            in2 => \N__15659\,
            in3 => \N__14822\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21614\,
            ce => 'H',
            sr => \N__21340\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_1_c2_1_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101101111000"
        )
    port map (
            in0 => \N__14259\,
            in1 => \N__14118\,
            in2 => \N__14482\,
            in3 => \N__14609\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_1_c2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_1_c2_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100000101"
        )
    port map (
            in0 => \N__14610\,
            in1 => \_gnd_net_\,
            in2 => \N__14819\,
            in3 => \N__14812\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_1_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum1_i_1_3_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001000101011"
        )
    port map (
            in0 => \N__14627\,
            in1 => \N__14119\,
            in2 => \N__14618\,
            in3 => \N__14611\,
            lcout => \this_vga_signals.mult1_un54_sum1_i_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_address_buffer_q_esr_5_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001001001101"
        )
    port map (
            in0 => \N__14477\,
            in1 => \N__14297\,
            in2 => \N__14126\,
            in3 => \N__13961\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21583\,
            ce => \N__15317\,
            sr => \N__15211\
        );

    \this_vga_signals.M_address_buffer_q_esr_13_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100100"
        )
    port map (
            in0 => \N__15446\,
            in1 => \N__15410\,
            in2 => \N__15392\,
            in3 => \N__15344\,
            lcout => \M_this_vga_signals_address_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21584\,
            ce => \N__15316\,
            sr => \N__15215\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15098\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21589\,
            ce => \N__15011\,
            sr => \N__14958\
        );

    \this_start_data_delay.M_last_q_RNI9P6N1_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__15978\,
            in1 => \N__21395\,
            in2 => \N__15740\,
            in3 => \N__19023\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_state_q_srsts_i_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_2_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001110000"
        )
    port map (
            in0 => \N__15620\,
            in1 => \N__15979\,
            in2 => \N__14900\,
            in3 => \N__18771\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_1_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001001111"
        )
    port map (
            in0 => \N__15616\,
            in1 => \N__15739\,
            in2 => \N__14897\,
            in3 => \N__21389\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_i_a2_0_1_1_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__21747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19996\,
            lcout => \this_start_data_delay.N_389_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.dma_i_a2_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19995\,
            in1 => \N__15975\,
            in2 => \_gnd_net_\,
            in3 => \N__19014\,
            lcout => port_dmab_c,
            ltout => \port_dmab_c_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI7S6U1_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21746\,
            in1 => \N__21387\,
            in2 => \N__14828\,
            in3 => \N__18740\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNINC2J4_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__21388\,
            in1 => \N__15976\,
            in2 => \N__14825\,
            in3 => \N__15615\,
            lcout => \this_start_data_delay.M_this_state_q_srsts_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_i_a2_1_9_1_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15712\,
            in1 => \N__15697\,
            in2 => \N__15686\,
            in3 => \N__15670\,
            lcout => \this_start_data_delay.M_this_state_q_srsts_i_a2_1_9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_i_a2_1_6_1_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15658\,
            in2 => \_gnd_net_\,
            in3 => \N__15640\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_state_q_srsts_i_a2_1_6Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_i_a2_1_1_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15629\,
            in1 => \N__15545\,
            in2 => \N__15623\,
            in3 => \N__15488\,
            lcout => \this_start_data_delay.N_413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_i_a2_1_8_1_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15601\,
            in1 => \N__15586\,
            in2 => \N__15574\,
            in3 => \N__15556\,
            lcout => \this_start_data_delay.M_this_state_q_srsts_i_a2_1_8Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_i_a2_1_7_1_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15538\,
            in1 => \N__15526\,
            in2 => \N__15515\,
            in3 => \N__15499\,
            lcout => \this_start_data_delay.M_this_state_q_srsts_i_a2_1_7Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI20CE_0_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21393\,
            lcout => \M_this_state_q_RNI20CEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15798\,
            in2 => \_gnd_net_\,
            in3 => \N__15776\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__15799\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15464\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15800\,
            in2 => \_gnd_net_\,
            in3 => \N__15806\,
            lcout => \M_this_state_q_nss_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15797\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_0_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15766\,
            lcout => \M_this_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_11_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__15722\,
            in1 => \N__21782\,
            in2 => \N__18051\,
            in3 => \N__17471\,
            lcout => \M_this_internal_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21601\,
            ce => 'H',
            sr => \N__21342\
        );

    \this_start_data_delay.M_this_state_q_srsts_0_a2_1_0_4_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__15946\,
            in1 => \N__21394\,
            in2 => \N__20039\,
            in3 => \N__19015\,
            lcout => \this_start_data_delay.M_this_state_q_srsts_0_a2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15749\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI8LQ11_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__15853\,
            in1 => \N__15876\,
            in2 => \N__15839\,
            in3 => \N__15977\,
            lcout => \this_start_data_delay.N_353_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBJQQ_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__15877\,
            in1 => \N__15834\,
            in2 => \_gnd_net_\,
            in3 => \N__15851\,
            lcout => \M_this_start_data_delay_out_0\,
            ltout => \M_this_start_data_delay_out_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_11_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001111111"
        )
    port map (
            in0 => \N__18938\,
            in1 => \N__17737\,
            in2 => \N__15725\,
            in3 => \N__20634\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNICHCU_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__15878\,
            in1 => \N__15835\,
            in2 => \N__15920\,
            in3 => \N__15852\,
            lcout => \this_start_data_delay.N_352_0\,
            ltout => \this_start_data_delay.N_352_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011111111"
        )
    port map (
            in0 => \N__16073\,
            in1 => \N__15896\,
            in2 => \N__15890\,
            in3 => \N__15887\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__15875\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15854\,
            lcout => \this_start_data_delay.M_last_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIILOC1_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__15824\,
            in1 => \N__15945\,
            in2 => \_gnd_net_\,
            in3 => \N__21391\,
            lcout => \this_start_data_delay.N_398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_4_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011101010101"
        )
    port map (
            in0 => \N__16896\,
            in1 => \N__17722\,
            in2 => \N__18937\,
            in3 => \N__18761\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_1_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011011111"
        )
    port map (
            in0 => \N__18791\,
            in1 => \N__17721\,
            in2 => \N__18270\,
            in3 => \N__16290\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIHI621_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21392\,
            in2 => \_gnd_net_\,
            in3 => \N__18790\,
            lcout => \this_start_data_delay.N_407\,
            ltout => \this_start_data_delay.N_407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_6_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__16001\,
            in1 => \N__15995\,
            in2 => \N__15818\,
            in3 => \N__16092\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21619\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_1_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001110100001100"
        )
    port map (
            in0 => \N__21718\,
            in1 => \N__18013\,
            in2 => \N__15815\,
            in3 => \N__16271\,
            lcout => \M_this_internal_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21624\,
            ce => 'H',
            sr => \N__21341\
        );

    \this_start_data_delay.M_this_internal_address_q_3s2_LC_18_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__15994\,
            in1 => \N__17726\,
            in2 => \_gnd_net_\,
            in3 => \N__21717\,
            lcout => \M_this_internal_address_q_3_sm0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_5_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011011111"
        )
    port map (
            in0 => \N__18793\,
            in1 => \N__17746\,
            in2 => \N__18226\,
            in3 => \N__16765\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_7_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__17748\,
            in1 => \N__16632\,
            in2 => \N__18980\,
            in3 => \N__18794\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_3_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100110011"
        )
    port map (
            in0 => \N__17747\,
            in1 => \N__17035\,
            in2 => \N__19520\,
            in3 => \N__18792\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_13_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__17734\,
            in1 => \N__20550\,
            in2 => \N__20942\,
            in3 => \N__18738\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_12_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__17735\,
            in1 => \N__20730\,
            in2 => \N__18227\,
            in3 => \N__18737\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI95RM1_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__15983\,
            in1 => \N__18683\,
            in2 => \N__15947\,
            in3 => \N__18736\,
            lcout => \N_346_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_9_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__17736\,
            in1 => \N__16497\,
            in2 => \N__20977\,
            in3 => \N__18739\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_4_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010100110000"
        )
    port map (
            in0 => \N__21836\,
            in1 => \N__15926\,
            in2 => \N__18082\,
            in3 => \N__16877\,
            lcout => \M_this_internal_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21616\,
            ce => 'H',
            sr => \N__21343\
        );

    \M_this_internal_address_q_2_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100110000"
        )
    port map (
            in0 => \N__16112\,
            in1 => \N__21838\,
            in2 => \N__16133\,
            in3 => \N__18069\,
            lcout => \M_this_internal_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21616\,
            ce => 'H',
            sr => \N__21343\
        );

    \M_this_internal_address_q_9_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010100110000"
        )
    port map (
            in0 => \N__21837\,
            in1 => \N__16118\,
            in2 => \N__18083\,
            in3 => \N__16478\,
            lcout => \M_this_internal_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21616\,
            ce => 'H',
            sr => \N__21343\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_10_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__17719\,
            in1 => \N__17196\,
            in2 => \N__19519\,
            in3 => \N__18762\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_2_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100110011"
        )
    port map (
            in0 => \N__17720\,
            in1 => \N__16152\,
            in2 => \N__20984\,
            in3 => \N__18763\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_5_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__16061\,
            in1 => \N__16105\,
            in2 => \N__17745\,
            in3 => \N__16093\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__16106\,
            in1 => \N__16094\,
            in2 => \N__19053\,
            in3 => \N__16079\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_d29_LC_19_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17491\,
            in1 => \N__16023\,
            in2 => \N__16055\,
            in3 => \N__21201\,
            lcout => \this_start_data_delay.M_this_state_dZ0Z29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_0_a2_3_4_LC_19_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111111111111"
        )
    port map (
            in0 => \N__16053\,
            in1 => \N__16025\,
            in2 => \N__21206\,
            in3 => \N__17492\,
            lcout => \this_start_data_delay.N_396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_d27_LC_19_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__17489\,
            in1 => \N__16022\,
            in2 => \N__16054\,
            in3 => \N__21197\,
            lcout => \this_start_data_delay.M_this_state_dZ0Z27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_d28_LC_19_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16052\,
            in1 => \N__16024\,
            in2 => \N__21205\,
            in3 => \N__17490\,
            lcout => \this_start_data_delay.M_this_state_dZ0Z28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_13_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16466\,
            lcout => \this_vram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_12_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16457\,
            lcout => \this_vram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_5_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__16445\,
            in1 => \N__21857\,
            in2 => \N__18073\,
            in3 => \N__16745\,
            lcout => \M_this_internal_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => 'H',
            sr => \N__21346\
        );

    \M_this_internal_address_q_3_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101010000"
        )
    port map (
            in0 => \N__21856\,
            in1 => \N__16439\,
            in2 => \N__17012\,
            in3 => \N__18046\,
            lcout => \M_this_internal_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => 'H',
            sr => \N__21346\
        );

    \M_this_internal_address_q_7_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__18045\,
            in1 => \N__21858\,
            in2 => \N__16433\,
            in3 => \N__16613\,
            lcout => \M_this_internal_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => 'H',
            sr => \N__21346\
        );

    \M_this_internal_address_q_0_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101000100"
        )
    port map (
            in0 => \N__21855\,
            in1 => \N__16406\,
            in2 => \N__17324\,
            in3 => \N__18050\,
            lcout => \M_this_internal_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21609\,
            ce => 'H',
            sr => \N__21346\
        );

    \M_this_internal_address_q_RNI6EA12_0_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17343\,
            in2 => \N__16421\,
            in3 => \N__16420\,
            lcout => \M_this_internal_address_q_RNI6EA12Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_20_21_0_\,
            carryout => \un1_M_this_internal_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_0_c_RNI4MQI_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16303\,
            in2 => \_gnd_net_\,
            in3 => \N__16259\,
            lcout => \un1_M_this_internal_address_q_cry_0_c_RNI4MQIZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_0\,
            carryout => \un1_M_this_internal_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_1_c_RNI6PRI_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16153\,
            in2 => \_gnd_net_\,
            in3 => \N__16121\,
            lcout => \un1_M_this_internal_address_q_cry_1_c_RNI6PRIZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_1\,
            carryout => \un1_M_this_internal_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_2_c_RNI8SSI_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17031\,
            in2 => \_gnd_net_\,
            in3 => \N__17003\,
            lcout => \un1_M_this_internal_address_q_cry_2_c_RNI8SSIZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_2\,
            carryout => \un1_M_this_internal_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_3_c_RNIAVTI_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16897\,
            in2 => \_gnd_net_\,
            in3 => \N__16871\,
            lcout => \un1_M_this_internal_address_q_cry_3_c_RNIAVTIZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_3\,
            carryout => \un1_M_this_internal_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_4_c_RNIC2VI_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16764\,
            in2 => \_gnd_net_\,
            in3 => \N__16739\,
            lcout => \un1_M_this_internal_address_q_cry_4_c_RNIC2VIZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_4\,
            carryout => \un1_M_this_internal_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_5_c_RNIE50J_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17775\,
            in2 => \_gnd_net_\,
            in3 => \N__16736\,
            lcout => \un1_M_this_internal_address_q_cry_5_c_RNIE50JZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_5\,
            carryout => \un1_M_this_internal_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_6_c_RNIG81J_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16633\,
            in2 => \_gnd_net_\,
            in3 => \N__16607\,
            lcout => \un1_M_this_internal_address_q_cry_6_c_RNIG81JZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_6\,
            carryout => \un1_M_this_internal_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_7_c_RNIIB2J_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17539\,
            in2 => \_gnd_net_\,
            in3 => \N__16604\,
            lcout => \un1_M_this_internal_address_q_cry_7_c_RNIIB2JZ0\,
            ltout => OPEN,
            carryin => \bfn_20_22_0_\,
            carryout => \un1_M_this_internal_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_8_c_RNIKE3J_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16498\,
            in2 => \_gnd_net_\,
            in3 => \N__16472\,
            lcout => \un1_M_this_internal_address_q_cry_8_c_RNIKE3JZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_8\,
            carryout => \un1_M_this_internal_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_9_c_RNITQCI_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17197\,
            in2 => \_gnd_net_\,
            in3 => \N__16469\,
            lcout => \un1_M_this_internal_address_q_cry_9_c_RNITQCIZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_9\,
            carryout => \un1_M_this_internal_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_10_c_RNI6I0D_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20663\,
            in2 => \_gnd_net_\,
            in3 => \N__17459\,
            lcout => \un1_M_this_internal_address_q_cry_10_c_RNI6I0DZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_10\,
            carryout => \un1_M_this_internal_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_11_c_RNI8L1D_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20712\,
            in2 => \_gnd_net_\,
            in3 => \N__17456\,
            lcout => \un1_M_this_internal_address_q_cry_11_c_RNI8L1DZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_11\,
            carryout => \un1_M_this_internal_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_internal_address_q_cry_12_c_RNIAO2D_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20526\,
            in2 => \_gnd_net_\,
            in3 => \N__17453\,
            lcout => \un1_M_this_internal_address_q_cry_12_c_RNIAO2DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_0_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001111"
        )
    port map (
            in0 => \N__17741\,
            in1 => \N__18975\,
            in2 => \N__17356\,
            in3 => \N__18783\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_10_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__17312\,
            in1 => \N__21835\,
            in2 => \N__18080\,
            in3 => \N__17306\,
            lcout => \M_this_internal_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21626\,
            ce => 'H',
            sr => \N__21344\
        );

    \M_this_internal_address_q_12_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__17177\,
            in1 => \N__21859\,
            in2 => \N__18085\,
            in3 => \N__17168\,
            lcout => \M_this_internal_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21620\,
            ce => 'H',
            sr => \N__21347\
        );

    \M_this_internal_address_q_6_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__17756\,
            in1 => \N__21860\,
            in2 => \N__18086\,
            in3 => \N__17162\,
            lcout => \M_this_internal_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21620\,
            ce => 'H',
            sr => \N__21347\
        );

    \M_this_internal_address_q_13_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__17156\,
            in1 => \N__21820\,
            in2 => \N__18081\,
            in3 => \N__17144\,
            lcout => \M_this_internal_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21627\,
            ce => 'H',
            sr => \N__21345\
        );

    \M_this_internal_address_q_8_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010011110100"
        )
    port map (
            in0 => \N__21819\,
            in1 => \N__17138\,
            in2 => \N__18084\,
            in3 => \N__17519\,
            lcout => \M_this_internal_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21627\,
            ce => 'H',
            sr => \N__21345\
        );

    \M_this_state_q_3_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19030\,
            in2 => \_gnd_net_\,
            in3 => \N__18798\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21627\,
            ce => 'H',
            sr => \N__21345\
        );

    \this_vram.mem_mem_0_0_RNIQOI11_0_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19618\,
            in1 => \N__17972\,
            in2 => \_gnd_net_\,
            in3 => \N__17963\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI95PB2_11_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__18363\,
            in1 => \N__19212\,
            in2 => \N__17948\,
            in3 => \N__18512\,
            lcout => \this_vram.mem_DOUT_7_i_m2_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_11_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17945\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIDSEJ4_11_LC_22_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__19775\,
            in1 => \N__18473\,
            in2 => \N__18365\,
            in3 => \N__17936\,
            lcout => \M_this_vram_read_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_6_LC_22_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100110011"
        )
    port map (
            in0 => \N__17749\,
            in1 => \N__17776\,
            in2 => \N__20938\,
            in3 => \N__18800\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.M_this_internal_address_q_3_ns_1_8_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__17750\,
            in1 => \N__17538\,
            in2 => \N__18278\,
            in3 => \N__18797\,
            lcout => \this_vram.M_this_internal_address_q_3_ns_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_d27_2_LC_22_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__17513\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17501\,
            lcout => \this_start_data_delay.M_this_state_d27Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_wclke_3_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20759\,
            in1 => \N__20685\,
            in2 => \N__20595\,
            in3 => \N__20502\,
            lcout => \this_vram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_RNIU0N11_0_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19619\,
            in1 => \N__18542\,
            in2 => \_gnd_net_\,
            in3 => \N__18527\,
            lcout => \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_RNI05P11_0_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18506\,
            in1 => \N__18488\,
            in2 => \_gnd_net_\,
            in3 => \N__19628\,
            lcout => \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIKREJ4_11_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18351\,
            in1 => \N__19160\,
            in2 => \_gnd_net_\,
            in3 => \N__19277\,
            lcout => \M_this_vram_read_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI95PB2_0_11_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__19211\,
            in1 => \N__19097\,
            in2 => \N__19133\,
            in3 => \N__18350\,
            lcout => \this_vram.mem_DOUT_7_i_m2_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNID5PB2_11_LC_23_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__19199\,
            in1 => \N__19340\,
            in2 => \N__19637\,
            in3 => \N__18355\,
            lcout => OPEN,
            ltout => \this_vram.mem_DOUT_7_i_m2_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNILSEJ4_11_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__18359\,
            in1 => \N__19706\,
            in2 => \N__18422\,
            in3 => \N__19739\,
            lcout => \M_this_vram_read_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIDSEJ4_0_11_LC_23_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__19670\,
            in1 => \N__19526\,
            in2 => \N__18364\,
            in3 => \N__18323\,
            lcout => \M_this_vram_read_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIIUD53_LC_23_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__18274\,
            in1 => \N__20901\,
            in2 => \N__18219\,
            in3 => \N__20879\,
            lcout => \M_this_vram_write_data_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un23_i_o2_LC_23_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19054\,
            in2 => \_gnd_net_\,
            in3 => \N__19019\,
            lcout => \this_start_data_delay.N_351_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIDVQ81_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__19055\,
            in1 => \N__19965\,
            in2 => \_gnd_net_\,
            in3 => \N__18799\,
            lcout => \this_start_data_delay.un1_M_this_state_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI9MQ11_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19031\,
            in2 => \_gnd_net_\,
            in3 => \N__18795\,
            lcout => \M_this_vram_write_data_0_sqmuxa\,
            ltout => \M_this_vram_write_data_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIGSD53_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__18979\,
            in1 => \N__18933\,
            in2 => \N__18890\,
            in3 => \N__20876\,
            lcout => \M_this_vram_write_data_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIB2RF1_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__18796\,
            in1 => \N__19943\,
            in2 => \_gnd_net_\,
            in3 => \N__18682\,
            lcout => \M_this_vram_write_en_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_wclke_3_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__20762\,
            in1 => \N__20681\,
            in2 => \N__20597\,
            in3 => \N__20513\,
            lcout => \this_vram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_wclke_3_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__20760\,
            in1 => \N__20680\,
            in2 => \N__20596\,
            in3 => \N__20511\,
            lcout => \this_vram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_wclke_3_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__20512\,
            in1 => \N__20590\,
            in2 => \N__20687\,
            in3 => \N__20761\,
            lcout => \this_vram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_1_RNISOI11_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19622\,
            in1 => \N__18602\,
            in2 => \_gnd_net_\,
            in3 => \N__18590\,
            lcout => \this_vram.mem_mem_0_1_RNISOIZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_1_RNI7JS51_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__19616\,
            in1 => \N__19331\,
            in2 => \N__19213\,
            in3 => \N__19319\,
            lcout => OPEN,
            ltout => \this_vram.mem_DOUT_6_i_m2_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_1_RNI8NL72_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__19304\,
            in1 => \N__19295\,
            in2 => \N__19280\,
            in3 => \N__19209\,
            lcout => \this_vram.mem_N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_1_RNI5FQ51_LC_24_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__19617\,
            in1 => \N__19271\,
            in2 => \N__19214\,
            in3 => \N__19259\,
            lcout => OPEN,
            ltout => \this_vram.mem_DOUT_3_i_m2_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_1_RNI4FH72_LC_24_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__19244\,
            in1 => \N__19229\,
            in2 => \N__19217\,
            in3 => \N__19210\,
            lcout => \this_vram.mem_N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_RNIQOI11_LC_24_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19154\,
            in1 => \N__19615\,
            in2 => \_gnd_net_\,
            in3 => \N__19139\,
            lcout => \this_vram.mem_mem_0_0_RNIQOIZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_RNIU0N11_LC_24_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19620\,
            in1 => \N__19124\,
            in2 => \_gnd_net_\,
            in3 => \N__19112\,
            lcout => \this_vram.mem_mem_2_0_RNIU0NZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_0_wclke_3_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__20679\,
            in1 => \N__20751\,
            in2 => \N__20594\,
            in3 => \N__20510\,
            lcout => \this_vram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19070\,
            in1 => \N__19784\,
            in2 => \_gnd_net_\,
            in3 => \N__19621\,
            lcout => \this_vram.mem_mem_1_0_RNISSK11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_1_RNIUSK11_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19626\,
            in1 => \N__19766\,
            in2 => \_gnd_net_\,
            in3 => \N__19754\,
            lcout => \this_vram.mem_mem_1_1_RNIUSKZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_1_RNI25P11_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19627\,
            in1 => \N__19733\,
            in2 => \_gnd_net_\,
            in3 => \N__19718\,
            lcout => \this_vram.mem_mem_3_1_RNI25PZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_RNI05P11_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19700\,
            in1 => \N__19685\,
            in2 => \_gnd_net_\,
            in3 => \N__19625\,
            lcout => \this_vram.mem_mem_3_0_RNI05PZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_1_RNI01N11_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__19664\,
            in1 => \_gnd_net_\,
            in2 => \N__19652\,
            in3 => \N__19623\,
            lcout => \this_vram.mem_mem_2_1_RNI01NZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_RNISSK11_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19624\,
            in1 => \N__19553\,
            in2 => \_gnd_net_\,
            in3 => \N__19544\,
            lcout => \this_vram.mem_mem_1_0_RNISSKZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIM2E53_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__19506\,
            in1 => \N__20878\,
            in2 => \N__19463\,
            in3 => \N__20902\,
            lcout => \M_this_vram_write_data_0_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_5_0_wclke_3_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20734\,
            in1 => \N__20567\,
            in2 => \N__20664\,
            in3 => \N__20489\,
            lcout => \this_vram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIK0E53_LC_24_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__20970\,
            in1 => \N__20920\,
            in2 => \N__20903\,
            in3 => \N__20877\,
            lcout => \M_this_vram_write_data_0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_7_0_wclke_3_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__20488\,
            in1 => \N__20554\,
            in2 => \N__20686\,
            in3 => \N__20750\,
            lcout => \this_vram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_6_0_wclke_3_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20749\,
            in1 => \N__20675\,
            in2 => \N__20566\,
            in3 => \N__20487\,
            lcout => \this_vram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_24_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_0_LC_30_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21843\,
            in1 => \N__19888\,
            in2 => \N__20060\,
            in3 => \N__20059\,
            lcout => \M_this_external_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_30_23_0_\,
            carryout => \un1_M_this_external_address_q_cry_0\,
            clk => \N__21648\,
            ce => 'H',
            sr => \N__21350\
        );

    \M_this_external_address_q_1_LC_30_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21851\,
            in1 => \N__19867\,
            in2 => \_gnd_net_\,
            in3 => \N__19856\,
            lcout => \M_this_external_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_0\,
            carryout => \un1_M_this_external_address_q_cry_1\,
            clk => \N__21648\,
            ce => 'H',
            sr => \N__21350\
        );

    \M_this_external_address_q_2_LC_30_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21844\,
            in1 => \N__19837\,
            in2 => \_gnd_net_\,
            in3 => \N__19826\,
            lcout => \M_this_external_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_1\,
            carryout => \un1_M_this_external_address_q_cry_2\,
            clk => \N__21648\,
            ce => 'H',
            sr => \N__21350\
        );

    \M_this_external_address_q_3_LC_30_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21852\,
            in1 => \N__19813\,
            in2 => \_gnd_net_\,
            in3 => \N__19802\,
            lcout => \M_this_external_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_2\,
            carryout => \un1_M_this_external_address_q_cry_3\,
            clk => \N__21648\,
            ce => 'H',
            sr => \N__21350\
        );

    \M_this_external_address_q_4_LC_30_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21845\,
            in1 => \N__19795\,
            in2 => \_gnd_net_\,
            in3 => \N__21176\,
            lcout => \M_this_external_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_3\,
            carryout => \un1_M_this_external_address_q_cry_4\,
            clk => \N__21648\,
            ce => 'H',
            sr => \N__21350\
        );

    \M_this_external_address_q_5_LC_30_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21853\,
            in1 => \N__21166\,
            in2 => \_gnd_net_\,
            in3 => \N__21155\,
            lcout => \M_this_external_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_4\,
            carryout => \un1_M_this_external_address_q_cry_5\,
            clk => \N__21648\,
            ce => 'H',
            sr => \N__21350\
        );

    \M_this_external_address_q_6_LC_30_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21846\,
            in1 => \N__21145\,
            in2 => \_gnd_net_\,
            in3 => \N__21134\,
            lcout => \M_this_external_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_5\,
            carryout => \un1_M_this_external_address_q_cry_6\,
            clk => \N__21648\,
            ce => 'H',
            sr => \N__21350\
        );

    \M_this_external_address_q_7_LC_30_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21854\,
            in1 => \N__21118\,
            in2 => \_gnd_net_\,
            in3 => \N__21107\,
            lcout => \M_this_external_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_6\,
            carryout => \un1_M_this_external_address_q_cry_7\,
            clk => \N__21648\,
            ce => 'H',
            sr => \N__21350\
        );

    \M_this_external_address_q_8_LC_30_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21850\,
            in1 => \N__21085\,
            in2 => \_gnd_net_\,
            in3 => \N__21074\,
            lcout => \M_this_external_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_30_24_0_\,
            carryout => \un1_M_this_external_address_q_cry_8\,
            clk => \N__21651\,
            ce => 'H',
            sr => \N__21348\
        );

    \M_this_external_address_q_9_LC_30_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21841\,
            in1 => \N__21064\,
            in2 => \_gnd_net_\,
            in3 => \N__21053\,
            lcout => \M_this_external_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_8\,
            carryout => \un1_M_this_external_address_q_cry_9\,
            clk => \N__21651\,
            ce => 'H',
            sr => \N__21348\
        );

    \M_this_external_address_q_10_LC_30_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21847\,
            in1 => \N__21034\,
            in2 => \_gnd_net_\,
            in3 => \N__21023\,
            lcout => \M_this_external_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_9\,
            carryout => \un1_M_this_external_address_q_cry_10\,
            clk => \N__21651\,
            ce => 'H',
            sr => \N__21348\
        );

    \M_this_external_address_q_11_LC_30_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21839\,
            in1 => \N__21016\,
            in2 => \_gnd_net_\,
            in3 => \N__21005\,
            lcout => \M_this_external_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_10\,
            carryout => \un1_M_this_external_address_q_cry_11\,
            clk => \N__21651\,
            ce => 'H',
            sr => \N__21348\
        );

    \M_this_external_address_q_12_LC_30_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21848\,
            in1 => \N__20998\,
            in2 => \_gnd_net_\,
            in3 => \N__20987\,
            lcout => \M_this_external_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_11\,
            carryout => \un1_M_this_external_address_q_cry_12\,
            clk => \N__21651\,
            ce => 'H',
            sr => \N__21348\
        );

    \M_this_external_address_q_13_LC_30_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__21840\,
            in1 => \N__21898\,
            in2 => \_gnd_net_\,
            in3 => \N__21887\,
            lcout => \M_this_external_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_12\,
            carryout => \un1_M_this_external_address_q_cry_13\,
            clk => \N__21651\,
            ce => 'H',
            sr => \N__21348\
        );

    \M_this_external_address_q_14_LC_30_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21849\,
            in1 => \N__21874\,
            in2 => \_gnd_net_\,
            in3 => \N__21863\,
            lcout => \M_this_external_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_13\,
            carryout => \un1_M_this_external_address_q_cry_14\,
            clk => \N__21651\,
            ce => 'H',
            sr => \N__21348\
        );

    \M_this_external_address_q_15_LC_30_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__21842\,
            in1 => \N__21664\,
            in2 => \_gnd_net_\,
            in3 => \N__21680\,
            lcout => \M_this_external_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21651\,
            ce => 'H',
            sr => \N__21348\
        );

    \this_start_data_delay.M_this_state_d27_6_LC_32_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21266\,
            in1 => \N__21254\,
            in2 => \N__21242\,
            in3 => \N__21218\,
            lcout => \this_start_data_delay.M_this_state_d27Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
