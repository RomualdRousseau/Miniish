// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 3 2022 11:35:56

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    rgb,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    debug,
    clk);

    input [15:0] port_address;
    input [7:0] port_data;
    output [5:0] rgb;
    output vsync;
    output vblank;
    input rst_n;
    input port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    output debug;
    input clk;

    wire N__20690;
    wire N__20689;
    wire N__20688;
    wire N__20679;
    wire N__20678;
    wire N__20677;
    wire N__20670;
    wire N__20669;
    wire N__20668;
    wire N__20661;
    wire N__20660;
    wire N__20659;
    wire N__20652;
    wire N__20651;
    wire N__20650;
    wire N__20643;
    wire N__20642;
    wire N__20641;
    wire N__20634;
    wire N__20633;
    wire N__20632;
    wire N__20625;
    wire N__20624;
    wire N__20623;
    wire N__20616;
    wire N__20615;
    wire N__20614;
    wire N__20607;
    wire N__20606;
    wire N__20605;
    wire N__20598;
    wire N__20597;
    wire N__20596;
    wire N__20589;
    wire N__20588;
    wire N__20587;
    wire N__20580;
    wire N__20579;
    wire N__20578;
    wire N__20571;
    wire N__20570;
    wire N__20569;
    wire N__20562;
    wire N__20561;
    wire N__20560;
    wire N__20553;
    wire N__20552;
    wire N__20551;
    wire N__20544;
    wire N__20543;
    wire N__20542;
    wire N__20535;
    wire N__20534;
    wire N__20533;
    wire N__20526;
    wire N__20525;
    wire N__20524;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20508;
    wire N__20507;
    wire N__20506;
    wire N__20499;
    wire N__20498;
    wire N__20497;
    wire N__20490;
    wire N__20489;
    wire N__20488;
    wire N__20481;
    wire N__20480;
    wire N__20479;
    wire N__20472;
    wire N__20471;
    wire N__20470;
    wire N__20463;
    wire N__20462;
    wire N__20461;
    wire N__20454;
    wire N__20453;
    wire N__20452;
    wire N__20445;
    wire N__20444;
    wire N__20443;
    wire N__20436;
    wire N__20435;
    wire N__20434;
    wire N__20427;
    wire N__20426;
    wire N__20425;
    wire N__20418;
    wire N__20417;
    wire N__20416;
    wire N__20409;
    wire N__20408;
    wire N__20407;
    wire N__20400;
    wire N__20399;
    wire N__20398;
    wire N__20391;
    wire N__20390;
    wire N__20389;
    wire N__20372;
    wire N__20369;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20349;
    wire N__20344;
    wire N__20341;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20329;
    wire N__20328;
    wire N__20327;
    wire N__20326;
    wire N__20321;
    wire N__20320;
    wire N__20319;
    wire N__20318;
    wire N__20317;
    wire N__20314;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20285;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20273;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20228;
    wire N__20225;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20217;
    wire N__20212;
    wire N__20209;
    wire N__20208;
    wire N__20203;
    wire N__20200;
    wire N__20199;
    wire N__20194;
    wire N__20191;
    wire N__20190;
    wire N__20189;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20168;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20020;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20012;
    wire N__20009;
    wire N__20008;
    wire N__20007;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19999;
    wire N__19996;
    wire N__19995;
    wire N__19994;
    wire N__19993;
    wire N__19990;
    wire N__19987;
    wire N__19986;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19890;
    wire N__19887;
    wire N__19884;
    wire N__19877;
    wire N__19874;
    wire N__19865;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19633;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19622;
    wire N__19621;
    wire N__19620;
    wire N__19619;
    wire N__19614;
    wire N__19611;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19593;
    wire N__19590;
    wire N__19585;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19567;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19522;
    wire N__19521;
    wire N__19520;
    wire N__19519;
    wire N__19518;
    wire N__19517;
    wire N__19516;
    wire N__19515;
    wire N__19514;
    wire N__19513;
    wire N__19504;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19486;
    wire N__19475;
    wire N__19474;
    wire N__19473;
    wire N__19472;
    wire N__19471;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19457;
    wire N__19454;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19376;
    wire N__19373;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19349;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19325;
    wire N__19324;
    wire N__19319;
    wire N__19318;
    wire N__19317;
    wire N__19316;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19308;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19286;
    wire N__19279;
    wire N__19274;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19253;
    wire N__19244;
    wire N__19243;
    wire N__19240;
    wire N__19239;
    wire N__19238;
    wire N__19237;
    wire N__19234;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19222;
    wire N__19221;
    wire N__19218;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19204;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19185;
    wire N__19182;
    wire N__19177;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19157;
    wire N__19156;
    wire N__19155;
    wire N__19152;
    wire N__19151;
    wire N__19150;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19112;
    wire N__19107;
    wire N__19104;
    wire N__19097;
    wire N__19094;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19082;
    wire N__19081;
    wire N__19078;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19058;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19035;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19001;
    wire N__18998;
    wire N__18997;
    wire N__18996;
    wire N__18993;
    wire N__18990;
    wire N__18989;
    wire N__18986;
    wire N__18981;
    wire N__18978;
    wire N__18977;
    wire N__18976;
    wire N__18973;
    wire N__18968;
    wire N__18965;
    wire N__18964;
    wire N__18961;
    wire N__18960;
    wire N__18957;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18943;
    wire N__18940;
    wire N__18935;
    wire N__18930;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18691;
    wire N__18690;
    wire N__18689;
    wire N__18688;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18677;
    wire N__18674;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18666;
    wire N__18665;
    wire N__18658;
    wire N__18655;
    wire N__18654;
    wire N__18651;
    wire N__18650;
    wire N__18647;
    wire N__18646;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18634;
    wire N__18633;
    wire N__18628;
    wire N__18625;
    wire N__18624;
    wire N__18623;
    wire N__18622;
    wire N__18619;
    wire N__18614;
    wire N__18611;
    wire N__18610;
    wire N__18609;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18595;
    wire N__18594;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18582;
    wire N__18581;
    wire N__18578;
    wire N__18577;
    wire N__18576;
    wire N__18575;
    wire N__18572;
    wire N__18567;
    wire N__18564;
    wire N__18563;
    wire N__18562;
    wire N__18559;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18541;
    wire N__18538;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18522;
    wire N__18521;
    wire N__18520;
    wire N__18519;
    wire N__18516;
    wire N__18515;
    wire N__18514;
    wire N__18511;
    wire N__18508;
    wire N__18505;
    wire N__18502;
    wire N__18499;
    wire N__18496;
    wire N__18495;
    wire N__18488;
    wire N__18485;
    wire N__18478;
    wire N__18471;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18426;
    wire N__18415;
    wire N__18410;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18392;
    wire N__18389;
    wire N__18384;
    wire N__18375;
    wire N__18362;
    wire N__18361;
    wire N__18358;
    wire N__18357;
    wire N__18356;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18348;
    wire N__18347;
    wire N__18346;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18320;
    wire N__18315;
    wire N__18312;
    wire N__18311;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18301;
    wire N__18294;
    wire N__18289;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18079;
    wire N__18076;
    wire N__18073;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17980;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17951;
    wire N__17948;
    wire N__17947;
    wire N__17944;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17848;
    wire N__17845;
    wire N__17842;
    wire N__17841;
    wire N__17838;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17830;
    wire N__17827;
    wire N__17824;
    wire N__17819;
    wire N__17816;
    wire N__17811;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17799;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17767;
    wire N__17764;
    wire N__17761;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17740;
    wire N__17739;
    wire N__17738;
    wire N__17737;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17727;
    wire N__17724;
    wire N__17721;
    wire N__17716;
    wire N__17713;
    wire N__17712;
    wire N__17711;
    wire N__17710;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17688;
    wire N__17687;
    wire N__17686;
    wire N__17685;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17665;
    wire N__17658;
    wire N__17653;
    wire N__17646;
    wire N__17641;
    wire N__17638;
    wire N__17627;
    wire N__17626;
    wire N__17625;
    wire N__17624;
    wire N__17623;
    wire N__17620;
    wire N__17619;
    wire N__17616;
    wire N__17615;
    wire N__17614;
    wire N__17613;
    wire N__17612;
    wire N__17609;
    wire N__17608;
    wire N__17607;
    wire N__17606;
    wire N__17605;
    wire N__17604;
    wire N__17599;
    wire N__17592;
    wire N__17589;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17570;
    wire N__17569;
    wire N__17568;
    wire N__17567;
    wire N__17562;
    wire N__17557;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17520;
    wire N__17507;
    wire N__17504;
    wire N__17503;
    wire N__17502;
    wire N__17501;
    wire N__17500;
    wire N__17499;
    wire N__17496;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17486;
    wire N__17485;
    wire N__17484;
    wire N__17483;
    wire N__17482;
    wire N__17481;
    wire N__17480;
    wire N__17479;
    wire N__17478;
    wire N__17477;
    wire N__17472;
    wire N__17469;
    wire N__17464;
    wire N__17457;
    wire N__17454;
    wire N__17453;
    wire N__17452;
    wire N__17451;
    wire N__17446;
    wire N__17443;
    wire N__17434;
    wire N__17431;
    wire N__17426;
    wire N__17421;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17407;
    wire N__17404;
    wire N__17401;
    wire N__17396;
    wire N__17393;
    wire N__17378;
    wire N__17377;
    wire N__17376;
    wire N__17375;
    wire N__17374;
    wire N__17373;
    wire N__17372;
    wire N__17371;
    wire N__17370;
    wire N__17369;
    wire N__17368;
    wire N__17367;
    wire N__17366;
    wire N__17365;
    wire N__17364;
    wire N__17363;
    wire N__17362;
    wire N__17361;
    wire N__17360;
    wire N__17359;
    wire N__17358;
    wire N__17357;
    wire N__17356;
    wire N__17355;
    wire N__17354;
    wire N__17353;
    wire N__17352;
    wire N__17351;
    wire N__17350;
    wire N__17349;
    wire N__17348;
    wire N__17347;
    wire N__17346;
    wire N__17345;
    wire N__17344;
    wire N__17343;
    wire N__17342;
    wire N__17341;
    wire N__17340;
    wire N__17339;
    wire N__17338;
    wire N__17337;
    wire N__17336;
    wire N__17335;
    wire N__17334;
    wire N__17333;
    wire N__17332;
    wire N__17331;
    wire N__17330;
    wire N__17329;
    wire N__17328;
    wire N__17327;
    wire N__17326;
    wire N__17325;
    wire N__17324;
    wire N__17323;
    wire N__17322;
    wire N__17321;
    wire N__17320;
    wire N__17319;
    wire N__17318;
    wire N__17317;
    wire N__17316;
    wire N__17315;
    wire N__17314;
    wire N__17313;
    wire N__17312;
    wire N__17311;
    wire N__17310;
    wire N__17309;
    wire N__17308;
    wire N__17307;
    wire N__17306;
    wire N__17305;
    wire N__17304;
    wire N__17303;
    wire N__17302;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17140;
    wire N__17137;
    wire N__17136;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17111;
    wire N__17108;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17100;
    wire N__17095;
    wire N__17092;
    wire N__17091;
    wire N__17086;
    wire N__17083;
    wire N__17082;
    wire N__17077;
    wire N__17074;
    wire N__17073;
    wire N__17072;
    wire N__17067;
    wire N__17064;
    wire N__17063;
    wire N__17060;
    wire N__17055;
    wire N__17052;
    wire N__17049;
    wire N__17044;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17032;
    wire N__17029;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17015;
    wire N__17012;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17000;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16988;
    wire N__16985;
    wire N__16984;
    wire N__16981;
    wire N__16978;
    wire N__16977;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16894;
    wire N__16893;
    wire N__16888;
    wire N__16887;
    wire N__16884;
    wire N__16881;
    wire N__16878;
    wire N__16875;
    wire N__16870;
    wire N__16867;
    wire N__16864;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16834;
    wire N__16831;
    wire N__16830;
    wire N__16827;
    wire N__16824;
    wire N__16821;
    wire N__16818;
    wire N__16815;
    wire N__16810;
    wire N__16807;
    wire N__16804;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16782;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16772;
    wire N__16767;
    wire N__16764;
    wire N__16761;
    wire N__16760;
    wire N__16755;
    wire N__16752;
    wire N__16749;
    wire N__16748;
    wire N__16747;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16732;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16713;
    wire N__16708;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16567;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16546;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16422;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16406;
    wire N__16405;
    wire N__16402;
    wire N__16399;
    wire N__16396;
    wire N__16393;
    wire N__16390;
    wire N__16387;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16344;
    wire N__16343;
    wire N__16342;
    wire N__16341;
    wire N__16340;
    wire N__16339;
    wire N__16338;
    wire N__16337;
    wire N__16336;
    wire N__16335;
    wire N__16334;
    wire N__16333;
    wire N__16332;
    wire N__16327;
    wire N__16322;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16302;
    wire N__16297;
    wire N__16296;
    wire N__16295;
    wire N__16294;
    wire N__16293;
    wire N__16292;
    wire N__16291;
    wire N__16290;
    wire N__16289;
    wire N__16288;
    wire N__16287;
    wire N__16286;
    wire N__16285;
    wire N__16284;
    wire N__16283;
    wire N__16282;
    wire N__16281;
    wire N__16280;
    wire N__16279;
    wire N__16276;
    wire N__16265;
    wire N__16260;
    wire N__16257;
    wire N__16246;
    wire N__16243;
    wire N__16236;
    wire N__16229;
    wire N__16222;
    wire N__16217;
    wire N__16214;
    wire N__16207;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16052;
    wire N__16049;
    wire N__16046;
    wire N__16045;
    wire N__16042;
    wire N__16041;
    wire N__16038;
    wire N__16035;
    wire N__16032;
    wire N__16027;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15913;
    wire N__15910;
    wire N__15909;
    wire N__15906;
    wire N__15903;
    wire N__15900;
    wire N__15895;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15854;
    wire N__15851;
    wire N__15848;
    wire N__15845;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15791;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15731;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15714;
    wire N__15711;
    wire N__15708;
    wire N__15705;
    wire N__15702;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15611;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15599;
    wire N__15596;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15584;
    wire N__15583;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15573;
    wire N__15570;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15511;
    wire N__15510;
    wire N__15509;
    wire N__15508;
    wire N__15507;
    wire N__15506;
    wire N__15505;
    wire N__15504;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15473;
    wire N__15472;
    wire N__15471;
    wire N__15470;
    wire N__15469;
    wire N__15468;
    wire N__15467;
    wire N__15466;
    wire N__15465;
    wire N__15464;
    wire N__15463;
    wire N__15462;
    wire N__15459;
    wire N__15456;
    wire N__15453;
    wire N__15450;
    wire N__15447;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15289;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15161;
    wire N__15160;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15125;
    wire N__15122;
    wire N__15119;
    wire N__15116;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15092;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14950;
    wire N__14949;
    wire N__14946;
    wire N__14943;
    wire N__14940;
    wire N__14937;
    wire N__14934;
    wire N__14929;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14800;
    wire N__14799;
    wire N__14796;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14779;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14752;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14593;
    wire N__14590;
    wire N__14589;
    wire N__14586;
    wire N__14583;
    wire N__14580;
    wire N__14577;
    wire N__14574;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14558;
    wire N__14555;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14473;
    wire N__14470;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14358;
    wire N__14357;
    wire N__14354;
    wire N__14353;
    wire N__14352;
    wire N__14351;
    wire N__14350;
    wire N__14349;
    wire N__14348;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14333;
    wire N__14330;
    wire N__14327;
    wire N__14322;
    wire N__14319;
    wire N__14300;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14289;
    wire N__14288;
    wire N__14287;
    wire N__14286;
    wire N__14285;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14268;
    wire N__14263;
    wire N__14252;
    wire N__14249;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14180;
    wire N__14177;
    wire N__14174;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14131;
    wire N__14126;
    wire N__14123;
    wire N__14122;
    wire N__14119;
    wire N__14116;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14069;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14051;
    wire N__14050;
    wire N__14049;
    wire N__14048;
    wire N__14043;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14033;
    wire N__14030;
    wire N__14025;
    wire N__14022;
    wire N__14017;
    wire N__14012;
    wire N__14009;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13822;
    wire N__13821;
    wire N__13820;
    wire N__13819;
    wire N__13818;
    wire N__13817;
    wire N__13816;
    wire N__13815;
    wire N__13814;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13806;
    wire N__13803;
    wire N__13802;
    wire N__13799;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13785;
    wire N__13784;
    wire N__13781;
    wire N__13778;
    wire N__13777;
    wire N__13776;
    wire N__13775;
    wire N__13774;
    wire N__13773;
    wire N__13772;
    wire N__13771;
    wire N__13770;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13762;
    wire N__13761;
    wire N__13760;
    wire N__13757;
    wire N__13752;
    wire N__13749;
    wire N__13748;
    wire N__13739;
    wire N__13734;
    wire N__13733;
    wire N__13730;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13710;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13698;
    wire N__13695;
    wire N__13690;
    wire N__13687;
    wire N__13682;
    wire N__13677;
    wire N__13674;
    wire N__13671;
    wire N__13666;
    wire N__13657;
    wire N__13654;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13633;
    wire N__13630;
    wire N__13625;
    wire N__13614;
    wire N__13611;
    wire N__13604;
    wire N__13599;
    wire N__13592;
    wire N__13583;
    wire N__13580;
    wire N__13579;
    wire N__13578;
    wire N__13577;
    wire N__13576;
    wire N__13575;
    wire N__13574;
    wire N__13571;
    wire N__13566;
    wire N__13565;
    wire N__13564;
    wire N__13563;
    wire N__13560;
    wire N__13557;
    wire N__13556;
    wire N__13555;
    wire N__13554;
    wire N__13553;
    wire N__13552;
    wire N__13549;
    wire N__13546;
    wire N__13541;
    wire N__13532;
    wire N__13529;
    wire N__13524;
    wire N__13519;
    wire N__13516;
    wire N__13513;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13489;
    wire N__13488;
    wire N__13487;
    wire N__13486;
    wire N__13483;
    wire N__13482;
    wire N__13479;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13471;
    wire N__13470;
    wire N__13467;
    wire N__13466;
    wire N__13465;
    wire N__13464;
    wire N__13463;
    wire N__13458;
    wire N__13455;
    wire N__13454;
    wire N__13453;
    wire N__13452;
    wire N__13451;
    wire N__13450;
    wire N__13449;
    wire N__13448;
    wire N__13447;
    wire N__13444;
    wire N__13441;
    wire N__13438;
    wire N__13433;
    wire N__13430;
    wire N__13425;
    wire N__13422;
    wire N__13419;
    wire N__13414;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13402;
    wire N__13401;
    wire N__13400;
    wire N__13399;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13378;
    wire N__13373;
    wire N__13368;
    wire N__13363;
    wire N__13360;
    wire N__13355;
    wire N__13350;
    wire N__13349;
    wire N__13346;
    wire N__13337;
    wire N__13334;
    wire N__13329;
    wire N__13324;
    wire N__13319;
    wire N__13316;
    wire N__13301;
    wire N__13300;
    wire N__13299;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13288;
    wire N__13287;
    wire N__13284;
    wire N__13283;
    wire N__13282;
    wire N__13281;
    wire N__13280;
    wire N__13279;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13245;
    wire N__13242;
    wire N__13237;
    wire N__13234;
    wire N__13211;
    wire N__13210;
    wire N__13207;
    wire N__13204;
    wire N__13201;
    wire N__13198;
    wire N__13193;
    wire N__13190;
    wire N__13189;
    wire N__13186;
    wire N__13183;
    wire N__13180;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13088;
    wire N__13085;
    wire N__13084;
    wire N__13083;
    wire N__13082;
    wire N__13081;
    wire N__13078;
    wire N__13077;
    wire N__13076;
    wire N__13073;
    wire N__13072;
    wire N__13071;
    wire N__13068;
    wire N__13063;
    wire N__13062;
    wire N__13059;
    wire N__13054;
    wire N__13051;
    wire N__13046;
    wire N__13045;
    wire N__13044;
    wire N__13043;
    wire N__13042;
    wire N__13041;
    wire N__13036;
    wire N__13035;
    wire N__13032;
    wire N__13027;
    wire N__13022;
    wire N__13017;
    wire N__13010;
    wire N__13007;
    wire N__13004;
    wire N__12989;
    wire N__12988;
    wire N__12987;
    wire N__12986;
    wire N__12983;
    wire N__12982;
    wire N__12981;
    wire N__12980;
    wire N__12979;
    wire N__12978;
    wire N__12977;
    wire N__12976;
    wire N__12975;
    wire N__12972;
    wire N__12969;
    wire N__12964;
    wire N__12961;
    wire N__12958;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12950;
    wire N__12949;
    wire N__12946;
    wire N__12945;
    wire N__12942;
    wire N__12933;
    wire N__12930;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12916;
    wire N__12913;
    wire N__12908;
    wire N__12907;
    wire N__12904;
    wire N__12901;
    wire N__12898;
    wire N__12891;
    wire N__12888;
    wire N__12881;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12862;
    wire N__12859;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12832;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12815;
    wire N__12814;
    wire N__12813;
    wire N__12812;
    wire N__12809;
    wire N__12808;
    wire N__12807;
    wire N__12806;
    wire N__12805;
    wire N__12804;
    wire N__12803;
    wire N__12802;
    wire N__12801;
    wire N__12800;
    wire N__12799;
    wire N__12798;
    wire N__12797;
    wire N__12796;
    wire N__12795;
    wire N__12794;
    wire N__12791;
    wire N__12790;
    wire N__12787;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12775;
    wire N__12772;
    wire N__12767;
    wire N__12760;
    wire N__12751;
    wire N__12744;
    wire N__12741;
    wire N__12734;
    wire N__12713;
    wire N__12712;
    wire N__12711;
    wire N__12710;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12676;
    wire N__12675;
    wire N__12674;
    wire N__12673;
    wire N__12672;
    wire N__12671;
    wire N__12668;
    wire N__12667;
    wire N__12664;
    wire N__12663;
    wire N__12662;
    wire N__12661;
    wire N__12660;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12652;
    wire N__12651;
    wire N__12650;
    wire N__12643;
    wire N__12638;
    wire N__12637;
    wire N__12634;
    wire N__12629;
    wire N__12628;
    wire N__12627;
    wire N__12626;
    wire N__12625;
    wire N__12624;
    wire N__12621;
    wire N__12620;
    wire N__12615;
    wire N__12612;
    wire N__12607;
    wire N__12604;
    wire N__12603;
    wire N__12602;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12596;
    wire N__12593;
    wire N__12590;
    wire N__12589;
    wire N__12586;
    wire N__12581;
    wire N__12578;
    wire N__12569;
    wire N__12564;
    wire N__12561;
    wire N__12554;
    wire N__12547;
    wire N__12540;
    wire N__12535;
    wire N__12532;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12484;
    wire N__12483;
    wire N__12482;
    wire N__12481;
    wire N__12478;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12466;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12448;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12356;
    wire N__12353;
    wire N__12350;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12338;
    wire N__12335;
    wire N__12332;
    wire N__12329;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12319;
    wire N__12318;
    wire N__12317;
    wire N__12316;
    wire N__12315;
    wire N__12314;
    wire N__12313;
    wire N__12310;
    wire N__12309;
    wire N__12308;
    wire N__12303;
    wire N__12302;
    wire N__12301;
    wire N__12300;
    wire N__12299;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12289;
    wire N__12284;
    wire N__12281;
    wire N__12276;
    wire N__12273;
    wire N__12266;
    wire N__12261;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12232;
    wire N__12231;
    wire N__12228;
    wire N__12223;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12185;
    wire N__12182;
    wire N__12179;
    wire N__12176;
    wire N__12173;
    wire N__12170;
    wire N__12167;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12038;
    wire N__12035;
    wire N__12034;
    wire N__12033;
    wire N__12032;
    wire N__12031;
    wire N__12030;
    wire N__12029;
    wire N__12026;
    wire N__12025;
    wire N__12024;
    wire N__12023;
    wire N__12022;
    wire N__12021;
    wire N__12018;
    wire N__12017;
    wire N__12014;
    wire N__12013;
    wire N__12012;
    wire N__12009;
    wire N__12004;
    wire N__12001;
    wire N__12000;
    wire N__11997;
    wire N__11996;
    wire N__11995;
    wire N__11994;
    wire N__11993;
    wire N__11990;
    wire N__11989;
    wire N__11986;
    wire N__11983;
    wire N__11978;
    wire N__11973;
    wire N__11970;
    wire N__11965;
    wire N__11960;
    wire N__11955;
    wire N__11954;
    wire N__11953;
    wire N__11950;
    wire N__11943;
    wire N__11940;
    wire N__11935;
    wire N__11930;
    wire N__11925;
    wire N__11916;
    wire N__11913;
    wire N__11910;
    wire N__11901;
    wire N__11896;
    wire N__11893;
    wire N__11882;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11870;
    wire N__11869;
    wire N__11866;
    wire N__11865;
    wire N__11864;
    wire N__11861;
    wire N__11856;
    wire N__11853;
    wire N__11852;
    wire N__11851;
    wire N__11848;
    wire N__11847;
    wire N__11846;
    wire N__11845;
    wire N__11844;
    wire N__11841;
    wire N__11840;
    wire N__11839;
    wire N__11838;
    wire N__11837;
    wire N__11836;
    wire N__11835;
    wire N__11834;
    wire N__11833;
    wire N__11832;
    wire N__11831;
    wire N__11828;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11810;
    wire N__11807;
    wire N__11802;
    wire N__11795;
    wire N__11792;
    wire N__11783;
    wire N__11762;
    wire N__11761;
    wire N__11760;
    wire N__11757;
    wire N__11756;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11748;
    wire N__11747;
    wire N__11744;
    wire N__11743;
    wire N__11742;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11728;
    wire N__11725;
    wire N__11724;
    wire N__11723;
    wire N__11722;
    wire N__11719;
    wire N__11714;
    wire N__11711;
    wire N__11708;
    wire N__11701;
    wire N__11698;
    wire N__11693;
    wire N__11678;
    wire N__11677;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11623;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11615;
    wire N__11614;
    wire N__11613;
    wire N__11612;
    wire N__11611;
    wire N__11608;
    wire N__11603;
    wire N__11600;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11576;
    wire N__11573;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11565;
    wire N__11564;
    wire N__11563;
    wire N__11562;
    wire N__11557;
    wire N__11554;
    wire N__11547;
    wire N__11540;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11525;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11462;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11435;
    wire N__11432;
    wire N__11429;
    wire N__11426;
    wire N__11423;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11394;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11382;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11264;
    wire N__11261;
    wire N__11258;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11047;
    wire N__11046;
    wire N__11043;
    wire N__11038;
    wire N__11035;
    wire N__11030;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11026;
    wire N__11025;
    wire N__11024;
    wire N__11023;
    wire N__11020;
    wire N__11017;
    wire N__11016;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11004;
    wire N__11003;
    wire N__11002;
    wire N__10999;
    wire N__10998;
    wire N__10997;
    wire N__10994;
    wire N__10993;
    wire N__10992;
    wire N__10987;
    wire N__10986;
    wire N__10983;
    wire N__10978;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10959;
    wire N__10956;
    wire N__10951;
    wire N__10948;
    wire N__10943;
    wire N__10922;
    wire N__10921;
    wire N__10918;
    wire N__10917;
    wire N__10914;
    wire N__10913;
    wire N__10910;
    wire N__10905;
    wire N__10904;
    wire N__10903;
    wire N__10900;
    wire N__10895;
    wire N__10890;
    wire N__10887;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10871;
    wire N__10870;
    wire N__10869;
    wire N__10868;
    wire N__10865;
    wire N__10864;
    wire N__10857;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10828;
    wire N__10827;
    wire N__10824;
    wire N__10823;
    wire N__10822;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10814;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10791;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10748;
    wire N__10747;
    wire N__10746;
    wire N__10745;
    wire N__10744;
    wire N__10743;
    wire N__10742;
    wire N__10741;
    wire N__10740;
    wire N__10739;
    wire N__10736;
    wire N__10735;
    wire N__10734;
    wire N__10733;
    wire N__10732;
    wire N__10731;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10704;
    wire N__10701;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10689;
    wire N__10684;
    wire N__10673;
    wire N__10670;
    wire N__10669;
    wire N__10668;
    wire N__10667;
    wire N__10666;
    wire N__10665;
    wire N__10664;
    wire N__10661;
    wire N__10648;
    wire N__10645;
    wire N__10638;
    wire N__10633;
    wire N__10630;
    wire N__10619;
    wire N__10616;
    wire N__10615;
    wire N__10612;
    wire N__10609;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10591;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10570;
    wire N__10569;
    wire N__10568;
    wire N__10567;
    wire N__10562;
    wire N__10557;
    wire N__10554;
    wire N__10547;
    wire N__10546;
    wire N__10545;
    wire N__10540;
    wire N__10539;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10531;
    wire N__10528;
    wire N__10523;
    wire N__10522;
    wire N__10521;
    wire N__10520;
    wire N__10519;
    wire N__10518;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10494;
    wire N__10491;
    wire N__10488;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10339;
    wire N__10336;
    wire N__10335;
    wire N__10334;
    wire N__10333;
    wire N__10330;
    wire N__10327;
    wire N__10320;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10306;
    wire N__10303;
    wire N__10300;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10243;
    wire N__10242;
    wire N__10241;
    wire N__10240;
    wire N__10239;
    wire N__10236;
    wire N__10235;
    wire N__10234;
    wire N__10231;
    wire N__10226;
    wire N__10225;
    wire N__10224;
    wire N__10223;
    wire N__10222;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10208;
    wire N__10203;
    wire N__10196;
    wire N__10193;
    wire N__10178;
    wire N__10175;
    wire N__10174;
    wire N__10169;
    wire N__10166;
    wire N__10165;
    wire N__10162;
    wire N__10161;
    wire N__10160;
    wire N__10159;
    wire N__10158;
    wire N__10151;
    wire N__10150;
    wire N__10149;
    wire N__10144;
    wire N__10143;
    wire N__10142;
    wire N__10141;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10130;
    wire N__10129;
    wire N__10128;
    wire N__10125;
    wire N__10122;
    wire N__10117;
    wire N__10112;
    wire N__10107;
    wire N__10102;
    wire N__10097;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10033;
    wire N__10028;
    wire N__10027;
    wire N__10026;
    wire N__10025;
    wire N__10024;
    wire N__10023;
    wire N__10016;
    wire N__10013;
    wire N__10012;
    wire N__10011;
    wire N__10006;
    wire N__10003;
    wire N__10002;
    wire N__10001;
    wire N__10000;
    wire N__9999;
    wire N__9998;
    wire N__9997;
    wire N__9996;
    wire N__9995;
    wire N__9992;
    wire N__9987;
    wire N__9982;
    wire N__9977;
    wire N__9968;
    wire N__9963;
    wire N__9950;
    wire N__9947;
    wire N__9946;
    wire N__9945;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9933;
    wire N__9926;
    wire N__9925;
    wire N__9922;
    wire N__9921;
    wire N__9920;
    wire N__9919;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9907;
    wire N__9902;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9862;
    wire N__9859;
    wire N__9856;
    wire N__9853;
    wire N__9850;
    wire N__9845;
    wire N__9842;
    wire N__9841;
    wire N__9836;
    wire N__9833;
    wire N__9832;
    wire N__9831;
    wire N__9826;
    wire N__9825;
    wire N__9824;
    wire N__9823;
    wire N__9822;
    wire N__9821;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9806;
    wire N__9799;
    wire N__9788;
    wire N__9785;
    wire N__9782;
    wire N__9781;
    wire N__9780;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9766;
    wire N__9765;
    wire N__9764;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9752;
    wire N__9747;
    wire N__9742;
    wire N__9731;
    wire N__9728;
    wire N__9727;
    wire N__9726;
    wire N__9725;
    wire N__9724;
    wire N__9721;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9694;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9669;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9634;
    wire N__9633;
    wire N__9630;
    wire N__9627;
    wire N__9622;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9601;
    wire N__9600;
    wire N__9599;
    wire N__9598;
    wire N__9597;
    wire N__9586;
    wire N__9583;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9571;
    wire N__9568;
    wire N__9565;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9478;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9433;
    wire N__9430;
    wire N__9429;
    wire N__9428;
    wire N__9425;
    wire N__9424;
    wire N__9423;
    wire N__9422;
    wire N__9417;
    wire N__9408;
    wire N__9405;
    wire N__9398;
    wire N__9395;
    wire N__9394;
    wire N__9393;
    wire N__9392;
    wire N__9391;
    wire N__9390;
    wire N__9387;
    wire N__9384;
    wire N__9383;
    wire N__9378;
    wire N__9369;
    wire N__9366;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9220;
    wire N__9217;
    wire N__9216;
    wire N__9215;
    wire N__9214;
    wire N__9211;
    wire N__9210;
    wire N__9209;
    wire N__9206;
    wire N__9201;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9189;
    wire N__9184;
    wire N__9181;
    wire N__9170;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9158;
    wire N__9155;
    wire N__9154;
    wire N__9149;
    wire N__9146;
    wire N__9145;
    wire N__9144;
    wire N__9143;
    wire N__9142;
    wire N__9141;
    wire N__9136;
    wire N__9127;
    wire N__9122;
    wire N__9119;
    wire N__9118;
    wire N__9117;
    wire N__9114;
    wire N__9113;
    wire N__9108;
    wire N__9103;
    wire N__9098;
    wire N__9097;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9013;
    wire N__9012;
    wire N__9009;
    wire N__9008;
    wire N__9007;
    wire N__9004;
    wire N__9003;
    wire N__9002;
    wire N__9001;
    wire N__9000;
    wire N__8997;
    wire N__8996;
    wire N__8993;
    wire N__8988;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8967;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8899;
    wire N__8898;
    wire N__8897;
    wire N__8896;
    wire N__8895;
    wire N__8894;
    wire N__8893;
    wire N__8890;
    wire N__8885;
    wire N__8874;
    wire N__8867;
    wire N__8866;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8851;
    wire N__8848;
    wire N__8847;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8836;
    wire N__8833;
    wire N__8832;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8808;
    wire N__8801;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8777;
    wire N__8776;
    wire N__8775;
    wire N__8774;
    wire N__8773;
    wire N__8770;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8755;
    wire N__8752;
    wire N__8749;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8730;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8707;
    wire N__8704;
    wire N__8701;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8671;
    wire N__8670;
    wire N__8667;
    wire N__8666;
    wire N__8665;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8648;
    wire N__8647;
    wire N__8646;
    wire N__8643;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8625;
    wire N__8622;
    wire N__8617;
    wire N__8614;
    wire N__8597;
    wire N__8596;
    wire N__8593;
    wire N__8592;
    wire N__8591;
    wire N__8590;
    wire N__8589;
    wire N__8588;
    wire N__8587;
    wire N__8584;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8558;
    wire N__8553;
    wire N__8540;
    wire N__8539;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8531;
    wire N__8530;
    wire N__8529;
    wire N__8526;
    wire N__8525;
    wire N__8524;
    wire N__8523;
    wire N__8522;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8514;
    wire N__8513;
    wire N__8512;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8494;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8470;
    wire N__8465;
    wire N__8462;
    wire N__8455;
    wire N__8438;
    wire N__8435;
    wire N__8434;
    wire N__8433;
    wire N__8430;
    wire N__8429;
    wire N__8428;
    wire N__8427;
    wire N__8426;
    wire N__8425;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8393;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8371;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8348;
    wire N__8345;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8330;
    wire N__8329;
    wire N__8328;
    wire N__8325;
    wire N__8324;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8309;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8261;
    wire N__8258;
    wire N__8257;
    wire N__8256;
    wire N__8253;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8236;
    wire N__8233;
    wire N__8230;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8218;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8198;
    wire N__8195;
    wire N__8194;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8162;
    wire N__8159;
    wire N__8158;
    wire N__8155;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8139;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8116;
    wire N__8115;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8071;
    wire N__8068;
    wire N__8067;
    wire N__8066;
    wire N__8065;
    wire N__8064;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8049;
    wire N__8044;
    wire N__8041;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8023;
    wire N__8022;
    wire N__8017;
    wire N__8014;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7999;
    wire N__7998;
    wire N__7995;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7975;
    wire N__7970;
    wire N__7969;
    wire N__7966;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7940;
    wire N__7937;
    wire N__7936;
    wire N__7935;
    wire N__7934;
    wire N__7931;
    wire N__7924;
    wire N__7923;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7911;
    wire N__7904;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7858;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7846;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7816;
    wire N__7815;
    wire N__7810;
    wire N__7807;
    wire N__7802;
    wire N__7799;
    wire N__7798;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7770;
    wire N__7765;
    wire N__7760;
    wire N__7757;
    wire N__7756;
    wire N__7755;
    wire N__7752;
    wire N__7747;
    wire N__7742;
    wire N__7741;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7706;
    wire N__7705;
    wire N__7704;
    wire N__7703;
    wire N__7700;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7684;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7645;
    wire N__7642;
    wire N__7641;
    wire N__7640;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7619;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7597;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7574;
    wire N__7571;
    wire N__7570;
    wire N__7569;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7471;
    wire N__7468;
    wire N__7465;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7450;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7397;
    wire N__7396;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7388;
    wire N__7385;
    wire N__7382;
    wire N__7379;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7316;
    wire N__7315;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7273;
    wire N__7272;
    wire N__7271;
    wire N__7266;
    wire N__7263;
    wire N__7262;
    wire N__7261;
    wire N__7258;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7242;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire VCCG0;
    wire GNDG0;
    wire port_rw_c_i;
    wire port_nmib_c_i;
    wire \this_vga_signals.N_29_cascade_ ;
    wire \this_vga_signals.N_40_cascade_ ;
    wire \this_vga_signals.N_20 ;
    wire \this_vga_signals.N_18_cascade_ ;
    wire this_vga_signals_N_274_i;
    wire \this_vga_signals.hvisible_i_a2_0_3_0_cascade_ ;
    wire \this_vga_signals.M_hstate_qZ0Z_1 ;
    wire \this_vga_signals.N_49_cascade_ ;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire \this_vga_signals.N_32 ;
    wire \this_vga_signals.M_hstate_qZ0Z_0 ;
    wire \this_vga_signals.N_26 ;
    wire \this_vga_signals.N_26_cascade_ ;
    wire \this_vga_signals.N_51 ;
    wire \this_vga_signals.N_273 ;
    wire \this_vga_signals.N_2_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.N_70_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_1_0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.m44_0_0 ;
    wire \this_vga_signals.M_vcounter_q_RNIQE2J1Z0Z_9_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fast_RNI3BJLZ0Z_4 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1 ;
    wire \this_vga_signals.mult1_un40_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_2_cascade_ ;
    wire bfn_9_23_0_;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7NZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8NZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_7 ;
    wire bfn_9_24_0_;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_8 ;
    wire bfn_10_17_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_10_18_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_9 ;
    wire \this_vga_signals.M_hstate_d_0_sqmuxa ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_10 ;
    wire \this_vga_signals.g1_0_0_a2_0_cascade_ ;
    wire \this_vga_signals.g0_11_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KANZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.N_2 ;
    wire \this_vga_signals.i9_mux_cascade_ ;
    wire \this_vga_signals.i9_mux ;
    wire \this_vga_signals.address_1_c5_i ;
    wire port_nmib_c;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_9 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCNZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBNZ0 ;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire \this_vga_signals.address_1_c4_cascade_ ;
    wire \this_vga_signals.N_70 ;
    wire \this_vga_signals.SUM_0 ;
    wire \this_vga_signals.mult1_un40_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_c ;
    wire \this_vga_signals.mult1_un40_sum_axbxc1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un47_sum_c3_cascade_ ;
    wire \this_vga_signals.N_13_0 ;
    wire \this_vga_signals.if_i1_mux ;
    wire \this_vga_signals.M_vcounter_q_RNO_0Z0Z_3 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_ ;
    wire \this_vga_signals.address_m24_ns_1Z0Z_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c3 ;
    wire \this_vga_signals.mult1_un54_sum_c2_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_RNO_0Z0Z_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire bfn_11_17_0_;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire \this_vga_signals.un12_address_cry_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.un12_address_cry_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.un12_address_cry_2 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.un12_address_cry_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.un12_address_cry_4 ;
    wire \this_vga_signals.un12_address_cry_5 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.un12_address_cry_6 ;
    wire \this_vga_signals.un12_address_cry_7 ;
    wire bfn_11_18_0_;
    wire \this_vga_signals.un12_address_cry_8 ;
    wire \this_vga_signals.un12_address_cry_9 ;
    wire \this_vga_signals.un12_address_cry_10 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.N_49 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_11 ;
    wire N_16;
    wire \this_vga_signals.mult1_un61_sum_ac0_7_0_3_1_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_7_0_3_2 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.N_27 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.hvisible_i_a2_2_0 ;
    wire rgb_c_4;
    wire \this_vga_signals.m30_3 ;
    wire \this_vga_signals.m30_4_cascade_ ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.N_3_0_cascade_ ;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire rgb_c_0;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.address_m1_1_1 ;
    wire \this_vga_signals.mult1_un54_sum_c2 ;
    wire \this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c3_1 ;
    wire \this_vga_signals.mult1_un61_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un61_sum_c2 ;
    wire \this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2 ;
    wire \this_vga_signals.address_i3_mux_i ;
    wire \this_vga_signals.address_m27_ns_1_cascade_ ;
    wire \this_vga_signals.address_i2_mux_3_cascade_ ;
    wire \this_vga_signals.address_i2_mux_2 ;
    wire \this_vga_signals.M_vcounter_q_RNO_0Z0Z_1 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_8_cascade_ ;
    wire \this_vga_signals.g1_1_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_10 ;
    wire \this_vga_signals.M_hcounter_q_i_11 ;
    wire \this_vga_signals.un12_address_cry_9_THRU_CO ;
    wire \this_vga_signals.un12_address_cry_9_c_RNIVF1R ;
    wire \this_vga_signals.un12_address_cry_10_c_RNINP5K ;
    wire \this_vga_signals.un12_address_cry_9_c_RNIVF1R_cascade_ ;
    wire \this_vga_signals.un12_address_cry_9_c_RNIEJOE ;
    wire \this_vga_signals.mult1_un47_sum_c5_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb3_x1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb3_cascade_ ;
    wire \this_vga_signals.if_m5_sn ;
    wire \this_vga_signals.if_m5_rn_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c5_cascade_ ;
    wire M_this_vga_signals_address_4;
    wire \this_vga_signals.mult1_un61_sum_ac0_7_0_3 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c4 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_7_0_4_cascade_ ;
    wire \this_vga_signals.if_m4_0_1_cascade_ ;
    wire \this_vga_signals.G_12_0_x3_0_cascade_ ;
    wire vsync_c;
    wire \this_vga_signals.N_52_cascade_ ;
    wire \this_vga_signals.N_76_mux ;
    wire \this_vga_signals.N_76_mux_cascade_ ;
    wire \this_vga_signals.N_72_mux ;
    wire \this_vga_signals.N_55_cascade_ ;
    wire \this_vga_signals.M_vstate_q_RNO_1Z0Z_0_cascade_ ;
    wire \this_vga_signals.M_vstate_q_RNO_2Z0Z_0 ;
    wire \this_vga_signals.M_vstate_qZ0Z_1 ;
    wire \this_vga_signals.m35_e_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c2 ;
    wire \this_vga_signals.address_N_9_0_cascade_ ;
    wire \this_vga_signals.address_N_10_0 ;
    wire \this_vga_signals.address_N_3 ;
    wire \this_vga_signals.M_vcounter_q_RNITV8S_2Z0Z_0 ;
    wire \this_vga_signals.M_vcounter_q_RNI8OSG6BZ0Z_2_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb1_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3 ;
    wire \this_vga_signals.address_m35_1 ;
    wire \this_vga_signals.N_75_mux ;
    wire \this_vga_signals.N_84 ;
    wire \this_vga_signals.M_vcounter_q_RNO_0Z0Z_2 ;
    wire \this_vga_signals.address_m31_1 ;
    wire \this_vga_signals.address_i2_mux_4 ;
    wire \this_vga_signals.M_vcounter_q_RNITV8S_1Z0Z_0 ;
    wire \this_vga_signals.address_N_9_0 ;
    wire \this_vga_signals.address_N_33_cascade_ ;
    wire \this_vga_signals.address_N_34 ;
    wire \this_vga_signals.g1_1 ;
    wire \this_vga_signals.mult1_un61_sum_axb3_0_cascade_ ;
    wire \this_vga_signals.g0_4_0_1_cascade_ ;
    wire \this_vga_signals.g1_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_axb3_out ;
    wire \this_vga_signals.mult1_un54_sum_axb4 ;
    wire \this_vga_signals.mult1_un47_sum_c5 ;
    wire \this_vga_signals.mult1_un61_sum_axb4_x0 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_7_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb4_x1 ;
    wire \this_vga_signals.mult1_un61_sum_axb4_i_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_5_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb4_i ;
    wire \this_vga_signals.g0_6_0_0_1 ;
    wire this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_;
    wire \this_vga_signals.mult1_un61_sum_axb3 ;
    wire \this_vga_signals.if_m4_0_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc5 ;
    wire \this_vga_signals.un12_address_cry_7_c_RNI32HB ;
    wire \this_vga_signals.if_m2_3_0 ;
    wire \this_vga_signals.mult1_un61_sum_axb3_1 ;
    wire \this_vga_signals.G_12_0_3_1 ;
    wire \this_vga_signals.N_9_cascade_ ;
    wire \this_vga_signals.G_12_0_3_cascade_ ;
    wire \this_vga_signals.if_m4_0_1 ;
    wire this_vga_signals_un17_address_if_N_8_mux_cascade_;
    wire \this_vga_signals.N_10_0 ;
    wire N_6_i_cascade_;
    wire \this_vga_signals.N_18_0 ;
    wire \this_vga_signals.g0_6_1 ;
    wire \this_vga_signals.G_12_0_x3_0 ;
    wire N_11_0_cascade_;
    wire \this_vga_signals.N_5_i ;
    wire \this_vga_signals.G_12_0_1 ;
    wire \this_vga_signals.N_25 ;
    wire \this_vga_signals.M_vstate_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.N_275 ;
    wire \this_vga_signals.if_N_9_i_i_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_ ;
    wire M_this_vga_signals_address_8;
    wire \this_vga_signals.address_m6_0_1_cascade_ ;
    wire \this_vga_signals.address_mZ0Z1 ;
    wire \this_vga_signals.address_i2_mux_cascade_ ;
    wire \this_vga_signals.address_N_11 ;
    wire \this_vga_signals.address_i2_mux_0 ;
    wire \this_vga_signals.address_m21_ns_1_cascade_ ;
    wire \this_vga_signals.address_i2_mux_1 ;
    wire \this_vga_signals.address_N_22_cascade_ ;
    wire \this_vga_signals.address_N_36 ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.mult1_un61_sum_axb1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_0 ;
    wire \this_vga_signals.if_m16_0_o4 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.address_N_40 ;
    wire \this_vga_signals.if_m4_0_1_0_0 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc5_1_N_3L3_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc5_1_N_2L1 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5_cascade_ ;
    wire \this_vga_signals.N_21_0 ;
    wire \this_vga_signals.g0_6_0_0_2 ;
    wire \this_vga_signals.if_N_8_mux_2_2 ;
    wire \this_vga_signals.mult1_un82_sum_axb3_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_4 ;
    wire \this_vga_signals.g0_i_x4_4_a3_1 ;
    wire \this_vga_signals.if_m1_0 ;
    wire \this_vga_signals.if_N_3_3_i ;
    wire this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5_cascade_;
    wire \this_vga_signals.if_N_3_2_i_cascade_ ;
    wire M_this_vga_signals_address_3;
    wire \this_vga_signals.mult1_un61_sum_ac0_7_0_4 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_5 ;
    wire \this_vga_signals.N_12 ;
    wire \this_vga_signals.g0_0_0_a2_1_0_cascade_ ;
    wire \this_vga_signals.if_N_3_2_i_3_1_cascade_ ;
    wire \this_vga_signals.N_31 ;
    wire \this_vga_signals.N_20_i_i ;
    wire \this_vga_signals.N_20_i_i_cascade_ ;
    wire \this_vga_signals.N_26_i_i ;
    wire \this_vga_signals.mult1_un47_sum_c3 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_1 ;
    wire \this_vga_signals.mult1_un68_sum_c3 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0 ;
    wire M_this_vga_signals_address_9;
    wire \this_vga_signals.mult1_un54_sum_ac0_7 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_8 ;
    wire M_this_vga_signals_address_6;
    wire \this_vga_signals.N_4 ;
    wire \this_vram.M_this_vram_read_data_1_cascade_ ;
    wire rgb_c_2;
    wire \this_vga_signals.g0_4 ;
    wire \this_vga_signals.if_N_8_mux_2_2_1 ;
    wire \this_vga_signals.N_3_1_0_1_cascade_ ;
    wire \this_vga_signals.g1_2_0_0 ;
    wire \this_vga_signals.g0_0_0_0 ;
    wire \this_vga_signals.if_m1_0_0 ;
    wire \this_vga_signals.N_21 ;
    wire \this_vga_signals.g0_3 ;
    wire \this_vga_signals.N_20_i_i_0 ;
    wire \this_vga_signals.g0_0_a3_3 ;
    wire \this_vga_signals.mult1_un82_sum_ac0_7_0_1_0 ;
    wire \this_vga_signals.N_11_cascade_ ;
    wire \this_vga_signals.g0_0_a3_2 ;
    wire \this_vga_signals.g0_0_a3_5_cascade_ ;
    wire \this_vga_signals.g0_i_x4_4_a3 ;
    wire \this_vga_signals.N_3_3_0 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_1 ;
    wire \this_vga_signals.g0_0_1_0 ;
    wire \this_vga_signals.g1_5_0_0_cascade_ ;
    wire \this_vga_signals.r_N_2_0_0_0 ;
    wire \this_vga_signals.g0_1_0 ;
    wire \this_vga_signals.g0_1_2_cascade_ ;
    wire this_vga_signals_un17_address_if_N_8_mux;
    wire \this_vga_signals.g0_3_0_a2_1_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_ac0_7_0_1_2 ;
    wire \this_vga_signals.if_N_8_mux_2_0 ;
    wire this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5;
    wire \this_vga_signals.if_N_3_2_i ;
    wire \this_vga_signals.g1_0_0_0 ;
    wire this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0;
    wire \this_vga_signals.g0_6_0 ;
    wire \this_vga_signals.g1_2_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5 ;
    wire \this_vga_signals.g1_5_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb3 ;
    wire \this_vga_signals.g0_0_1_1 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_2_cascade_ ;
    wire \this_vga_signals.g1_0_0_0_0 ;
    wire \this_vga_signals.g0_0_3_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_ac0_7_0_1_4 ;
    wire \this_vga_signals.g0_6 ;
    wire \this_vga_signals.g0_13 ;
    wire \this_vga_signals.if_N_3_2_i_0 ;
    wire \this_vga_signals.g0_0_0_a2_1 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_0 ;
    wire \this_vga_signals.g1_2_cascade_ ;
    wire \this_vga_signals.r_N_2_0_0_2_cascade_ ;
    wire \this_vga_signals.N_3_1_1 ;
    wire \this_vga_signals.g0_3_1 ;
    wire \this_vga_signals.mult1_un68_sum_c5 ;
    wire \this_vga_signals.un12_address_cry_3_c_RNIRLCB ;
    wire \this_vga_signals.g0_5_3_cascade_ ;
    wire \this_vga_signals.un12_address_cry_2_c_RNIPIBB ;
    wire \this_vga_signals.un12_address_cry_1_c_RNINFAB ;
    wire \this_vga_signals.mult1_un96_sum_c5_0_1_0_1_cascade_ ;
    wire \this_vga_signals.N_3_1_2 ;
    wire \this_vga_signals.g1_0_0_0_1 ;
    wire \this_vga_signals.mult1_un96_sum_c5_cascade_ ;
    wire \this_vga_signals.g2_0 ;
    wire \this_vga_signals.mult1_un96_sum_axbxc5_2 ;
    wire \this_vga_signals.g1_0_3_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_c5_0_0_0_0 ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.g1_0_0 ;
    wire \this_vga_signals.if_N_3_2_i_1 ;
    wire \this_vga_signals.un12_address_cry_4_c_RNITODB ;
    wire \this_vga_signals.mult1_un75_sum_axbxc5 ;
    wire \this_vga_signals.mult1_un82_sum_ac0_7_0_1_3 ;
    wire \this_vga_signals.un12_address_cry_5_c_RNIVREB ;
    wire this_vga_signals_un17_address_if_m2_2_0;
    wire \this_vga_signals.g0_38 ;
    wire \this_vga_signals.N_4_0_1 ;
    wire \this_vga_signals.if_N_3_2_i_2_0 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_0 ;
    wire port_clk_c;
    wire this_start_data_delay_this_edge_detector_M_last_q;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_0 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_3 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_1 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_2 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_5 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_1 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_2 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_3 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_4 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_10 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_9 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_6 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_4 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_5 ;
    wire \this_vga_signals.mult1_un61_sum_c3 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1 ;
    wire M_this_vga_signals_address_10;
    wire \this_vram.M_this_vram_read_data_0 ;
    wire \this_vram.N_17_0 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_11 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_12 ;
    wire debug_d;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_13 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_14 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_15 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_16 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_17 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_18 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_7 ;
    wire \this_start_data_delay.this_delay.M_pipe_qZ0Z_8 ;
    wire \this_start_data_delay.this_edge_detector.N_215 ;
    wire \this_start_data_delay.this_edge_detector.N_212 ;
    wire \this_start_data_delay.this_edge_detector.N_219 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_8 ;
    wire port_data_c_5;
    wire \this_start_data_delay.this_edge_detector.N_222 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_6 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_7 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_9 ;
    wire bfn_19_23_0_;
    wire un1_M_current_address_q_cry_0;
    wire M_current_address_qZ0Z_2;
    wire un1_M_current_address_q_cry_1_c_RNI4TBNZ0;
    wire un1_M_current_address_q_cry_1;
    wire un1_M_current_address_q_cry_2;
    wire un1_M_current_address_q_cry_3_c_RNI83ENZ0;
    wire un1_M_current_address_q_cry_3;
    wire M_current_address_qZ0Z_5;
    wire un1_M_current_address_q_cry_4_c_RNIA6FNZ0;
    wire un1_M_current_address_q_cry_4;
    wire un1_M_current_address_q_cry_5;
    wire un1_M_current_address_q_cry_6;
    wire un1_M_current_address_q_cry_7;
    wire un1_M_current_address_q_cry_7_c_RNIGFINZ0;
    wire bfn_19_24_0_;
    wire M_current_address_qZ0Z_9;
    wire un1_M_current_address_q_cry_8_c_RNIIIJNZ0;
    wire un1_M_current_address_q_cry_8;
    wire un1_M_current_address_q_cry_9;
    wire un1_M_current_address_q_cry_10;
    wire un1_M_current_address_q_cry_11_c_RNI6NLHZ0;
    wire un1_M_current_address_q_cry_11;
    wire un1_M_current_address_q_cry_12;
    wire N_177_0;
    wire un1_M_current_address_q_cry_9_c_RNIRDIMZ0;
    wire un1_M_current_address_q_cry_0_c_RNI2QANZ0;
    wire un1_M_current_address_q_cry_12_c_RNI8QMHZ0;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_12 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_10 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_11 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_13 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_14 ;
    wire M_current_address_q_RNIHDTUZ0Z_0;
    wire un1_M_current_address_q_cry_5_c_RNIC9GNZ0;
    wire un1_M_current_address_q_cry_6_c_RNIECHNZ0;
    wire un1_M_current_address_q_cry_10_c_RNI4KKHZ0;
    wire un1_M_current_address_q_cry_2_c_RNI60DNZ0;
    wire N_339_g;
    wire M_current_address_qZ0Z_6;
    wire \this_start_data_delay.this_edge_detector.N_216 ;
    wire M_current_address_qZ0Z_3;
    wire \this_start_data_delay.this_edge_detector.N_213 ;
    wire M_current_address_qZ0Z_8;
    wire \this_start_data_delay.this_edge_detector.N_218 ;
    wire M_current_address_qZ0Z_10;
    wire \this_start_data_delay.this_edge_detector.N_220 ;
    wire \this_start_data_delay.this_edge_detector.N_221 ;
    wire port_data_c_6;
    wire \this_start_data_delay.this_edge_detector.N_223 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_15 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_16 ;
    wire M_current_address_qZ0Z_7;
    wire \this_start_data_delay.this_edge_detector.N_217 ;
    wire M_current_address_qZ0Z_0;
    wire \this_start_data_delay.this_edge_detector.N_210 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_17 ;
    wire \this_start_address_delay.this_delay.M_pipe_qZ0Z_18 ;
    wire M_this_start_address_delay_out_0;
    wire M_state_q_ns_1_0__N_24_mux_cascade_;
    wire M_state_q_ns_1_0__N_10_cascade_;
    wire M_current_address_qZ0Z_1;
    wire \this_start_data_delay.this_edge_detector.N_211 ;
    wire M_current_address_qZ0Z_4;
    wire port_data_c_4;
    wire \this_start_data_delay.this_edge_detector.N_214 ;
    wire M_state_qZ0Z_0;
    wire port_address_c_1;
    wire M_state_q_ns_1_0__N_24_mux;
    wire port_address_c_0;
    wire M_this_reset_cond_out_0;
    wire M_this_start_data_delay_out_0;
    wire M_state_q_ns_1_0__i12_mux_cascade_;
    wire M_state_qZ0Z_1;
    wire clk_c_g;
    wire port_data_c_0;
    wire M_this_vram_write_data_0;
    wire \this_vram.mem_WE_8 ;
    wire \this_vram.mem_N_91 ;
    wire \this_vram.mem_N_88 ;
    wire N_16_0;
    wire port_address_c_4;
    wire port_address_c_7;
    wire port_enb_c;
    wire port_address_c_2;
    wire M_state_q_ns_1_0__m7Z0Z_5;
    wire port_data_c_1;
    wire M_this_vram_write_data_1;
    wire \this_vram.mem_out_bus2_1 ;
    wire \this_vram.mem_out_bus6_1 ;
    wire \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0 ;
    wire \this_vram.mem_WE_14 ;
    wire \this_vram.mem_WE_10 ;
    wire M_this_vram_read_data_3;
    wire \this_vram.mem_out_bus4_1 ;
    wire \this_vram.mem_out_bus0_1 ;
    wire \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0 ;
    wire \this_vram.mem_out_bus7_3 ;
    wire \this_vram.mem_out_bus3_3 ;
    wire \this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_ ;
    wire \this_vram.mem_N_102 ;
    wire \this_vram.mem_radregZ0Z_11 ;
    wire M_this_vram_read_data_2;
    wire \this_vram.mem_WE_12 ;
    wire \this_vram.mem_N_109 ;
    wire CONSTANT_ONE_NET;
    wire \this_vga_signals.mult1_un61_sum_axbxc5 ;
    wire M_this_vga_signals_address_5;
    wire \this_vram.mem_out_bus1_2 ;
    wire \this_vram.mem_out_bus5_2 ;
    wire \this_vram.mem_out_bus1_1 ;
    wire \this_vram.mem_out_bus5_1 ;
    wire \this_vram.mem_mem_1_0_RNISSK11Z0Z_0 ;
    wire \this_vram.mem_out_bus6_0 ;
    wire \this_vram.mem_out_bus2_0 ;
    wire \this_vram.mem_mem_2_0_RNIU0NZ0Z11_cascade_ ;
    wire \this_vram.mem_N_112 ;
    wire \this_vram.mem_out_bus4_0 ;
    wire \this_vram.mem_out_bus0_0 ;
    wire \this_vram.mem_mem_0_0_RNIQOIZ0Z11 ;
    wire \this_vram.mem_out_bus3_2 ;
    wire \this_vram.mem_out_bus7_2 ;
    wire \this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_ ;
    wire \this_vram.mem_mem_1_1_RNIUSKZ0Z11 ;
    wire \this_vram.mem_N_95 ;
    wire \this_vram.mem_out_bus5_3 ;
    wire \this_vram.mem_out_bus1_3 ;
    wire \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0 ;
    wire \this_vram.mem_out_bus3_0 ;
    wire \this_vram.mem_out_bus7_0 ;
    wire \this_vram.mem_mem_3_0_RNI05PZ0Z11 ;
    wire \this_vram.mem_out_bus6_3 ;
    wire \this_vram.mem_out_bus2_3 ;
    wire \this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_ ;
    wire \this_vram.mem_N_105 ;
    wire \this_vram.mem_out_bus0_3 ;
    wire \this_vram.mem_out_bus4_3 ;
    wire \this_vram.mem_mem_0_1_RNISOI11Z0Z_0 ;
    wire \this_vram.mem_out_bus2_2 ;
    wire \this_vram.mem_out_bus6_2 ;
    wire \this_vram.mem_out_bus0_2 ;
    wire \this_vram.mem_out_bus4_2 ;
    wire \this_vram.mem_mem_2_1_RNI01NZ0Z11 ;
    wire \this_vram.mem_mem_0_1_RNISOIZ0Z11_cascade_ ;
    wire \this_vram.mem_radregZ0Z_12 ;
    wire \this_vram.mem_N_98 ;
    wire \this_vram.mem_out_bus1_0 ;
    wire \this_vram.mem_out_bus5_0 ;
    wire \this_vram.mem_mem_1_0_RNISSKZ0Z11 ;
    wire \this_vram.mem_radregZ0Z_13 ;
    wire \this_vram.mem_out_bus7_1 ;
    wire \this_vram.mem_out_bus3_1 ;
    wire \this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ;
    wire \this_vram.mem_WE_6 ;
    wire \this_vram.mem_WE_4 ;
    wire \this_vram.mem_WE_2 ;
    wire M_current_address_qZ0Z_12;
    wire M_current_address_qZ0Z_11;
    wire M_current_address_qZ0Z_13;
    wire \this_vram.mem_WE_0 ;
    wire port_data_c_2;
    wire M_this_vram_write_data_2;
    wire port_data_c_3;
    wire M_this_vram_write_en_0_sqmuxa;
    wire M_this_vram_write_data_3;
    wire \this_vga_signals.g0_7 ;
    wire \this_vga_signals.mult1_un89_sum_c5 ;
    wire M_this_vga_signals_address_1;
    wire \this_vga_signals.rgb72 ;
    wire \this_vga_signals.mult1_un82_sum_c5 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc5_1_i ;
    wire M_this_vga_signals_address_2;
    wire port_rw_c;
    wire port_address_c_6;
    wire port_address_c_5;
    wire port_address_c_3;
    wire M_state_q_ns_1_0__m7Z0Z_4;
    wire _gnd_net_;

    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,\this_vram.mem_out_bus0_1 ,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,\this_vram.mem_out_bus0_0 ,dangling_wire_11,dangling_wire_12,dangling_wire_13}),
            .RADDR({N__14252,N__11510,N__10451,N__11156,N__12218,N__18278,N__9338,N__11342,N__19814,N__20120,N__13949}),
            .WADDR({N__16013,N__14900,N__16145,N__15821,N__15386,N__15050,N__16529,N__15263,N__14687,N__16661,N__15686}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,N__16793,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__17111,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .RCLKE(),
            .RCLK(N__17302),
            .RE(N__18695),
            .WCLKE(N__17984),
            .WCLK(N__17303),
            .WE(N__18610));
    defparam \this_vram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,\this_vram.mem_out_bus0_3 ,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,\this_vram.mem_out_bus0_2 ,dangling_wire_55,dangling_wire_56,dangling_wire_57}),
            .RADDR({N__14246,N__11504,N__10445,N__11150,N__12212,N__18272,N__9332,N__11336,N__19808,N__20114,N__13943}),
            .WADDR({N__16007,N__14894,N__16139,N__15815,N__15380,N__15044,N__16523,N__15257,N__14681,N__16655,N__15680}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,N__20228,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,N__18996,dangling_wire_85,dangling_wire_86,dangling_wire_87}),
            .RCLKE(),
            .RCLK(N__17304),
            .RE(N__18691),
            .WCLKE(N__17980),
            .WCLK(N__17305),
            .WE(N__18688));
    defparam \this_vram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,\this_vram.mem_out_bus1_1 ,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,\this_vram.mem_out_bus1_0 ,dangling_wire_99,dangling_wire_100,dangling_wire_101}),
            .RADDR({N__14240,N__11498,N__10439,N__11144,N__12206,N__18266,N__9326,N__11330,N__19802,N__20108,N__13937}),
            .WADDR({N__16001,N__14888,N__16133,N__15809,N__15374,N__15038,N__16517,N__15251,N__14675,N__16649,N__15674}),
            .MASK({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .WDATA({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__16789,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__17107,dangling_wire_129,dangling_wire_130,dangling_wire_131}),
            .RCLKE(),
            .RCLK(N__17306),
            .RE(N__18690),
            .WCLKE(N__17771),
            .WCLK(N__17307),
            .WE(N__18687));
    defparam \this_vram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,\this_vram.mem_out_bus1_3 ,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,\this_vram.mem_out_bus1_2 ,dangling_wire_143,dangling_wire_144,dangling_wire_145}),
            .RADDR({N__14234,N__11492,N__10433,N__11138,N__12200,N__18260,N__9320,N__11324,N__19796,N__20102,N__13931}),
            .WADDR({N__15995,N__14882,N__16127,N__15803,N__15368,N__15032,N__16511,N__15245,N__14669,N__16643,N__15668}),
            .MASK({dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161}),
            .WDATA({dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,N__20224,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,N__19001,dangling_wire_173,dangling_wire_174,dangling_wire_175}),
            .RCLKE(),
            .RCLK(N__17308),
            .RE(N__18666),
            .WCLKE(N__17767),
            .WCLK(N__17309),
            .WE(N__18677));
    defparam \this_vram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,\this_vram.mem_out_bus2_1 ,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,\this_vram.mem_out_bus2_0 ,dangling_wire_187,dangling_wire_188,dangling_wire_189}),
            .RADDR({N__14228,N__11486,N__10427,N__11132,N__12194,N__18254,N__9314,N__11318,N__19790,N__20096,N__13925}),
            .WADDR({N__15989,N__14876,N__16121,N__15797,N__15362,N__15026,N__16505,N__15239,N__14663,N__16637,N__15662}),
            .MASK({dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205}),
            .WDATA({dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,N__16782,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,N__17100,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .RCLKE(),
            .RCLK(N__17311),
            .RE(N__18665),
            .WCLKE(N__17951),
            .WCLK(N__17310),
            .WE(N__18609));
    defparam \this_vram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,\this_vram.mem_out_bus2_3 ,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,\this_vram.mem_out_bus2_2 ,dangling_wire_231,dangling_wire_232,dangling_wire_233}),
            .RADDR({N__14222,N__11480,N__10421,N__11126,N__12188,N__18248,N__9308,N__11312,N__19784,N__20090,N__13919}),
            .WADDR({N__15983,N__14870,N__16115,N__15791,N__15356,N__15020,N__16499,N__15233,N__14657,N__16631,N__15656}),
            .MASK({dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249}),
            .WDATA({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,N__20217,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,N__18997,dangling_wire_261,dangling_wire_262,dangling_wire_263}),
            .RCLKE(),
            .RCLK(N__17313),
            .RE(N__18634),
            .WCLKE(N__17947),
            .WCLK(N__17314),
            .WE(N__18654));
    defparam \this_vram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,\this_vram.mem_out_bus3_1 ,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,\this_vram.mem_out_bus3_0 ,dangling_wire_275,dangling_wire_276,dangling_wire_277}),
            .RADDR({N__14216,N__11474,N__10415,N__11120,N__12182,N__18242,N__9302,N__11306,N__19778,N__20084,N__13913}),
            .WADDR({N__15977,N__14864,N__16109,N__15785,N__15350,N__15014,N__16493,N__15227,N__14651,N__16625,N__15650}),
            .MASK({dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293}),
            .WDATA({dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,N__16772,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,N__17091,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .RCLKE(),
            .RCLK(N__17321),
            .RE(N__18633),
            .WCLKE(N__17036),
            .WCLK(N__17322),
            .WE(N__18563));
    defparam \this_vram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,\this_vram.mem_out_bus3_3 ,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,\this_vram.mem_out_bus3_2 ,dangling_wire_319,dangling_wire_320,dangling_wire_321}),
            .RADDR({N__14210,N__11468,N__10409,N__11114,N__12176,N__18236,N__9296,N__11300,N__19772,N__20078,N__13907}),
            .WADDR({N__15971,N__14858,N__16103,N__15779,N__15344,N__15008,N__16487,N__15221,N__14645,N__16619,N__15644}),
            .MASK({dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337}),
            .WDATA({dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,N__20208,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,N__18989,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .RCLKE(),
            .RCLK(N__17334),
            .RE(N__18595),
            .WCLKE(N__17032),
            .WCLK(N__17335),
            .WE(N__18624));
    defparam \this_vram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,\this_vram.mem_out_bus4_1 ,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,\this_vram.mem_out_bus4_0 ,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .RADDR({N__14204,N__11462,N__10403,N__11108,N__12170,N__18230,N__9290,N__11294,N__19766,N__20072,N__13901}),
            .WADDR({N__15965,N__14852,N__16097,N__15773,N__15338,N__15002,N__16481,N__15215,N__14639,N__16613,N__15638}),
            .MASK({dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381}),
            .WDATA({dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,N__16760,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,N__17082,dangling_wire_393,dangling_wire_394,dangling_wire_395}),
            .RCLKE(),
            .RCLK(N__17344),
            .RE(N__18594),
            .WCLKE(N__19403),
            .WCLK(N__17345),
            .WE(N__18575));
    defparam \this_vram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,\this_vram.mem_out_bus4_3 ,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,\this_vram.mem_out_bus4_2 ,dangling_wire_407,dangling_wire_408,dangling_wire_409}),
            .RADDR({N__14198,N__11456,N__10397,N__11102,N__12164,N__18224,N__9284,N__11288,N__19760,N__20066,N__13895}),
            .WADDR({N__15959,N__14846,N__16091,N__15767,N__15332,N__14996,N__16475,N__15209,N__14633,N__16607,N__15632}),
            .MASK({dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425}),
            .WDATA({dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,N__20199,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,N__18977,dangling_wire_437,dangling_wire_438,dangling_wire_439}),
            .RCLKE(),
            .RCLK(N__17355),
            .RE(N__18515),
            .WCLKE(N__19399),
            .WCLK(N__17356),
            .WE(N__18562));
    defparam \this_vram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,\this_vram.mem_out_bus5_1 ,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,\this_vram.mem_out_bus5_0 ,dangling_wire_451,dangling_wire_452,dangling_wire_453}),
            .RADDR({N__14192,N__11450,N__10391,N__11096,N__12158,N__18218,N__9278,N__11282,N__19754,N__20060,N__13889}),
            .WADDR({N__15953,N__14840,N__16085,N__15761,N__15326,N__14990,N__16469,N__15203,N__14627,N__16601,N__15626}),
            .MASK({dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469}),
            .WDATA({dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,N__16748,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,N__17073,dangling_wire_481,dangling_wire_482,dangling_wire_483}),
            .RCLKE(),
            .RCLK(N__17366),
            .RE(N__18514),
            .WCLKE(N__19376),
            .WCLK(N__17367),
            .WE(N__18495));
    defparam \this_vram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,\this_vram.mem_out_bus5_3 ,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,\this_vram.mem_out_bus5_2 ,dangling_wire_495,dangling_wire_496,dangling_wire_497}),
            .RADDR({N__14186,N__11444,N__10385,N__11090,N__12152,N__18212,N__9272,N__11276,N__19748,N__20054,N__13883}),
            .WADDR({N__15947,N__14834,N__16079,N__15755,N__15320,N__14984,N__16463,N__15197,N__14621,N__16595,N__15620}),
            .MASK({dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513}),
            .WDATA({dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,N__20189,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,N__18964,dangling_wire_525,dangling_wire_526,dangling_wire_527}),
            .RCLKE(),
            .RCLK(N__17369),
            .RE(N__18519),
            .WCLKE(N__19372),
            .WCLK(N__17370),
            .WE(N__18521));
    defparam \this_vram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,\this_vram.mem_out_bus6_1 ,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,\this_vram.mem_out_bus6_0 ,dangling_wire_539,dangling_wire_540,dangling_wire_541}),
            .RADDR({N__14180,N__11438,N__10379,N__11084,N__12146,N__18206,N__9266,N__11270,N__19742,N__20048,N__13877}),
            .WADDR({N__15941,N__14828,N__16073,N__15749,N__15314,N__14978,N__16457,N__15191,N__14615,N__16589,N__15614}),
            .MASK({dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557}),
            .WDATA({dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,N__16732,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,N__17063,dangling_wire_569,dangling_wire_570,dangling_wire_571}),
            .RCLKE(),
            .RCLK(N__17371),
            .RE(N__18520),
            .WCLKE(N__19348),
            .WCLK(N__17372),
            .WE(N__18522));
    defparam \this_vram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,\this_vram.mem_out_bus6_3 ,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,\this_vram.mem_out_bus6_2 ,dangling_wire_583,dangling_wire_584,dangling_wire_585}),
            .RADDR({N__14174,N__11432,N__10373,N__11078,N__12140,N__18200,N__9260,N__11264,N__19736,N__20042,N__13871}),
            .WADDR({N__15935,N__14822,N__16067,N__15743,N__15308,N__14972,N__16451,N__15185,N__14609,N__16583,N__15608}),
            .MASK({dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601}),
            .WDATA({dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,N__20168,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,N__18960,dangling_wire_613,dangling_wire_614,dangling_wire_615}),
            .RCLKE(),
            .RCLK(N__17373),
            .RE(N__18576),
            .WCLKE(N__19349),
            .WCLK(N__17374),
            .WE(N__18581));
    defparam \this_vram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,\this_vram.mem_out_bus7_1 ,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,\this_vram.mem_out_bus7_0 ,dangling_wire_627,dangling_wire_628,dangling_wire_629}),
            .RADDR({N__14168,N__11426,N__10367,N__11072,N__12134,N__18194,N__9254,N__11258,N__19730,N__20036,N__13865}),
            .WADDR({N__15929,N__14816,N__16061,N__15737,N__15302,N__14966,N__16445,N__15179,N__14603,N__16577,N__15602}),
            .MASK({dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645}),
            .WDATA({dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,N__16747,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,N__17072,dangling_wire_657,dangling_wire_658,dangling_wire_659}),
            .RCLKE(),
            .RCLK(N__17375),
            .RE(N__18577),
            .WCLKE(N__19057),
            .WCLK(N__17376),
            .WE(N__18582));
    defparam \this_vram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,\this_vram.mem_out_bus7_3 ,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,\this_vram.mem_out_bus7_2 ,dangling_wire_671,dangling_wire_672,dangling_wire_673}),
            .RADDR({N__14162,N__11420,N__10361,N__11066,N__12128,N__18188,N__9248,N__11252,N__19724,N__20030,N__13859}),
            .WADDR({N__15923,N__14810,N__16055,N__15731,N__15296,N__14960,N__16439,N__15173,N__14597,N__16571,N__15596}),
            .MASK({dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689}),
            .WDATA({dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,N__20190,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,N__18976,dangling_wire_701,dangling_wire_702,dangling_wire_703}),
            .RCLKE(),
            .RCLK(N__17377),
            .RE(N__18623),
            .WCLKE(N__19058),
            .WCLK(N__17378),
            .WE(N__18622));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__20688),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__20690),
            .DIN(N__20689),
            .DOUT(N__20688),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__20690),
            .PADOUT(N__20689),
            .PADIN(N__20688),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_iopad (
            .OE(N__20679),
            .DIN(N__20678),
            .DOUT(N__20677),
            .PACKAGEPIN(debug));
    defparam debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_preio (
            .PADOEN(N__20679),
            .PADOUT(N__20678),
            .PADIN(N__20677),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14453),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__20670),
            .DIN(N__20669),
            .DOUT(N__20668),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__20670),
            .PADOUT(N__20669),
            .PADIN(N__20668),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8300),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__20661),
            .DIN(N__20660),
            .DOUT(N__20659),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__20661),
            .PADOUT(N__20660),
            .PADIN(N__20659),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7298),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_0_iopad (
            .OE(N__20652),
            .DIN(N__20651),
            .DOUT(N__20650),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_0_preio (
            .PADOEN(N__20652),
            .PADOUT(N__20651),
            .PADIN(N__20650),
            .CLOCKENABLE(),
            .DIN0(port_address_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_1_iopad (
            .OE(N__20643),
            .DIN(N__20642),
            .DOUT(N__20641),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_1_preio (
            .PADOEN(N__20643),
            .PADOUT(N__20642),
            .PADIN(N__20641),
            .CLOCKENABLE(),
            .DIN0(port_address_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_2_iopad (
            .OE(N__20634),
            .DIN(N__20633),
            .DOUT(N__20632),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_2_preio (
            .PADOEN(N__20634),
            .PADOUT(N__20633),
            .PADIN(N__20632),
            .CLOCKENABLE(),
            .DIN0(port_address_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_3_iopad (
            .OE(N__20625),
            .DIN(N__20624),
            .DOUT(N__20623),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_3_preio (
            .PADOEN(N__20625),
            .PADOUT(N__20624),
            .PADIN(N__20623),
            .CLOCKENABLE(),
            .DIN0(port_address_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_4_iopad (
            .OE(N__20616),
            .DIN(N__20615),
            .DOUT(N__20614),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_4_preio (
            .PADOEN(N__20616),
            .PADOUT(N__20615),
            .PADIN(N__20614),
            .CLOCKENABLE(),
            .DIN0(port_address_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_5_iopad (
            .OE(N__20607),
            .DIN(N__20606),
            .DOUT(N__20605),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_5_preio (
            .PADOEN(N__20607),
            .PADOUT(N__20606),
            .PADIN(N__20605),
            .CLOCKENABLE(),
            .DIN0(port_address_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_6_iopad (
            .OE(N__20598),
            .DIN(N__20597),
            .DOUT(N__20596),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_6_preio (
            .PADOEN(N__20598),
            .PADOUT(N__20597),
            .PADIN(N__20596),
            .CLOCKENABLE(),
            .DIN0(port_address_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_ibuf_7_iopad (
            .OE(N__20589),
            .DIN(N__20588),
            .DOUT(N__20587),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_address_ibuf_7_preio (
            .PADOEN(N__20589),
            .PADOUT(N__20588),
            .PADIN(N__20587),
            .CLOCKENABLE(),
            .DIN0(port_address_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__20580),
            .DIN(N__20579),
            .DOUT(N__20578),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__20580),
            .PADOUT(N__20579),
            .PADIN(N__20578),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__20571),
            .DIN(N__20570),
            .DOUT(N__20569),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__20571),
            .PADOUT(N__20570),
            .PADIN(N__20569),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__20562),
            .DIN(N__20561),
            .DOUT(N__20560),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__20562),
            .PADOUT(N__20561),
            .PADIN(N__20560),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__20553),
            .DIN(N__20552),
            .DOUT(N__20551),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__20553),
            .PADOUT(N__20552),
            .PADIN(N__20551),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__20544),
            .DIN(N__20543),
            .DOUT(N__20542),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__20544),
            .PADOUT(N__20543),
            .PADIN(N__20542),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__20535),
            .DIN(N__20534),
            .DOUT(N__20533),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__20535),
            .PADOUT(N__20534),
            .PADIN(N__20533),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__20526),
            .DIN(N__20525),
            .DOUT(N__20524),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__20526),
            .PADOUT(N__20525),
            .PADIN(N__20524),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__20517),
            .DIN(N__20516),
            .DOUT(N__20515),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__20517),
            .PADOUT(N__20516),
            .PADIN(N__20515),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__20508),
            .DIN(N__20507),
            .DOUT(N__20506),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__20508),
            .PADOUT(N__20507),
            .PADIN(N__20506),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7217),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__20499),
            .DIN(N__20498),
            .DOUT(N__20497),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__20499),
            .PADOUT(N__20498),
            .PADIN(N__20497),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__18689),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__20490),
            .DIN(N__20489),
            .DOUT(N__20488),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__20490),
            .PADOUT(N__20489),
            .PADIN(N__20488),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__20481),
            .DIN(N__20480),
            .DOUT(N__20479),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__20481),
            .PADOUT(N__20480),
            .PADIN(N__20479),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7802),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_ibuf_iopad (
            .OE(N__20472),
            .DIN(N__20471),
            .DOUT(N__20470),
            .PACKAGEPIN(port_rw));
    defparam port_rw_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_rw_ibuf_preio (
            .PADOEN(N__20472),
            .PADOUT(N__20471),
            .PADIN(N__20470),
            .CLOCKENABLE(),
            .DIN0(port_rw_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__20463),
            .DIN(N__20462),
            .DOUT(N__20461),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__20463),
            .PADOUT(N__20462),
            .PADIN(N__20461),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__9050),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__20454),
            .DIN(N__20453),
            .DOUT(N__20452),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__20454),
            .PADOUT(N__20453),
            .PADIN(N__20452),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__9040),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__20445),
            .DIN(N__20444),
            .DOUT(N__20443),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__20445),
            .PADOUT(N__20444),
            .PADIN(N__20443),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12088),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__20436),
            .DIN(N__20435),
            .DOUT(N__20434),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__20436),
            .PADOUT(N__20435),
            .PADIN(N__20434),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12098),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__20427),
            .DIN(N__20426),
            .DOUT(N__20425),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__20427),
            .PADOUT(N__20426),
            .PADIN(N__20425),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8707),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__20418),
            .DIN(N__20417),
            .DOUT(N__20416),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__20418),
            .PADOUT(N__20417),
            .PADIN(N__20416),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8714),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__20409),
            .DIN(N__20408),
            .DOUT(N__20407),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__20409),
            .PADOUT(N__20408),
            .PADIN(N__20407),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__20400),
            .DIN(N__20399),
            .DOUT(N__20398),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__20400),
            .PADOUT(N__20399),
            .PADIN(N__20398),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7211),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__20391),
            .DIN(N__20390),
            .DOUT(N__20389),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__20391),
            .PADOUT(N__20390),
            .PADIN(N__20389),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__9515),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__4905 (
            .O(N__20372),
            .I(N__20369));
    InMux I__4904 (
            .O(N__20369),
            .I(N__20365));
    CascadeMux I__4903 (
            .O(N__20368),
            .I(N__20362));
    LocalMux I__4902 (
            .O(N__20365),
            .I(N__20359));
    InMux I__4901 (
            .O(N__20362),
            .I(N__20356));
    Span4Mux_v I__4900 (
            .O(N__20359),
            .I(N__20353));
    LocalMux I__4899 (
            .O(N__20356),
            .I(N__20350));
    Span4Mux_v I__4898 (
            .O(N__20353),
            .I(N__20344));
    Span4Mux_v I__4897 (
            .O(N__20350),
            .I(N__20344));
    InMux I__4896 (
            .O(N__20349),
            .I(N__20341));
    Sp12to4 I__4895 (
            .O(N__20344),
            .I(N__20336));
    LocalMux I__4894 (
            .O(N__20341),
            .I(N__20336));
    Span12Mux_h I__4893 (
            .O(N__20336),
            .I(N__20333));
    Odrv12 I__4892 (
            .O(N__20333),
            .I(port_data_c_3));
    InMux I__4891 (
            .O(N__20330),
            .I(N__20321));
    InMux I__4890 (
            .O(N__20329),
            .I(N__20321));
    InMux I__4889 (
            .O(N__20328),
            .I(N__20314));
    InMux I__4888 (
            .O(N__20327),
            .I(N__20310));
    InMux I__4887 (
            .O(N__20326),
            .I(N__20307));
    LocalMux I__4886 (
            .O(N__20321),
            .I(N__20304));
    InMux I__4885 (
            .O(N__20320),
            .I(N__20301));
    InMux I__4884 (
            .O(N__20319),
            .I(N__20298));
    InMux I__4883 (
            .O(N__20318),
            .I(N__20295));
    InMux I__4882 (
            .O(N__20317),
            .I(N__20292));
    LocalMux I__4881 (
            .O(N__20314),
            .I(N__20289));
    InMux I__4880 (
            .O(N__20313),
            .I(N__20286));
    LocalMux I__4879 (
            .O(N__20310),
            .I(N__20281));
    LocalMux I__4878 (
            .O(N__20307),
            .I(N__20278));
    Span4Mux_v I__4877 (
            .O(N__20304),
            .I(N__20273));
    LocalMux I__4876 (
            .O(N__20301),
            .I(N__20273));
    LocalMux I__4875 (
            .O(N__20298),
            .I(N__20262));
    LocalMux I__4874 (
            .O(N__20295),
            .I(N__20262));
    LocalMux I__4873 (
            .O(N__20292),
            .I(N__20262));
    Span4Mux_v I__4872 (
            .O(N__20289),
            .I(N__20262));
    LocalMux I__4871 (
            .O(N__20286),
            .I(N__20262));
    InMux I__4870 (
            .O(N__20285),
            .I(N__20259));
    InMux I__4869 (
            .O(N__20284),
            .I(N__20256));
    Span4Mux_v I__4868 (
            .O(N__20281),
            .I(N__20253));
    Span4Mux_h I__4867 (
            .O(N__20278),
            .I(N__20250));
    Span4Mux_v I__4866 (
            .O(N__20273),
            .I(N__20245));
    Span4Mux_v I__4865 (
            .O(N__20262),
            .I(N__20245));
    LocalMux I__4864 (
            .O(N__20259),
            .I(N__20242));
    LocalMux I__4863 (
            .O(N__20256),
            .I(N__20239));
    Odrv4 I__4862 (
            .O(N__20253),
            .I(M_this_vram_write_en_0_sqmuxa));
    Odrv4 I__4861 (
            .O(N__20250),
            .I(M_this_vram_write_en_0_sqmuxa));
    Odrv4 I__4860 (
            .O(N__20245),
            .I(M_this_vram_write_en_0_sqmuxa));
    Odrv12 I__4859 (
            .O(N__20242),
            .I(M_this_vram_write_en_0_sqmuxa));
    Odrv4 I__4858 (
            .O(N__20239),
            .I(M_this_vram_write_en_0_sqmuxa));
    InMux I__4857 (
            .O(N__20228),
            .I(N__20225));
    LocalMux I__4856 (
            .O(N__20225),
            .I(N__20221));
    InMux I__4855 (
            .O(N__20224),
            .I(N__20218));
    Span4Mux_v I__4854 (
            .O(N__20221),
            .I(N__20212));
    LocalMux I__4853 (
            .O(N__20218),
            .I(N__20212));
    InMux I__4852 (
            .O(N__20217),
            .I(N__20209));
    Span4Mux_v I__4851 (
            .O(N__20212),
            .I(N__20203));
    LocalMux I__4850 (
            .O(N__20209),
            .I(N__20203));
    InMux I__4849 (
            .O(N__20208),
            .I(N__20200));
    Span4Mux_v I__4848 (
            .O(N__20203),
            .I(N__20194));
    LocalMux I__4847 (
            .O(N__20200),
            .I(N__20194));
    InMux I__4846 (
            .O(N__20199),
            .I(N__20191));
    Span4Mux_v I__4845 (
            .O(N__20194),
            .I(N__20184));
    LocalMux I__4844 (
            .O(N__20191),
            .I(N__20184));
    InMux I__4843 (
            .O(N__20190),
            .I(N__20181));
    InMux I__4842 (
            .O(N__20189),
            .I(N__20178));
    Span4Mux_v I__4841 (
            .O(N__20184),
            .I(N__20175));
    LocalMux I__4840 (
            .O(N__20181),
            .I(N__20172));
    LocalMux I__4839 (
            .O(N__20178),
            .I(N__20169));
    Span4Mux_v I__4838 (
            .O(N__20175),
            .I(N__20163));
    Span4Mux_s2_v I__4837 (
            .O(N__20172),
            .I(N__20163));
    Span4Mux_h I__4836 (
            .O(N__20169),
            .I(N__20160));
    InMux I__4835 (
            .O(N__20168),
            .I(N__20157));
    Odrv4 I__4834 (
            .O(N__20163),
            .I(M_this_vram_write_data_3));
    Odrv4 I__4833 (
            .O(N__20160),
            .I(M_this_vram_write_data_3));
    LocalMux I__4832 (
            .O(N__20157),
            .I(M_this_vram_write_data_3));
    InMux I__4831 (
            .O(N__20150),
            .I(N__20147));
    LocalMux I__4830 (
            .O(N__20147),
            .I(N__20144));
    Span12Mux_s10_h I__4829 (
            .O(N__20144),
            .I(N__20141));
    Span12Mux_v I__4828 (
            .O(N__20141),
            .I(N__20138));
    Odrv12 I__4827 (
            .O(N__20138),
            .I(\this_vga_signals.g0_7 ));
    InMux I__4826 (
            .O(N__20135),
            .I(N__20132));
    LocalMux I__4825 (
            .O(N__20132),
            .I(N__20129));
    Span12Mux_h I__4824 (
            .O(N__20129),
            .I(N__20126));
    Span12Mux_v I__4823 (
            .O(N__20126),
            .I(N__20123));
    Odrv12 I__4822 (
            .O(N__20123),
            .I(\this_vga_signals.mult1_un89_sum_c5 ));
    CascadeMux I__4821 (
            .O(N__20120),
            .I(N__20117));
    CascadeBuf I__4820 (
            .O(N__20117),
            .I(N__20114));
    CascadeMux I__4819 (
            .O(N__20114),
            .I(N__20111));
    CascadeBuf I__4818 (
            .O(N__20111),
            .I(N__20108));
    CascadeMux I__4817 (
            .O(N__20108),
            .I(N__20105));
    CascadeBuf I__4816 (
            .O(N__20105),
            .I(N__20102));
    CascadeMux I__4815 (
            .O(N__20102),
            .I(N__20099));
    CascadeBuf I__4814 (
            .O(N__20099),
            .I(N__20096));
    CascadeMux I__4813 (
            .O(N__20096),
            .I(N__20093));
    CascadeBuf I__4812 (
            .O(N__20093),
            .I(N__20090));
    CascadeMux I__4811 (
            .O(N__20090),
            .I(N__20087));
    CascadeBuf I__4810 (
            .O(N__20087),
            .I(N__20084));
    CascadeMux I__4809 (
            .O(N__20084),
            .I(N__20081));
    CascadeBuf I__4808 (
            .O(N__20081),
            .I(N__20078));
    CascadeMux I__4807 (
            .O(N__20078),
            .I(N__20075));
    CascadeBuf I__4806 (
            .O(N__20075),
            .I(N__20072));
    CascadeMux I__4805 (
            .O(N__20072),
            .I(N__20069));
    CascadeBuf I__4804 (
            .O(N__20069),
            .I(N__20066));
    CascadeMux I__4803 (
            .O(N__20066),
            .I(N__20063));
    CascadeBuf I__4802 (
            .O(N__20063),
            .I(N__20060));
    CascadeMux I__4801 (
            .O(N__20060),
            .I(N__20057));
    CascadeBuf I__4800 (
            .O(N__20057),
            .I(N__20054));
    CascadeMux I__4799 (
            .O(N__20054),
            .I(N__20051));
    CascadeBuf I__4798 (
            .O(N__20051),
            .I(N__20048));
    CascadeMux I__4797 (
            .O(N__20048),
            .I(N__20045));
    CascadeBuf I__4796 (
            .O(N__20045),
            .I(N__20042));
    CascadeMux I__4795 (
            .O(N__20042),
            .I(N__20039));
    CascadeBuf I__4794 (
            .O(N__20039),
            .I(N__20036));
    CascadeMux I__4793 (
            .O(N__20036),
            .I(N__20033));
    CascadeBuf I__4792 (
            .O(N__20033),
            .I(N__20030));
    CascadeMux I__4791 (
            .O(N__20030),
            .I(N__20027));
    InMux I__4790 (
            .O(N__20027),
            .I(N__20024));
    LocalMux I__4789 (
            .O(N__20024),
            .I(M_this_vga_signals_address_1));
    InMux I__4788 (
            .O(N__20021),
            .I(N__20016));
    CascadeMux I__4787 (
            .O(N__20020),
            .I(N__20013));
    InMux I__4786 (
            .O(N__20019),
            .I(N__20009));
    LocalMux I__4785 (
            .O(N__20016),
            .I(N__20003));
    InMux I__4784 (
            .O(N__20013),
            .I(N__20000));
    CascadeMux I__4783 (
            .O(N__20012),
            .I(N__19996));
    LocalMux I__4782 (
            .O(N__20009),
            .I(N__19990));
    InMux I__4781 (
            .O(N__20008),
            .I(N__19987));
    InMux I__4780 (
            .O(N__20007),
            .I(N__19982));
    InMux I__4779 (
            .O(N__20006),
            .I(N__19979));
    Span4Mux_v I__4778 (
            .O(N__20003),
            .I(N__19976));
    LocalMux I__4777 (
            .O(N__20000),
            .I(N__19973));
    InMux I__4776 (
            .O(N__19999),
            .I(N__19970));
    InMux I__4775 (
            .O(N__19996),
            .I(N__19967));
    InMux I__4774 (
            .O(N__19995),
            .I(N__19964));
    InMux I__4773 (
            .O(N__19994),
            .I(N__19961));
    InMux I__4772 (
            .O(N__19993),
            .I(N__19958));
    Span4Mux_h I__4771 (
            .O(N__19990),
            .I(N__19953));
    LocalMux I__4770 (
            .O(N__19987),
            .I(N__19953));
    InMux I__4769 (
            .O(N__19986),
            .I(N__19950));
    CascadeMux I__4768 (
            .O(N__19985),
            .I(N__19947));
    LocalMux I__4767 (
            .O(N__19982),
            .I(N__19943));
    LocalMux I__4766 (
            .O(N__19979),
            .I(N__19940));
    Sp12to4 I__4765 (
            .O(N__19976),
            .I(N__19937));
    Span4Mux_h I__4764 (
            .O(N__19973),
            .I(N__19934));
    LocalMux I__4763 (
            .O(N__19970),
            .I(N__19931));
    LocalMux I__4762 (
            .O(N__19967),
            .I(N__19928));
    LocalMux I__4761 (
            .O(N__19964),
            .I(N__19917));
    LocalMux I__4760 (
            .O(N__19961),
            .I(N__19917));
    LocalMux I__4759 (
            .O(N__19958),
            .I(N__19917));
    Span4Mux_h I__4758 (
            .O(N__19953),
            .I(N__19917));
    LocalMux I__4757 (
            .O(N__19950),
            .I(N__19917));
    InMux I__4756 (
            .O(N__19947),
            .I(N__19914));
    InMux I__4755 (
            .O(N__19946),
            .I(N__19911));
    Span12Mux_v I__4754 (
            .O(N__19943),
            .I(N__19908));
    Span4Mux_v I__4753 (
            .O(N__19940),
            .I(N__19905));
    Span12Mux_h I__4752 (
            .O(N__19937),
            .I(N__19902));
    Sp12to4 I__4751 (
            .O(N__19934),
            .I(N__19899));
    Span4Mux_h I__4750 (
            .O(N__19931),
            .I(N__19890));
    Span4Mux_h I__4749 (
            .O(N__19928),
            .I(N__19890));
    Span4Mux_v I__4748 (
            .O(N__19917),
            .I(N__19890));
    LocalMux I__4747 (
            .O(N__19914),
            .I(N__19890));
    LocalMux I__4746 (
            .O(N__19911),
            .I(N__19887));
    Span12Mux_h I__4745 (
            .O(N__19908),
            .I(N__19884));
    Sp12to4 I__4744 (
            .O(N__19905),
            .I(N__19877));
    Span12Mux_v I__4743 (
            .O(N__19902),
            .I(N__19877));
    Span12Mux_v I__4742 (
            .O(N__19899),
            .I(N__19877));
    Span4Mux_h I__4741 (
            .O(N__19890),
            .I(N__19874));
    Odrv4 I__4740 (
            .O(N__19887),
            .I(\this_vga_signals.rgb72 ));
    Odrv12 I__4739 (
            .O(N__19884),
            .I(\this_vga_signals.rgb72 ));
    Odrv12 I__4738 (
            .O(N__19877),
            .I(\this_vga_signals.rgb72 ));
    Odrv4 I__4737 (
            .O(N__19874),
            .I(\this_vga_signals.rgb72 ));
    InMux I__4736 (
            .O(N__19865),
            .I(N__19861));
    InMux I__4735 (
            .O(N__19864),
            .I(N__19858));
    LocalMux I__4734 (
            .O(N__19861),
            .I(N__19855));
    LocalMux I__4733 (
            .O(N__19858),
            .I(N__19852));
    Span12Mux_s7_v I__4732 (
            .O(N__19855),
            .I(N__19849));
    Span12Mux_h I__4731 (
            .O(N__19852),
            .I(N__19846));
    Span12Mux_h I__4730 (
            .O(N__19849),
            .I(N__19843));
    Span12Mux_v I__4729 (
            .O(N__19846),
            .I(N__19840));
    Odrv12 I__4728 (
            .O(N__19843),
            .I(\this_vga_signals.mult1_un82_sum_c5 ));
    Odrv12 I__4727 (
            .O(N__19840),
            .I(\this_vga_signals.mult1_un82_sum_c5 ));
    InMux I__4726 (
            .O(N__19835),
            .I(N__19832));
    LocalMux I__4725 (
            .O(N__19832),
            .I(N__19829));
    Span12Mux_s10_v I__4724 (
            .O(N__19829),
            .I(N__19826));
    Span12Mux_h I__4723 (
            .O(N__19826),
            .I(N__19822));
    InMux I__4722 (
            .O(N__19825),
            .I(N__19819));
    Odrv12 I__4721 (
            .O(N__19822),
            .I(\this_vga_signals.mult1_un82_sum_axbxc5_1_i ));
    LocalMux I__4720 (
            .O(N__19819),
            .I(\this_vga_signals.mult1_un82_sum_axbxc5_1_i ));
    CascadeMux I__4719 (
            .O(N__19814),
            .I(N__19811));
    CascadeBuf I__4718 (
            .O(N__19811),
            .I(N__19808));
    CascadeMux I__4717 (
            .O(N__19808),
            .I(N__19805));
    CascadeBuf I__4716 (
            .O(N__19805),
            .I(N__19802));
    CascadeMux I__4715 (
            .O(N__19802),
            .I(N__19799));
    CascadeBuf I__4714 (
            .O(N__19799),
            .I(N__19796));
    CascadeMux I__4713 (
            .O(N__19796),
            .I(N__19793));
    CascadeBuf I__4712 (
            .O(N__19793),
            .I(N__19790));
    CascadeMux I__4711 (
            .O(N__19790),
            .I(N__19787));
    CascadeBuf I__4710 (
            .O(N__19787),
            .I(N__19784));
    CascadeMux I__4709 (
            .O(N__19784),
            .I(N__19781));
    CascadeBuf I__4708 (
            .O(N__19781),
            .I(N__19778));
    CascadeMux I__4707 (
            .O(N__19778),
            .I(N__19775));
    CascadeBuf I__4706 (
            .O(N__19775),
            .I(N__19772));
    CascadeMux I__4705 (
            .O(N__19772),
            .I(N__19769));
    CascadeBuf I__4704 (
            .O(N__19769),
            .I(N__19766));
    CascadeMux I__4703 (
            .O(N__19766),
            .I(N__19763));
    CascadeBuf I__4702 (
            .O(N__19763),
            .I(N__19760));
    CascadeMux I__4701 (
            .O(N__19760),
            .I(N__19757));
    CascadeBuf I__4700 (
            .O(N__19757),
            .I(N__19754));
    CascadeMux I__4699 (
            .O(N__19754),
            .I(N__19751));
    CascadeBuf I__4698 (
            .O(N__19751),
            .I(N__19748));
    CascadeMux I__4697 (
            .O(N__19748),
            .I(N__19745));
    CascadeBuf I__4696 (
            .O(N__19745),
            .I(N__19742));
    CascadeMux I__4695 (
            .O(N__19742),
            .I(N__19739));
    CascadeBuf I__4694 (
            .O(N__19739),
            .I(N__19736));
    CascadeMux I__4693 (
            .O(N__19736),
            .I(N__19733));
    CascadeBuf I__4692 (
            .O(N__19733),
            .I(N__19730));
    CascadeMux I__4691 (
            .O(N__19730),
            .I(N__19727));
    CascadeBuf I__4690 (
            .O(N__19727),
            .I(N__19724));
    CascadeMux I__4689 (
            .O(N__19724),
            .I(N__19721));
    InMux I__4688 (
            .O(N__19721),
            .I(N__19718));
    LocalMux I__4687 (
            .O(N__19718),
            .I(M_this_vga_signals_address_2));
    InMux I__4686 (
            .O(N__19715),
            .I(N__19712));
    LocalMux I__4685 (
            .O(N__19712),
            .I(N__19709));
    Span12Mux_s10_h I__4684 (
            .O(N__19709),
            .I(N__19706));
    Span12Mux_h I__4683 (
            .O(N__19706),
            .I(N__19702));
    InMux I__4682 (
            .O(N__19705),
            .I(N__19699));
    Odrv12 I__4681 (
            .O(N__19702),
            .I(port_rw_c));
    LocalMux I__4680 (
            .O(N__19699),
            .I(port_rw_c));
    InMux I__4679 (
            .O(N__19694),
            .I(N__19691));
    LocalMux I__4678 (
            .O(N__19691),
            .I(N__19688));
    Span12Mux_v I__4677 (
            .O(N__19688),
            .I(N__19685));
    Odrv12 I__4676 (
            .O(N__19685),
            .I(port_address_c_6));
    CascadeMux I__4675 (
            .O(N__19682),
            .I(N__19679));
    InMux I__4674 (
            .O(N__19679),
            .I(N__19676));
    LocalMux I__4673 (
            .O(N__19676),
            .I(port_address_c_5));
    InMux I__4672 (
            .O(N__19673),
            .I(N__19670));
    LocalMux I__4671 (
            .O(N__19670),
            .I(N__19667));
    Span12Mux_v I__4670 (
            .O(N__19667),
            .I(N__19664));
    Odrv12 I__4669 (
            .O(N__19664),
            .I(port_address_c_3));
    InMux I__4668 (
            .O(N__19661),
            .I(N__19658));
    LocalMux I__4667 (
            .O(N__19658),
            .I(N__19655));
    Span4Mux_h I__4666 (
            .O(N__19655),
            .I(N__19652));
    Span4Mux_h I__4665 (
            .O(N__19652),
            .I(N__19649));
    Span4Mux_h I__4664 (
            .O(N__19649),
            .I(N__19646));
    Odrv4 I__4663 (
            .O(N__19646),
            .I(M_state_q_ns_1_0__m7Z0Z_4));
    InMux I__4662 (
            .O(N__19643),
            .I(N__19640));
    LocalMux I__4661 (
            .O(N__19640),
            .I(\this_vram.mem_mem_2_1_RNI01NZ0Z11 ));
    CascadeMux I__4660 (
            .O(N__19637),
            .I(\this_vram.mem_mem_0_1_RNISOIZ0Z11_cascade_ ));
    InMux I__4659 (
            .O(N__19634),
            .I(N__19629));
    InMux I__4658 (
            .O(N__19633),
            .I(N__19626));
    InMux I__4657 (
            .O(N__19632),
            .I(N__19623));
    LocalMux I__4656 (
            .O(N__19629),
            .I(N__19614));
    LocalMux I__4655 (
            .O(N__19626),
            .I(N__19614));
    LocalMux I__4654 (
            .O(N__19623),
            .I(N__19611));
    InMux I__4653 (
            .O(N__19622),
            .I(N__19607));
    InMux I__4652 (
            .O(N__19621),
            .I(N__19604));
    InMux I__4651 (
            .O(N__19620),
            .I(N__19601));
    InMux I__4650 (
            .O(N__19619),
            .I(N__19598));
    Span4Mux_v I__4649 (
            .O(N__19614),
            .I(N__19593));
    Span4Mux_v I__4648 (
            .O(N__19611),
            .I(N__19593));
    InMux I__4647 (
            .O(N__19610),
            .I(N__19590));
    LocalMux I__4646 (
            .O(N__19607),
            .I(N__19585));
    LocalMux I__4645 (
            .O(N__19604),
            .I(N__19585));
    LocalMux I__4644 (
            .O(N__19601),
            .I(N__19576));
    LocalMux I__4643 (
            .O(N__19598),
            .I(N__19576));
    Sp12to4 I__4642 (
            .O(N__19593),
            .I(N__19576));
    LocalMux I__4641 (
            .O(N__19590),
            .I(N__19576));
    Sp12to4 I__4640 (
            .O(N__19585),
            .I(N__19573));
    Span12Mux_h I__4639 (
            .O(N__19576),
            .I(N__19570));
    Span12Mux_v I__4638 (
            .O(N__19573),
            .I(N__19567));
    Odrv12 I__4637 (
            .O(N__19570),
            .I(\this_vram.mem_radregZ0Z_12 ));
    Odrv12 I__4636 (
            .O(N__19567),
            .I(\this_vram.mem_radregZ0Z_12 ));
    InMux I__4635 (
            .O(N__19562),
            .I(N__19559));
    LocalMux I__4634 (
            .O(N__19559),
            .I(\this_vram.mem_N_98 ));
    InMux I__4633 (
            .O(N__19556),
            .I(N__19553));
    LocalMux I__4632 (
            .O(N__19553),
            .I(N__19550));
    Span12Mux_h I__4631 (
            .O(N__19550),
            .I(N__19547));
    Span12Mux_v I__4630 (
            .O(N__19547),
            .I(N__19544));
    Odrv12 I__4629 (
            .O(N__19544),
            .I(\this_vram.mem_out_bus1_0 ));
    InMux I__4628 (
            .O(N__19541),
            .I(N__19538));
    LocalMux I__4627 (
            .O(N__19538),
            .I(N__19535));
    Span4Mux_v I__4626 (
            .O(N__19535),
            .I(N__19532));
    Odrv4 I__4625 (
            .O(N__19532),
            .I(\this_vram.mem_out_bus5_0 ));
    InMux I__4624 (
            .O(N__19529),
            .I(N__19526));
    LocalMux I__4623 (
            .O(N__19526),
            .I(\this_vram.mem_mem_1_0_RNISSKZ0Z11 ));
    InMux I__4622 (
            .O(N__19523),
            .I(N__19504));
    InMux I__4621 (
            .O(N__19522),
            .I(N__19504));
    InMux I__4620 (
            .O(N__19521),
            .I(N__19504));
    InMux I__4619 (
            .O(N__19520),
            .I(N__19504));
    InMux I__4618 (
            .O(N__19519),
            .I(N__19497));
    InMux I__4617 (
            .O(N__19518),
            .I(N__19497));
    InMux I__4616 (
            .O(N__19517),
            .I(N__19497));
    InMux I__4615 (
            .O(N__19516),
            .I(N__19494));
    InMux I__4614 (
            .O(N__19515),
            .I(N__19491));
    InMux I__4613 (
            .O(N__19514),
            .I(N__19486));
    InMux I__4612 (
            .O(N__19513),
            .I(N__19486));
    LocalMux I__4611 (
            .O(N__19504),
            .I(N__19475));
    LocalMux I__4610 (
            .O(N__19497),
            .I(N__19475));
    LocalMux I__4609 (
            .O(N__19494),
            .I(N__19475));
    LocalMux I__4608 (
            .O(N__19491),
            .I(N__19475));
    LocalMux I__4607 (
            .O(N__19486),
            .I(N__19475));
    Span4Mux_v I__4606 (
            .O(N__19475),
            .I(N__19467));
    InMux I__4605 (
            .O(N__19474),
            .I(N__19464));
    InMux I__4604 (
            .O(N__19473),
            .I(N__19457));
    InMux I__4603 (
            .O(N__19472),
            .I(N__19457));
    InMux I__4602 (
            .O(N__19471),
            .I(N__19457));
    InMux I__4601 (
            .O(N__19470),
            .I(N__19454));
    Sp12to4 I__4600 (
            .O(N__19467),
            .I(N__19445));
    LocalMux I__4599 (
            .O(N__19464),
            .I(N__19445));
    LocalMux I__4598 (
            .O(N__19457),
            .I(N__19445));
    LocalMux I__4597 (
            .O(N__19454),
            .I(N__19445));
    Span12Mux_h I__4596 (
            .O(N__19445),
            .I(N__19442));
    Odrv12 I__4595 (
            .O(N__19442),
            .I(\this_vram.mem_radregZ0Z_13 ));
    InMux I__4594 (
            .O(N__19439),
            .I(N__19436));
    LocalMux I__4593 (
            .O(N__19436),
            .I(N__19433));
    Span4Mux_v I__4592 (
            .O(N__19433),
            .I(N__19430));
    Span4Mux_v I__4591 (
            .O(N__19430),
            .I(N__19427));
    Odrv4 I__4590 (
            .O(N__19427),
            .I(\this_vram.mem_out_bus7_1 ));
    InMux I__4589 (
            .O(N__19424),
            .I(N__19421));
    LocalMux I__4588 (
            .O(N__19421),
            .I(N__19418));
    Span4Mux_v I__4587 (
            .O(N__19418),
            .I(N__19415));
    Odrv4 I__4586 (
            .O(N__19415),
            .I(\this_vram.mem_out_bus3_1 ));
    InMux I__4585 (
            .O(N__19412),
            .I(N__19409));
    LocalMux I__4584 (
            .O(N__19409),
            .I(N__19406));
    Odrv4 I__4583 (
            .O(N__19406),
            .I(\this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ));
    CEMux I__4582 (
            .O(N__19403),
            .I(N__19400));
    LocalMux I__4581 (
            .O(N__19400),
            .I(N__19396));
    CEMux I__4580 (
            .O(N__19399),
            .I(N__19393));
    Span4Mux_v I__4579 (
            .O(N__19396),
            .I(N__19390));
    LocalMux I__4578 (
            .O(N__19393),
            .I(N__19387));
    Span4Mux_h I__4577 (
            .O(N__19390),
            .I(N__19384));
    Span4Mux_h I__4576 (
            .O(N__19387),
            .I(N__19381));
    Odrv4 I__4575 (
            .O(N__19384),
            .I(\this_vram.mem_WE_6 ));
    Odrv4 I__4574 (
            .O(N__19381),
            .I(\this_vram.mem_WE_6 ));
    CEMux I__4573 (
            .O(N__19376),
            .I(N__19373));
    LocalMux I__4572 (
            .O(N__19373),
            .I(N__19369));
    CEMux I__4571 (
            .O(N__19372),
            .I(N__19366));
    Span4Mux_v I__4570 (
            .O(N__19369),
            .I(N__19363));
    LocalMux I__4569 (
            .O(N__19366),
            .I(N__19360));
    Span4Mux_h I__4568 (
            .O(N__19363),
            .I(N__19357));
    Span4Mux_h I__4567 (
            .O(N__19360),
            .I(N__19354));
    Odrv4 I__4566 (
            .O(N__19357),
            .I(\this_vram.mem_WE_4 ));
    Odrv4 I__4565 (
            .O(N__19354),
            .I(\this_vram.mem_WE_4 ));
    CEMux I__4564 (
            .O(N__19349),
            .I(N__19345));
    CEMux I__4563 (
            .O(N__19348),
            .I(N__19342));
    LocalMux I__4562 (
            .O(N__19345),
            .I(N__19339));
    LocalMux I__4561 (
            .O(N__19342),
            .I(N__19336));
    Span4Mux_v I__4560 (
            .O(N__19339),
            .I(N__19333));
    Span4Mux_h I__4559 (
            .O(N__19336),
            .I(N__19330));
    Odrv4 I__4558 (
            .O(N__19333),
            .I(\this_vram.mem_WE_2 ));
    Odrv4 I__4557 (
            .O(N__19330),
            .I(\this_vram.mem_WE_2 ));
    InMux I__4556 (
            .O(N__19325),
            .I(N__19319));
    InMux I__4555 (
            .O(N__19324),
            .I(N__19319));
    LocalMux I__4554 (
            .O(N__19319),
            .I(N__19312));
    InMux I__4553 (
            .O(N__19318),
            .I(N__19309));
    InMux I__4552 (
            .O(N__19317),
            .I(N__19304));
    InMux I__4551 (
            .O(N__19316),
            .I(N__19301));
    InMux I__4550 (
            .O(N__19315),
            .I(N__19298));
    Span4Mux_h I__4549 (
            .O(N__19312),
            .I(N__19293));
    LocalMux I__4548 (
            .O(N__19309),
            .I(N__19293));
    InMux I__4547 (
            .O(N__19308),
            .I(N__19290));
    InMux I__4546 (
            .O(N__19307),
            .I(N__19287));
    LocalMux I__4545 (
            .O(N__19304),
            .I(N__19279));
    LocalMux I__4544 (
            .O(N__19301),
            .I(N__19279));
    LocalMux I__4543 (
            .O(N__19298),
            .I(N__19279));
    Span4Mux_h I__4542 (
            .O(N__19293),
            .I(N__19274));
    LocalMux I__4541 (
            .O(N__19290),
            .I(N__19274));
    LocalMux I__4540 (
            .O(N__19287),
            .I(N__19270));
    InMux I__4539 (
            .O(N__19286),
            .I(N__19267));
    Span12Mux_v I__4538 (
            .O(N__19279),
            .I(N__19264));
    Span4Mux_v I__4537 (
            .O(N__19274),
            .I(N__19261));
    InMux I__4536 (
            .O(N__19273),
            .I(N__19258));
    Span12Mux_h I__4535 (
            .O(N__19270),
            .I(N__19253));
    LocalMux I__4534 (
            .O(N__19267),
            .I(N__19253));
    Odrv12 I__4533 (
            .O(N__19264),
            .I(M_current_address_qZ0Z_12));
    Odrv4 I__4532 (
            .O(N__19261),
            .I(M_current_address_qZ0Z_12));
    LocalMux I__4531 (
            .O(N__19258),
            .I(M_current_address_qZ0Z_12));
    Odrv12 I__4530 (
            .O(N__19253),
            .I(M_current_address_qZ0Z_12));
    CascadeMux I__4529 (
            .O(N__19244),
            .I(N__19240));
    InMux I__4528 (
            .O(N__19243),
            .I(N__19234));
    InMux I__4527 (
            .O(N__19240),
            .I(N__19229));
    InMux I__4526 (
            .O(N__19239),
            .I(N__19229));
    InMux I__4525 (
            .O(N__19238),
            .I(N__19226));
    InMux I__4524 (
            .O(N__19237),
            .I(N__19223));
    LocalMux I__4523 (
            .O(N__19234),
            .I(N__19218));
    LocalMux I__4522 (
            .O(N__19229),
            .I(N__19211));
    LocalMux I__4521 (
            .O(N__19226),
            .I(N__19211));
    LocalMux I__4520 (
            .O(N__19223),
            .I(N__19211));
    InMux I__4519 (
            .O(N__19222),
            .I(N__19208));
    InMux I__4518 (
            .O(N__19221),
            .I(N__19205));
    Span4Mux_v I__4517 (
            .O(N__19218),
            .I(N__19200));
    Span4Mux_v I__4516 (
            .O(N__19211),
            .I(N__19197));
    LocalMux I__4515 (
            .O(N__19208),
            .I(N__19192));
    LocalMux I__4514 (
            .O(N__19205),
            .I(N__19192));
    InMux I__4513 (
            .O(N__19204),
            .I(N__19189));
    InMux I__4512 (
            .O(N__19203),
            .I(N__19186));
    Span4Mux_v I__4511 (
            .O(N__19200),
            .I(N__19182));
    Span4Mux_v I__4510 (
            .O(N__19197),
            .I(N__19177));
    Span4Mux_v I__4509 (
            .O(N__19192),
            .I(N__19177));
    LocalMux I__4508 (
            .O(N__19189),
            .I(N__19174));
    LocalMux I__4507 (
            .O(N__19186),
            .I(N__19171));
    InMux I__4506 (
            .O(N__19185),
            .I(N__19168));
    Odrv4 I__4505 (
            .O(N__19182),
            .I(M_current_address_qZ0Z_11));
    Odrv4 I__4504 (
            .O(N__19177),
            .I(M_current_address_qZ0Z_11));
    Odrv12 I__4503 (
            .O(N__19174),
            .I(M_current_address_qZ0Z_11));
    Odrv4 I__4502 (
            .O(N__19171),
            .I(M_current_address_qZ0Z_11));
    LocalMux I__4501 (
            .O(N__19168),
            .I(M_current_address_qZ0Z_11));
    CascadeMux I__4500 (
            .O(N__19157),
            .I(N__19152));
    CascadeMux I__4499 (
            .O(N__19156),
            .I(N__19146));
    CascadeMux I__4498 (
            .O(N__19155),
            .I(N__19143));
    InMux I__4497 (
            .O(N__19152),
            .I(N__19139));
    CascadeMux I__4496 (
            .O(N__19151),
            .I(N__19136));
    CascadeMux I__4495 (
            .O(N__19150),
            .I(N__19133));
    InMux I__4494 (
            .O(N__19149),
            .I(N__19128));
    InMux I__4493 (
            .O(N__19146),
            .I(N__19128));
    InMux I__4492 (
            .O(N__19143),
            .I(N__19125));
    CascadeMux I__4491 (
            .O(N__19142),
            .I(N__19122));
    LocalMux I__4490 (
            .O(N__19139),
            .I(N__19119));
    InMux I__4489 (
            .O(N__19136),
            .I(N__19116));
    InMux I__4488 (
            .O(N__19133),
            .I(N__19113));
    LocalMux I__4487 (
            .O(N__19128),
            .I(N__19107));
    LocalMux I__4486 (
            .O(N__19125),
            .I(N__19107));
    InMux I__4485 (
            .O(N__19122),
            .I(N__19104));
    Span4Mux_v I__4484 (
            .O(N__19119),
            .I(N__19097));
    LocalMux I__4483 (
            .O(N__19116),
            .I(N__19097));
    LocalMux I__4482 (
            .O(N__19113),
            .I(N__19097));
    CascadeMux I__4481 (
            .O(N__19112),
            .I(N__19094));
    Sp12to4 I__4480 (
            .O(N__19107),
            .I(N__19089));
    LocalMux I__4479 (
            .O(N__19104),
            .I(N__19089));
    Span4Mux_v I__4478 (
            .O(N__19097),
            .I(N__19086));
    InMux I__4477 (
            .O(N__19094),
            .I(N__19083));
    Span12Mux_v I__4476 (
            .O(N__19089),
            .I(N__19078));
    Sp12to4 I__4475 (
            .O(N__19086),
            .I(N__19073));
    LocalMux I__4474 (
            .O(N__19083),
            .I(N__19073));
    InMux I__4473 (
            .O(N__19082),
            .I(N__19070));
    InMux I__4472 (
            .O(N__19081),
            .I(N__19067));
    Odrv12 I__4471 (
            .O(N__19078),
            .I(M_current_address_qZ0Z_13));
    Odrv12 I__4470 (
            .O(N__19073),
            .I(M_current_address_qZ0Z_13));
    LocalMux I__4469 (
            .O(N__19070),
            .I(M_current_address_qZ0Z_13));
    LocalMux I__4468 (
            .O(N__19067),
            .I(M_current_address_qZ0Z_13));
    CEMux I__4467 (
            .O(N__19058),
            .I(N__19054));
    CEMux I__4466 (
            .O(N__19057),
            .I(N__19051));
    LocalMux I__4465 (
            .O(N__19054),
            .I(N__19046));
    LocalMux I__4464 (
            .O(N__19051),
            .I(N__19046));
    Span4Mux_v I__4463 (
            .O(N__19046),
            .I(N__19043));
    Span4Mux_h I__4462 (
            .O(N__19043),
            .I(N__19040));
    Odrv4 I__4461 (
            .O(N__19040),
            .I(\this_vram.mem_WE_0 ));
    CascadeMux I__4460 (
            .O(N__19037),
            .I(N__19032));
    CascadeMux I__4459 (
            .O(N__19036),
            .I(N__19029));
    InMux I__4458 (
            .O(N__19035),
            .I(N__19026));
    InMux I__4457 (
            .O(N__19032),
            .I(N__19021));
    InMux I__4456 (
            .O(N__19029),
            .I(N__19021));
    LocalMux I__4455 (
            .O(N__19026),
            .I(N__19018));
    LocalMux I__4454 (
            .O(N__19021),
            .I(N__19015));
    Span4Mux_v I__4453 (
            .O(N__19018),
            .I(N__19012));
    Span12Mux_h I__4452 (
            .O(N__19015),
            .I(N__19009));
    IoSpan4Mux I__4451 (
            .O(N__19012),
            .I(N__19006));
    Odrv12 I__4450 (
            .O(N__19009),
            .I(port_data_c_2));
    Odrv4 I__4449 (
            .O(N__19006),
            .I(port_data_c_2));
    InMux I__4448 (
            .O(N__19001),
            .I(N__18998));
    LocalMux I__4447 (
            .O(N__18998),
            .I(N__18993));
    InMux I__4446 (
            .O(N__18997),
            .I(N__18990));
    InMux I__4445 (
            .O(N__18996),
            .I(N__18986));
    Span4Mux_v I__4444 (
            .O(N__18993),
            .I(N__18981));
    LocalMux I__4443 (
            .O(N__18990),
            .I(N__18981));
    InMux I__4442 (
            .O(N__18989),
            .I(N__18978));
    LocalMux I__4441 (
            .O(N__18986),
            .I(N__18973));
    Span4Mux_v I__4440 (
            .O(N__18981),
            .I(N__18968));
    LocalMux I__4439 (
            .O(N__18978),
            .I(N__18968));
    InMux I__4438 (
            .O(N__18977),
            .I(N__18965));
    InMux I__4437 (
            .O(N__18976),
            .I(N__18961));
    Span12Mux_v I__4436 (
            .O(N__18973),
            .I(N__18957));
    Span4Mux_v I__4435 (
            .O(N__18968),
            .I(N__18952));
    LocalMux I__4434 (
            .O(N__18965),
            .I(N__18952));
    InMux I__4433 (
            .O(N__18964),
            .I(N__18949));
    LocalMux I__4432 (
            .O(N__18961),
            .I(N__18946));
    InMux I__4431 (
            .O(N__18960),
            .I(N__18943));
    Span12Mux_v I__4430 (
            .O(N__18957),
            .I(N__18940));
    Span4Mux_v I__4429 (
            .O(N__18952),
            .I(N__18935));
    LocalMux I__4428 (
            .O(N__18949),
            .I(N__18935));
    Span4Mux_s3_v I__4427 (
            .O(N__18946),
            .I(N__18930));
    LocalMux I__4426 (
            .O(N__18943),
            .I(N__18930));
    Odrv12 I__4425 (
            .O(N__18940),
            .I(M_this_vram_write_data_2));
    Odrv4 I__4424 (
            .O(N__18935),
            .I(M_this_vram_write_data_2));
    Odrv4 I__4423 (
            .O(N__18930),
            .I(M_this_vram_write_data_2));
    CascadeMux I__4422 (
            .O(N__18923),
            .I(\this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_ ));
    InMux I__4421 (
            .O(N__18920),
            .I(N__18917));
    LocalMux I__4420 (
            .O(N__18917),
            .I(\this_vram.mem_mem_1_1_RNIUSKZ0Z11 ));
    InMux I__4419 (
            .O(N__18914),
            .I(N__18911));
    LocalMux I__4418 (
            .O(N__18911),
            .I(N__18908));
    Span4Mux_v I__4417 (
            .O(N__18908),
            .I(N__18905));
    Odrv4 I__4416 (
            .O(N__18905),
            .I(\this_vram.mem_N_95 ));
    InMux I__4415 (
            .O(N__18902),
            .I(N__18899));
    LocalMux I__4414 (
            .O(N__18899),
            .I(N__18896));
    Span4Mux_v I__4413 (
            .O(N__18896),
            .I(N__18893));
    Odrv4 I__4412 (
            .O(N__18893),
            .I(\this_vram.mem_out_bus5_3 ));
    InMux I__4411 (
            .O(N__18890),
            .I(N__18887));
    LocalMux I__4410 (
            .O(N__18887),
            .I(N__18884));
    Span4Mux_v I__4409 (
            .O(N__18884),
            .I(N__18881));
    Span4Mux_v I__4408 (
            .O(N__18881),
            .I(N__18878));
    Odrv4 I__4407 (
            .O(N__18878),
            .I(\this_vram.mem_out_bus1_3 ));
    InMux I__4406 (
            .O(N__18875),
            .I(N__18872));
    LocalMux I__4405 (
            .O(N__18872),
            .I(\this_vram.mem_mem_1_1_RNIUSK11Z0Z_0 ));
    InMux I__4404 (
            .O(N__18869),
            .I(N__18866));
    LocalMux I__4403 (
            .O(N__18866),
            .I(N__18863));
    Odrv4 I__4402 (
            .O(N__18863),
            .I(\this_vram.mem_out_bus3_0 ));
    InMux I__4401 (
            .O(N__18860),
            .I(N__18857));
    LocalMux I__4400 (
            .O(N__18857),
            .I(N__18854));
    Sp12to4 I__4399 (
            .O(N__18854),
            .I(N__18851));
    Span12Mux_v I__4398 (
            .O(N__18851),
            .I(N__18848));
    Odrv12 I__4397 (
            .O(N__18848),
            .I(\this_vram.mem_out_bus7_0 ));
    InMux I__4396 (
            .O(N__18845),
            .I(N__18842));
    LocalMux I__4395 (
            .O(N__18842),
            .I(\this_vram.mem_mem_3_0_RNI05PZ0Z11 ));
    InMux I__4394 (
            .O(N__18839),
            .I(N__18836));
    LocalMux I__4393 (
            .O(N__18836),
            .I(N__18833));
    Sp12to4 I__4392 (
            .O(N__18833),
            .I(N__18830));
    Span12Mux_v I__4391 (
            .O(N__18830),
            .I(N__18827));
    Odrv12 I__4390 (
            .O(N__18827),
            .I(\this_vram.mem_out_bus6_3 ));
    InMux I__4389 (
            .O(N__18824),
            .I(N__18821));
    LocalMux I__4388 (
            .O(N__18821),
            .I(N__18818));
    Sp12to4 I__4387 (
            .O(N__18818),
            .I(N__18815));
    Span12Mux_v I__4386 (
            .O(N__18815),
            .I(N__18812));
    Odrv12 I__4385 (
            .O(N__18812),
            .I(\this_vram.mem_out_bus2_3 ));
    CascadeMux I__4384 (
            .O(N__18809),
            .I(\this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_ ));
    InMux I__4383 (
            .O(N__18806),
            .I(N__18803));
    LocalMux I__4382 (
            .O(N__18803),
            .I(\this_vram.mem_N_105 ));
    InMux I__4381 (
            .O(N__18800),
            .I(N__18797));
    LocalMux I__4380 (
            .O(N__18797),
            .I(N__18794));
    Sp12to4 I__4379 (
            .O(N__18794),
            .I(N__18791));
    Span12Mux_v I__4378 (
            .O(N__18791),
            .I(N__18788));
    Odrv12 I__4377 (
            .O(N__18788),
            .I(\this_vram.mem_out_bus0_3 ));
    InMux I__4376 (
            .O(N__18785),
            .I(N__18782));
    LocalMux I__4375 (
            .O(N__18782),
            .I(N__18779));
    Odrv4 I__4374 (
            .O(N__18779),
            .I(\this_vram.mem_out_bus4_3 ));
    InMux I__4373 (
            .O(N__18776),
            .I(N__18773));
    LocalMux I__4372 (
            .O(N__18773),
            .I(\this_vram.mem_mem_0_1_RNISOI11Z0Z_0 ));
    InMux I__4371 (
            .O(N__18770),
            .I(N__18767));
    LocalMux I__4370 (
            .O(N__18767),
            .I(N__18764));
    Span4Mux_h I__4369 (
            .O(N__18764),
            .I(N__18761));
    Span4Mux_v I__4368 (
            .O(N__18761),
            .I(N__18758));
    Odrv4 I__4367 (
            .O(N__18758),
            .I(\this_vram.mem_out_bus2_2 ));
    InMux I__4366 (
            .O(N__18755),
            .I(N__18752));
    LocalMux I__4365 (
            .O(N__18752),
            .I(N__18749));
    Span4Mux_v I__4364 (
            .O(N__18749),
            .I(N__18746));
    Span4Mux_v I__4363 (
            .O(N__18746),
            .I(N__18743));
    Odrv4 I__4362 (
            .O(N__18743),
            .I(\this_vram.mem_out_bus6_2 ));
    InMux I__4361 (
            .O(N__18740),
            .I(N__18737));
    LocalMux I__4360 (
            .O(N__18737),
            .I(N__18734));
    Sp12to4 I__4359 (
            .O(N__18734),
            .I(N__18731));
    Span12Mux_v I__4358 (
            .O(N__18731),
            .I(N__18728));
    Odrv12 I__4357 (
            .O(N__18728),
            .I(\this_vram.mem_out_bus0_2 ));
    InMux I__4356 (
            .O(N__18725),
            .I(N__18722));
    LocalMux I__4355 (
            .O(N__18722),
            .I(N__18719));
    Odrv4 I__4354 (
            .O(N__18719),
            .I(\this_vram.mem_out_bus4_2 ));
    InMux I__4353 (
            .O(N__18716),
            .I(N__18713));
    LocalMux I__4352 (
            .O(N__18713),
            .I(N__18710));
    Span4Mux_v I__4351 (
            .O(N__18710),
            .I(N__18706));
    InMux I__4350 (
            .O(N__18709),
            .I(N__18703));
    Sp12to4 I__4349 (
            .O(N__18706),
            .I(N__18698));
    LocalMux I__4348 (
            .O(N__18703),
            .I(N__18698));
    Odrv12 I__4347 (
            .O(N__18698),
            .I(\this_vram.mem_N_109 ));
    SRMux I__4346 (
            .O(N__18695),
            .I(N__18692));
    LocalMux I__4345 (
            .O(N__18692),
            .I(N__18684));
    SRMux I__4344 (
            .O(N__18691),
            .I(N__18681));
    SRMux I__4343 (
            .O(N__18690),
            .I(N__18678));
    IoInMux I__4342 (
            .O(N__18689),
            .I(N__18674));
    SRMux I__4341 (
            .O(N__18688),
            .I(N__18670));
    SRMux I__4340 (
            .O(N__18687),
            .I(N__18667));
    Span4Mux_s1_v I__4339 (
            .O(N__18684),
            .I(N__18658));
    LocalMux I__4338 (
            .O(N__18681),
            .I(N__18658));
    LocalMux I__4337 (
            .O(N__18678),
            .I(N__18658));
    SRMux I__4336 (
            .O(N__18677),
            .I(N__18655));
    LocalMux I__4335 (
            .O(N__18674),
            .I(N__18651));
    CascadeMux I__4334 (
            .O(N__18673),
            .I(N__18647));
    LocalMux I__4333 (
            .O(N__18670),
            .I(N__18641));
    LocalMux I__4332 (
            .O(N__18667),
            .I(N__18641));
    SRMux I__4331 (
            .O(N__18666),
            .I(N__18638));
    SRMux I__4330 (
            .O(N__18665),
            .I(N__18635));
    Span4Mux_v I__4329 (
            .O(N__18658),
            .I(N__18628));
    LocalMux I__4328 (
            .O(N__18655),
            .I(N__18628));
    SRMux I__4327 (
            .O(N__18654),
            .I(N__18625));
    Span4Mux_s2_h I__4326 (
            .O(N__18651),
            .I(N__18619));
    InMux I__4325 (
            .O(N__18650),
            .I(N__18614));
    InMux I__4324 (
            .O(N__18647),
            .I(N__18614));
    InMux I__4323 (
            .O(N__18646),
            .I(N__18611));
    Span4Mux_v I__4322 (
            .O(N__18641),
            .I(N__18602));
    LocalMux I__4321 (
            .O(N__18638),
            .I(N__18602));
    LocalMux I__4320 (
            .O(N__18635),
            .I(N__18602));
    SRMux I__4319 (
            .O(N__18634),
            .I(N__18599));
    SRMux I__4318 (
            .O(N__18633),
            .I(N__18596));
    Span4Mux_v I__4317 (
            .O(N__18628),
            .I(N__18589));
    LocalMux I__4316 (
            .O(N__18625),
            .I(N__18589));
    SRMux I__4315 (
            .O(N__18624),
            .I(N__18586));
    SRMux I__4314 (
            .O(N__18623),
            .I(N__18583));
    SRMux I__4313 (
            .O(N__18622),
            .I(N__18578));
    Sp12to4 I__4312 (
            .O(N__18619),
            .I(N__18572));
    LocalMux I__4311 (
            .O(N__18614),
            .I(N__18567));
    LocalMux I__4310 (
            .O(N__18611),
            .I(N__18567));
    SRMux I__4309 (
            .O(N__18610),
            .I(N__18564));
    SRMux I__4308 (
            .O(N__18609),
            .I(N__18559));
    Span4Mux_v I__4307 (
            .O(N__18602),
            .I(N__18552));
    LocalMux I__4306 (
            .O(N__18599),
            .I(N__18552));
    LocalMux I__4305 (
            .O(N__18596),
            .I(N__18552));
    SRMux I__4304 (
            .O(N__18595),
            .I(N__18549));
    SRMux I__4303 (
            .O(N__18594),
            .I(N__18546));
    Span4Mux_v I__4302 (
            .O(N__18589),
            .I(N__18541));
    LocalMux I__4301 (
            .O(N__18586),
            .I(N__18541));
    LocalMux I__4300 (
            .O(N__18583),
            .I(N__18538));
    SRMux I__4299 (
            .O(N__18582),
            .I(N__18535));
    SRMux I__4298 (
            .O(N__18581),
            .I(N__18532));
    LocalMux I__4297 (
            .O(N__18578),
            .I(N__18529));
    SRMux I__4296 (
            .O(N__18577),
            .I(N__18526));
    SRMux I__4295 (
            .O(N__18576),
            .I(N__18523));
    SRMux I__4294 (
            .O(N__18575),
            .I(N__18516));
    Span12Mux_s9_v I__4293 (
            .O(N__18572),
            .I(N__18511));
    Span4Mux_h I__4292 (
            .O(N__18567),
            .I(N__18508));
    LocalMux I__4291 (
            .O(N__18564),
            .I(N__18505));
    SRMux I__4290 (
            .O(N__18563),
            .I(N__18502));
    SRMux I__4289 (
            .O(N__18562),
            .I(N__18499));
    LocalMux I__4288 (
            .O(N__18559),
            .I(N__18496));
    Span4Mux_v I__4287 (
            .O(N__18552),
            .I(N__18488));
    LocalMux I__4286 (
            .O(N__18549),
            .I(N__18488));
    LocalMux I__4285 (
            .O(N__18546),
            .I(N__18488));
    Span4Mux_v I__4284 (
            .O(N__18541),
            .I(N__18485));
    Span4Mux_s2_v I__4283 (
            .O(N__18538),
            .I(N__18478));
    LocalMux I__4282 (
            .O(N__18535),
            .I(N__18478));
    LocalMux I__4281 (
            .O(N__18532),
            .I(N__18478));
    Span4Mux_s2_v I__4280 (
            .O(N__18529),
            .I(N__18471));
    LocalMux I__4279 (
            .O(N__18526),
            .I(N__18471));
    LocalMux I__4278 (
            .O(N__18523),
            .I(N__18471));
    SRMux I__4277 (
            .O(N__18522),
            .I(N__18468));
    SRMux I__4276 (
            .O(N__18521),
            .I(N__18465));
    SRMux I__4275 (
            .O(N__18520),
            .I(N__18462));
    SRMux I__4274 (
            .O(N__18519),
            .I(N__18459));
    LocalMux I__4273 (
            .O(N__18516),
            .I(N__18456));
    SRMux I__4272 (
            .O(N__18515),
            .I(N__18453));
    SRMux I__4271 (
            .O(N__18514),
            .I(N__18450));
    Span12Mux_h I__4270 (
            .O(N__18511),
            .I(N__18447));
    Span4Mux_h I__4269 (
            .O(N__18508),
            .I(N__18444));
    Span12Mux_s9_h I__4268 (
            .O(N__18505),
            .I(N__18441));
    LocalMux I__4267 (
            .O(N__18502),
            .I(N__18438));
    LocalMux I__4266 (
            .O(N__18499),
            .I(N__18435));
    Span12Mux_s9_h I__4265 (
            .O(N__18496),
            .I(N__18432));
    SRMux I__4264 (
            .O(N__18495),
            .I(N__18429));
    Span4Mux_v I__4263 (
            .O(N__18488),
            .I(N__18426));
    Span4Mux_v I__4262 (
            .O(N__18485),
            .I(N__18415));
    Span4Mux_v I__4261 (
            .O(N__18478),
            .I(N__18415));
    Span4Mux_v I__4260 (
            .O(N__18471),
            .I(N__18415));
    LocalMux I__4259 (
            .O(N__18468),
            .I(N__18415));
    LocalMux I__4258 (
            .O(N__18465),
            .I(N__18415));
    LocalMux I__4257 (
            .O(N__18462),
            .I(N__18410));
    LocalMux I__4256 (
            .O(N__18459),
            .I(N__18410));
    Span4Mux_h I__4255 (
            .O(N__18456),
            .I(N__18403));
    LocalMux I__4254 (
            .O(N__18453),
            .I(N__18403));
    LocalMux I__4253 (
            .O(N__18450),
            .I(N__18403));
    Span12Mux_v I__4252 (
            .O(N__18447),
            .I(N__18400));
    Span4Mux_h I__4251 (
            .O(N__18444),
            .I(N__18397));
    Span12Mux_v I__4250 (
            .O(N__18441),
            .I(N__18392));
    Span12Mux_s9_h I__4249 (
            .O(N__18438),
            .I(N__18392));
    Span4Mux_h I__4248 (
            .O(N__18435),
            .I(N__18389));
    Span12Mux_v I__4247 (
            .O(N__18432),
            .I(N__18384));
    LocalMux I__4246 (
            .O(N__18429),
            .I(N__18384));
    Span4Mux_v I__4245 (
            .O(N__18426),
            .I(N__18375));
    Span4Mux_v I__4244 (
            .O(N__18415),
            .I(N__18375));
    Span4Mux_v I__4243 (
            .O(N__18410),
            .I(N__18375));
    Span4Mux_v I__4242 (
            .O(N__18403),
            .I(N__18375));
    Odrv12 I__4241 (
            .O(N__18400),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4240 (
            .O(N__18397),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4239 (
            .O(N__18392),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4238 (
            .O(N__18389),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4237 (
            .O(N__18384),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4236 (
            .O(N__18375),
            .I(CONSTANT_ONE_NET));
    InMux I__4235 (
            .O(N__18362),
            .I(N__18358));
    CascadeMux I__4234 (
            .O(N__18361),
            .I(N__18352));
    LocalMux I__4233 (
            .O(N__18358),
            .I(N__18349));
    InMux I__4232 (
            .O(N__18357),
            .I(N__18342));
    InMux I__4231 (
            .O(N__18356),
            .I(N__18339));
    InMux I__4230 (
            .O(N__18355),
            .I(N__18334));
    InMux I__4229 (
            .O(N__18352),
            .I(N__18334));
    Span12Mux_h I__4228 (
            .O(N__18349),
            .I(N__18331));
    CascadeMux I__4227 (
            .O(N__18348),
            .I(N__18328));
    InMux I__4226 (
            .O(N__18347),
            .I(N__18325));
    InMux I__4225 (
            .O(N__18346),
            .I(N__18320));
    InMux I__4224 (
            .O(N__18345),
            .I(N__18320));
    LocalMux I__4223 (
            .O(N__18342),
            .I(N__18315));
    LocalMux I__4222 (
            .O(N__18339),
            .I(N__18315));
    LocalMux I__4221 (
            .O(N__18334),
            .I(N__18312));
    Span12Mux_v I__4220 (
            .O(N__18331),
            .I(N__18307));
    InMux I__4219 (
            .O(N__18328),
            .I(N__18304));
    LocalMux I__4218 (
            .O(N__18325),
            .I(N__18301));
    LocalMux I__4217 (
            .O(N__18320),
            .I(N__18294));
    Span4Mux_h I__4216 (
            .O(N__18315),
            .I(N__18294));
    Span4Mux_v I__4215 (
            .O(N__18312),
            .I(N__18294));
    InMux I__4214 (
            .O(N__18311),
            .I(N__18289));
    InMux I__4213 (
            .O(N__18310),
            .I(N__18289));
    Odrv12 I__4212 (
            .O(N__18307),
            .I(\this_vga_signals.mult1_un61_sum_axbxc5 ));
    LocalMux I__4211 (
            .O(N__18304),
            .I(\this_vga_signals.mult1_un61_sum_axbxc5 ));
    Odrv4 I__4210 (
            .O(N__18301),
            .I(\this_vga_signals.mult1_un61_sum_axbxc5 ));
    Odrv4 I__4209 (
            .O(N__18294),
            .I(\this_vga_signals.mult1_un61_sum_axbxc5 ));
    LocalMux I__4208 (
            .O(N__18289),
            .I(\this_vga_signals.mult1_un61_sum_axbxc5 ));
    CascadeMux I__4207 (
            .O(N__18278),
            .I(N__18275));
    CascadeBuf I__4206 (
            .O(N__18275),
            .I(N__18272));
    CascadeMux I__4205 (
            .O(N__18272),
            .I(N__18269));
    CascadeBuf I__4204 (
            .O(N__18269),
            .I(N__18266));
    CascadeMux I__4203 (
            .O(N__18266),
            .I(N__18263));
    CascadeBuf I__4202 (
            .O(N__18263),
            .I(N__18260));
    CascadeMux I__4201 (
            .O(N__18260),
            .I(N__18257));
    CascadeBuf I__4200 (
            .O(N__18257),
            .I(N__18254));
    CascadeMux I__4199 (
            .O(N__18254),
            .I(N__18251));
    CascadeBuf I__4198 (
            .O(N__18251),
            .I(N__18248));
    CascadeMux I__4197 (
            .O(N__18248),
            .I(N__18245));
    CascadeBuf I__4196 (
            .O(N__18245),
            .I(N__18242));
    CascadeMux I__4195 (
            .O(N__18242),
            .I(N__18239));
    CascadeBuf I__4194 (
            .O(N__18239),
            .I(N__18236));
    CascadeMux I__4193 (
            .O(N__18236),
            .I(N__18233));
    CascadeBuf I__4192 (
            .O(N__18233),
            .I(N__18230));
    CascadeMux I__4191 (
            .O(N__18230),
            .I(N__18227));
    CascadeBuf I__4190 (
            .O(N__18227),
            .I(N__18224));
    CascadeMux I__4189 (
            .O(N__18224),
            .I(N__18221));
    CascadeBuf I__4188 (
            .O(N__18221),
            .I(N__18218));
    CascadeMux I__4187 (
            .O(N__18218),
            .I(N__18215));
    CascadeBuf I__4186 (
            .O(N__18215),
            .I(N__18212));
    CascadeMux I__4185 (
            .O(N__18212),
            .I(N__18209));
    CascadeBuf I__4184 (
            .O(N__18209),
            .I(N__18206));
    CascadeMux I__4183 (
            .O(N__18206),
            .I(N__18203));
    CascadeBuf I__4182 (
            .O(N__18203),
            .I(N__18200));
    CascadeMux I__4181 (
            .O(N__18200),
            .I(N__18197));
    CascadeBuf I__4180 (
            .O(N__18197),
            .I(N__18194));
    CascadeMux I__4179 (
            .O(N__18194),
            .I(N__18191));
    CascadeBuf I__4178 (
            .O(N__18191),
            .I(N__18188));
    CascadeMux I__4177 (
            .O(N__18188),
            .I(N__18185));
    InMux I__4176 (
            .O(N__18185),
            .I(N__18182));
    LocalMux I__4175 (
            .O(N__18182),
            .I(N__18179));
    Odrv4 I__4174 (
            .O(N__18179),
            .I(M_this_vga_signals_address_5));
    InMux I__4173 (
            .O(N__18176),
            .I(N__18173));
    LocalMux I__4172 (
            .O(N__18173),
            .I(N__18170));
    Span4Mux_v I__4171 (
            .O(N__18170),
            .I(N__18167));
    Odrv4 I__4170 (
            .O(N__18167),
            .I(\this_vram.mem_out_bus1_2 ));
    InMux I__4169 (
            .O(N__18164),
            .I(N__18161));
    LocalMux I__4168 (
            .O(N__18161),
            .I(N__18158));
    Span4Mux_v I__4167 (
            .O(N__18158),
            .I(N__18155));
    Span4Mux_v I__4166 (
            .O(N__18155),
            .I(N__18152));
    Odrv4 I__4165 (
            .O(N__18152),
            .I(\this_vram.mem_out_bus5_2 ));
    InMux I__4164 (
            .O(N__18149),
            .I(N__18146));
    LocalMux I__4163 (
            .O(N__18146),
            .I(N__18143));
    Span4Mux_v I__4162 (
            .O(N__18143),
            .I(N__18140));
    Span4Mux_v I__4161 (
            .O(N__18140),
            .I(N__18137));
    Odrv4 I__4160 (
            .O(N__18137),
            .I(\this_vram.mem_out_bus1_1 ));
    InMux I__4159 (
            .O(N__18134),
            .I(N__18131));
    LocalMux I__4158 (
            .O(N__18131),
            .I(N__18128));
    Sp12to4 I__4157 (
            .O(N__18128),
            .I(N__18125));
    Odrv12 I__4156 (
            .O(N__18125),
            .I(\this_vram.mem_out_bus5_1 ));
    InMux I__4155 (
            .O(N__18122),
            .I(N__18119));
    LocalMux I__4154 (
            .O(N__18119),
            .I(N__18116));
    Span4Mux_v I__4153 (
            .O(N__18116),
            .I(N__18113));
    Odrv4 I__4152 (
            .O(N__18113),
            .I(\this_vram.mem_mem_1_0_RNISSK11Z0Z_0 ));
    InMux I__4151 (
            .O(N__18110),
            .I(N__18107));
    LocalMux I__4150 (
            .O(N__18107),
            .I(N__18104));
    Span4Mux_v I__4149 (
            .O(N__18104),
            .I(N__18101));
    Span4Mux_v I__4148 (
            .O(N__18101),
            .I(N__18098));
    Odrv4 I__4147 (
            .O(N__18098),
            .I(\this_vram.mem_out_bus6_0 ));
    InMux I__4146 (
            .O(N__18095),
            .I(N__18092));
    LocalMux I__4145 (
            .O(N__18092),
            .I(N__18089));
    Span4Mux_v I__4144 (
            .O(N__18089),
            .I(N__18086));
    Odrv4 I__4143 (
            .O(N__18086),
            .I(\this_vram.mem_out_bus2_0 ));
    CascadeMux I__4142 (
            .O(N__18083),
            .I(\this_vram.mem_mem_2_0_RNIU0NZ0Z11_cascade_ ));
    InMux I__4141 (
            .O(N__18080),
            .I(N__18076));
    InMux I__4140 (
            .O(N__18079),
            .I(N__18073));
    LocalMux I__4139 (
            .O(N__18076),
            .I(N__18068));
    LocalMux I__4138 (
            .O(N__18073),
            .I(N__18068));
    Span4Mux_v I__4137 (
            .O(N__18068),
            .I(N__18065));
    Span4Mux_h I__4136 (
            .O(N__18065),
            .I(N__18062));
    Odrv4 I__4135 (
            .O(N__18062),
            .I(\this_vram.mem_N_112 ));
    InMux I__4134 (
            .O(N__18059),
            .I(N__18056));
    LocalMux I__4133 (
            .O(N__18056),
            .I(N__18053));
    Odrv4 I__4132 (
            .O(N__18053),
            .I(\this_vram.mem_out_bus4_0 ));
    InMux I__4131 (
            .O(N__18050),
            .I(N__18047));
    LocalMux I__4130 (
            .O(N__18047),
            .I(N__18044));
    Sp12to4 I__4129 (
            .O(N__18044),
            .I(N__18041));
    Span12Mux_v I__4128 (
            .O(N__18041),
            .I(N__18038));
    Odrv12 I__4127 (
            .O(N__18038),
            .I(\this_vram.mem_out_bus0_0 ));
    InMux I__4126 (
            .O(N__18035),
            .I(N__18032));
    LocalMux I__4125 (
            .O(N__18032),
            .I(\this_vram.mem_mem_0_0_RNIQOIZ0Z11 ));
    InMux I__4124 (
            .O(N__18029),
            .I(N__18026));
    LocalMux I__4123 (
            .O(N__18026),
            .I(\this_vram.mem_out_bus3_2 ));
    InMux I__4122 (
            .O(N__18023),
            .I(N__18020));
    LocalMux I__4121 (
            .O(N__18020),
            .I(N__18017));
    Sp12to4 I__4120 (
            .O(N__18017),
            .I(N__18014));
    Span12Mux_v I__4119 (
            .O(N__18014),
            .I(N__18011));
    Odrv12 I__4118 (
            .O(N__18011),
            .I(\this_vram.mem_out_bus7_2 ));
    InMux I__4117 (
            .O(N__18008),
            .I(N__18005));
    LocalMux I__4116 (
            .O(N__18005),
            .I(N__18002));
    Span4Mux_h I__4115 (
            .O(N__18002),
            .I(N__17999));
    Sp12to4 I__4114 (
            .O(N__17999),
            .I(N__17996));
    Odrv12 I__4113 (
            .O(N__17996),
            .I(\this_vram.mem_out_bus6_1 ));
    InMux I__4112 (
            .O(N__17993),
            .I(N__17990));
    LocalMux I__4111 (
            .O(N__17990),
            .I(N__17987));
    Odrv4 I__4110 (
            .O(N__17987),
            .I(\this_vram.mem_mem_2_0_RNIU0N11Z0Z_0 ));
    CEMux I__4109 (
            .O(N__17984),
            .I(N__17981));
    LocalMux I__4108 (
            .O(N__17981),
            .I(N__17977));
    CEMux I__4107 (
            .O(N__17980),
            .I(N__17974));
    Span4Mux_h I__4106 (
            .O(N__17977),
            .I(N__17971));
    LocalMux I__4105 (
            .O(N__17974),
            .I(N__17968));
    Sp12to4 I__4104 (
            .O(N__17971),
            .I(N__17965));
    Span4Mux_h I__4103 (
            .O(N__17968),
            .I(N__17962));
    Span12Mux_v I__4102 (
            .O(N__17965),
            .I(N__17959));
    Sp12to4 I__4101 (
            .O(N__17962),
            .I(N__17956));
    Odrv12 I__4100 (
            .O(N__17959),
            .I(\this_vram.mem_WE_14 ));
    Odrv12 I__4099 (
            .O(N__17956),
            .I(\this_vram.mem_WE_14 ));
    CEMux I__4098 (
            .O(N__17951),
            .I(N__17948));
    LocalMux I__4097 (
            .O(N__17948),
            .I(N__17944));
    CEMux I__4096 (
            .O(N__17947),
            .I(N__17941));
    Span4Mux_v I__4095 (
            .O(N__17944),
            .I(N__17938));
    LocalMux I__4094 (
            .O(N__17941),
            .I(N__17935));
    Span4Mux_v I__4093 (
            .O(N__17938),
            .I(N__17932));
    Span4Mux_h I__4092 (
            .O(N__17935),
            .I(N__17929));
    Odrv4 I__4091 (
            .O(N__17932),
            .I(\this_vram.mem_WE_10 ));
    Odrv4 I__4090 (
            .O(N__17929),
            .I(\this_vram.mem_WE_10 ));
    InMux I__4089 (
            .O(N__17924),
            .I(N__17921));
    LocalMux I__4088 (
            .O(N__17921),
            .I(M_this_vram_read_data_3));
    InMux I__4087 (
            .O(N__17918),
            .I(N__17915));
    LocalMux I__4086 (
            .O(N__17915),
            .I(N__17912));
    Odrv4 I__4085 (
            .O(N__17912),
            .I(\this_vram.mem_out_bus4_1 ));
    InMux I__4084 (
            .O(N__17909),
            .I(N__17906));
    LocalMux I__4083 (
            .O(N__17906),
            .I(N__17903));
    Span12Mux_h I__4082 (
            .O(N__17903),
            .I(N__17900));
    Span12Mux_v I__4081 (
            .O(N__17900),
            .I(N__17897));
    Odrv12 I__4080 (
            .O(N__17897),
            .I(\this_vram.mem_out_bus0_1 ));
    InMux I__4079 (
            .O(N__17894),
            .I(N__17891));
    LocalMux I__4078 (
            .O(N__17891),
            .I(\this_vram.mem_mem_0_0_RNIQOI11Z0Z_0 ));
    InMux I__4077 (
            .O(N__17888),
            .I(N__17885));
    LocalMux I__4076 (
            .O(N__17885),
            .I(N__17882));
    Span4Mux_h I__4075 (
            .O(N__17882),
            .I(N__17879));
    Sp12to4 I__4074 (
            .O(N__17879),
            .I(N__17876));
    Span12Mux_v I__4073 (
            .O(N__17876),
            .I(N__17873));
    Odrv12 I__4072 (
            .O(N__17873),
            .I(\this_vram.mem_out_bus7_3 ));
    InMux I__4071 (
            .O(N__17870),
            .I(N__17867));
    LocalMux I__4070 (
            .O(N__17867),
            .I(N__17864));
    Span4Mux_v I__4069 (
            .O(N__17864),
            .I(N__17861));
    Odrv4 I__4068 (
            .O(N__17861),
            .I(\this_vram.mem_out_bus3_3 ));
    CascadeMux I__4067 (
            .O(N__17858),
            .I(\this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_ ));
    InMux I__4066 (
            .O(N__17855),
            .I(N__17852));
    LocalMux I__4065 (
            .O(N__17852),
            .I(\this_vram.mem_N_102 ));
    InMux I__4064 (
            .O(N__17849),
            .I(N__17845));
    InMux I__4063 (
            .O(N__17848),
            .I(N__17842));
    LocalMux I__4062 (
            .O(N__17845),
            .I(N__17838));
    LocalMux I__4061 (
            .O(N__17842),
            .I(N__17834));
    InMux I__4060 (
            .O(N__17841),
            .I(N__17831));
    Span4Mux_h I__4059 (
            .O(N__17838),
            .I(N__17827));
    InMux I__4058 (
            .O(N__17837),
            .I(N__17824));
    Span4Mux_h I__4057 (
            .O(N__17834),
            .I(N__17819));
    LocalMux I__4056 (
            .O(N__17831),
            .I(N__17819));
    InMux I__4055 (
            .O(N__17830),
            .I(N__17816));
    Span4Mux_h I__4054 (
            .O(N__17827),
            .I(N__17811));
    LocalMux I__4053 (
            .O(N__17824),
            .I(N__17811));
    Span4Mux_h I__4052 (
            .O(N__17819),
            .I(N__17806));
    LocalMux I__4051 (
            .O(N__17816),
            .I(N__17806));
    Span4Mux_h I__4050 (
            .O(N__17811),
            .I(N__17803));
    Span4Mux_h I__4049 (
            .O(N__17806),
            .I(N__17800));
    Span4Mux_h I__4048 (
            .O(N__17803),
            .I(N__17795));
    Span4Mux_v I__4047 (
            .O(N__17800),
            .I(N__17792));
    InMux I__4046 (
            .O(N__17799),
            .I(N__17789));
    InMux I__4045 (
            .O(N__17798),
            .I(N__17786));
    Odrv4 I__4044 (
            .O(N__17795),
            .I(\this_vram.mem_radregZ0Z_11 ));
    Odrv4 I__4043 (
            .O(N__17792),
            .I(\this_vram.mem_radregZ0Z_11 ));
    LocalMux I__4042 (
            .O(N__17789),
            .I(\this_vram.mem_radregZ0Z_11 ));
    LocalMux I__4041 (
            .O(N__17786),
            .I(\this_vram.mem_radregZ0Z_11 ));
    InMux I__4040 (
            .O(N__17777),
            .I(N__17774));
    LocalMux I__4039 (
            .O(N__17774),
            .I(M_this_vram_read_data_2));
    CEMux I__4038 (
            .O(N__17771),
            .I(N__17768));
    LocalMux I__4037 (
            .O(N__17768),
            .I(N__17764));
    CEMux I__4036 (
            .O(N__17767),
            .I(N__17761));
    Span4Mux_v I__4035 (
            .O(N__17764),
            .I(N__17756));
    LocalMux I__4034 (
            .O(N__17761),
            .I(N__17756));
    Span4Mux_v I__4033 (
            .O(N__17756),
            .I(N__17753));
    Span4Mux_v I__4032 (
            .O(N__17753),
            .I(N__17750));
    Span4Mux_v I__4031 (
            .O(N__17750),
            .I(N__17747));
    Odrv4 I__4030 (
            .O(N__17747),
            .I(\this_vram.mem_WE_12 ));
    InMux I__4029 (
            .O(N__17744),
            .I(N__17741));
    LocalMux I__4028 (
            .O(N__17741),
            .I(N__17734));
    InMux I__4027 (
            .O(N__17740),
            .I(N__17731));
    IoInMux I__4026 (
            .O(N__17739),
            .I(N__17728));
    InMux I__4025 (
            .O(N__17738),
            .I(N__17724));
    CascadeMux I__4024 (
            .O(N__17737),
            .I(N__17721));
    Span4Mux_h I__4023 (
            .O(N__17734),
            .I(N__17716));
    LocalMux I__4022 (
            .O(N__17731),
            .I(N__17716));
    LocalMux I__4021 (
            .O(N__17728),
            .I(N__17713));
    CascadeMux I__4020 (
            .O(N__17727),
            .I(N__17706));
    LocalMux I__4019 (
            .O(N__17724),
            .I(N__17703));
    InMux I__4018 (
            .O(N__17721),
            .I(N__17700));
    Sp12to4 I__4017 (
            .O(N__17716),
            .I(N__17697));
    Span4Mux_s2_v I__4016 (
            .O(N__17713),
            .I(N__17694));
    CascadeMux I__4015 (
            .O(N__17712),
            .I(N__17691));
    CascadeMux I__4014 (
            .O(N__17711),
            .I(N__17688));
    InMux I__4013 (
            .O(N__17710),
            .I(N__17682));
    InMux I__4012 (
            .O(N__17709),
            .I(N__17679));
    InMux I__4011 (
            .O(N__17706),
            .I(N__17676));
    Span4Mux_v I__4010 (
            .O(N__17703),
            .I(N__17673));
    LocalMux I__4009 (
            .O(N__17700),
            .I(N__17670));
    Span12Mux_v I__4008 (
            .O(N__17697),
            .I(N__17665));
    Sp12to4 I__4007 (
            .O(N__17694),
            .I(N__17665));
    InMux I__4006 (
            .O(N__17691),
            .I(N__17658));
    InMux I__4005 (
            .O(N__17688),
            .I(N__17658));
    InMux I__4004 (
            .O(N__17687),
            .I(N__17658));
    InMux I__4003 (
            .O(N__17686),
            .I(N__17653));
    InMux I__4002 (
            .O(N__17685),
            .I(N__17653));
    LocalMux I__4001 (
            .O(N__17682),
            .I(N__17646));
    LocalMux I__4000 (
            .O(N__17679),
            .I(N__17646));
    LocalMux I__3999 (
            .O(N__17676),
            .I(N__17646));
    Span4Mux_h I__3998 (
            .O(N__17673),
            .I(N__17641));
    Span4Mux_v I__3997 (
            .O(N__17670),
            .I(N__17641));
    Span12Mux_h I__3996 (
            .O(N__17665),
            .I(N__17638));
    LocalMux I__3995 (
            .O(N__17658),
            .I(M_this_reset_cond_out_0));
    LocalMux I__3994 (
            .O(N__17653),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__3993 (
            .O(N__17646),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__3992 (
            .O(N__17641),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__3991 (
            .O(N__17638),
            .I(M_this_reset_cond_out_0));
    CascadeMux I__3990 (
            .O(N__17627),
            .I(N__17620));
    CascadeMux I__3989 (
            .O(N__17626),
            .I(N__17616));
    InMux I__3988 (
            .O(N__17625),
            .I(N__17609));
    InMux I__3987 (
            .O(N__17624),
            .I(N__17599));
    InMux I__3986 (
            .O(N__17623),
            .I(N__17599));
    InMux I__3985 (
            .O(N__17620),
            .I(N__17592));
    InMux I__3984 (
            .O(N__17619),
            .I(N__17592));
    InMux I__3983 (
            .O(N__17616),
            .I(N__17592));
    InMux I__3982 (
            .O(N__17615),
            .I(N__17589));
    InMux I__3981 (
            .O(N__17614),
            .I(N__17584));
    InMux I__3980 (
            .O(N__17613),
            .I(N__17584));
    InMux I__3979 (
            .O(N__17612),
            .I(N__17581));
    LocalMux I__3978 (
            .O(N__17609),
            .I(N__17578));
    InMux I__3977 (
            .O(N__17608),
            .I(N__17575));
    InMux I__3976 (
            .O(N__17607),
            .I(N__17570));
    InMux I__3975 (
            .O(N__17606),
            .I(N__17570));
    InMux I__3974 (
            .O(N__17605),
            .I(N__17562));
    InMux I__3973 (
            .O(N__17604),
            .I(N__17562));
    LocalMux I__3972 (
            .O(N__17599),
            .I(N__17557));
    LocalMux I__3971 (
            .O(N__17592),
            .I(N__17557));
    LocalMux I__3970 (
            .O(N__17589),
            .I(N__17546));
    LocalMux I__3969 (
            .O(N__17584),
            .I(N__17546));
    LocalMux I__3968 (
            .O(N__17581),
            .I(N__17546));
    Span4Mux_v I__3967 (
            .O(N__17578),
            .I(N__17546));
    LocalMux I__3966 (
            .O(N__17575),
            .I(N__17546));
    LocalMux I__3965 (
            .O(N__17570),
            .I(N__17543));
    InMux I__3964 (
            .O(N__17569),
            .I(N__17540));
    InMux I__3963 (
            .O(N__17568),
            .I(N__17537));
    InMux I__3962 (
            .O(N__17567),
            .I(N__17534));
    LocalMux I__3961 (
            .O(N__17562),
            .I(N__17531));
    Span4Mux_v I__3960 (
            .O(N__17557),
            .I(N__17528));
    Span4Mux_h I__3959 (
            .O(N__17546),
            .I(N__17525));
    Span4Mux_v I__3958 (
            .O(N__17543),
            .I(N__17520));
    LocalMux I__3957 (
            .O(N__17540),
            .I(N__17520));
    LocalMux I__3956 (
            .O(N__17537),
            .I(M_this_start_data_delay_out_0));
    LocalMux I__3955 (
            .O(N__17534),
            .I(M_this_start_data_delay_out_0));
    Odrv12 I__3954 (
            .O(N__17531),
            .I(M_this_start_data_delay_out_0));
    Odrv4 I__3953 (
            .O(N__17528),
            .I(M_this_start_data_delay_out_0));
    Odrv4 I__3952 (
            .O(N__17525),
            .I(M_this_start_data_delay_out_0));
    Odrv4 I__3951 (
            .O(N__17520),
            .I(M_this_start_data_delay_out_0));
    CascadeMux I__3950 (
            .O(N__17507),
            .I(M_state_q_ns_1_0__i12_mux_cascade_));
    CascadeMux I__3949 (
            .O(N__17504),
            .I(N__17496));
    InMux I__3948 (
            .O(N__17503),
            .I(N__17493));
    InMux I__3947 (
            .O(N__17502),
            .I(N__17490));
    CascadeMux I__3946 (
            .O(N__17501),
            .I(N__17487));
    InMux I__3945 (
            .O(N__17500),
            .I(N__17472));
    InMux I__3944 (
            .O(N__17499),
            .I(N__17472));
    InMux I__3943 (
            .O(N__17496),
            .I(N__17469));
    LocalMux I__3942 (
            .O(N__17493),
            .I(N__17464));
    LocalMux I__3941 (
            .O(N__17490),
            .I(N__17464));
    InMux I__3940 (
            .O(N__17487),
            .I(N__17457));
    InMux I__3939 (
            .O(N__17486),
            .I(N__17457));
    InMux I__3938 (
            .O(N__17485),
            .I(N__17457));
    InMux I__3937 (
            .O(N__17484),
            .I(N__17454));
    InMux I__3936 (
            .O(N__17483),
            .I(N__17446));
    InMux I__3935 (
            .O(N__17482),
            .I(N__17446));
    InMux I__3934 (
            .O(N__17481),
            .I(N__17443));
    InMux I__3933 (
            .O(N__17480),
            .I(N__17434));
    InMux I__3932 (
            .O(N__17479),
            .I(N__17434));
    InMux I__3931 (
            .O(N__17478),
            .I(N__17434));
    InMux I__3930 (
            .O(N__17477),
            .I(N__17434));
    LocalMux I__3929 (
            .O(N__17472),
            .I(N__17431));
    LocalMux I__3928 (
            .O(N__17469),
            .I(N__17426));
    Span4Mux_h I__3927 (
            .O(N__17464),
            .I(N__17426));
    LocalMux I__3926 (
            .O(N__17457),
            .I(N__17421));
    LocalMux I__3925 (
            .O(N__17454),
            .I(N__17421));
    InMux I__3924 (
            .O(N__17453),
            .I(N__17418));
    InMux I__3923 (
            .O(N__17452),
            .I(N__17415));
    InMux I__3922 (
            .O(N__17451),
            .I(N__17412));
    LocalMux I__3921 (
            .O(N__17446),
            .I(N__17407));
    LocalMux I__3920 (
            .O(N__17443),
            .I(N__17407));
    LocalMux I__3919 (
            .O(N__17434),
            .I(N__17404));
    Span4Mux_h I__3918 (
            .O(N__17431),
            .I(N__17401));
    Span4Mux_v I__3917 (
            .O(N__17426),
            .I(N__17396));
    Span4Mux_h I__3916 (
            .O(N__17421),
            .I(N__17396));
    LocalMux I__3915 (
            .O(N__17418),
            .I(N__17393));
    LocalMux I__3914 (
            .O(N__17415),
            .I(M_state_qZ0Z_1));
    LocalMux I__3913 (
            .O(N__17412),
            .I(M_state_qZ0Z_1));
    Odrv4 I__3912 (
            .O(N__17407),
            .I(M_state_qZ0Z_1));
    Odrv4 I__3911 (
            .O(N__17404),
            .I(M_state_qZ0Z_1));
    Odrv4 I__3910 (
            .O(N__17401),
            .I(M_state_qZ0Z_1));
    Odrv4 I__3909 (
            .O(N__17396),
            .I(M_state_qZ0Z_1));
    Odrv12 I__3908 (
            .O(N__17393),
            .I(M_state_qZ0Z_1));
    ClkMux I__3907 (
            .O(N__17378),
            .I(N__17147));
    ClkMux I__3906 (
            .O(N__17377),
            .I(N__17147));
    ClkMux I__3905 (
            .O(N__17376),
            .I(N__17147));
    ClkMux I__3904 (
            .O(N__17375),
            .I(N__17147));
    ClkMux I__3903 (
            .O(N__17374),
            .I(N__17147));
    ClkMux I__3902 (
            .O(N__17373),
            .I(N__17147));
    ClkMux I__3901 (
            .O(N__17372),
            .I(N__17147));
    ClkMux I__3900 (
            .O(N__17371),
            .I(N__17147));
    ClkMux I__3899 (
            .O(N__17370),
            .I(N__17147));
    ClkMux I__3898 (
            .O(N__17369),
            .I(N__17147));
    ClkMux I__3897 (
            .O(N__17368),
            .I(N__17147));
    ClkMux I__3896 (
            .O(N__17367),
            .I(N__17147));
    ClkMux I__3895 (
            .O(N__17366),
            .I(N__17147));
    ClkMux I__3894 (
            .O(N__17365),
            .I(N__17147));
    ClkMux I__3893 (
            .O(N__17364),
            .I(N__17147));
    ClkMux I__3892 (
            .O(N__17363),
            .I(N__17147));
    ClkMux I__3891 (
            .O(N__17362),
            .I(N__17147));
    ClkMux I__3890 (
            .O(N__17361),
            .I(N__17147));
    ClkMux I__3889 (
            .O(N__17360),
            .I(N__17147));
    ClkMux I__3888 (
            .O(N__17359),
            .I(N__17147));
    ClkMux I__3887 (
            .O(N__17358),
            .I(N__17147));
    ClkMux I__3886 (
            .O(N__17357),
            .I(N__17147));
    ClkMux I__3885 (
            .O(N__17356),
            .I(N__17147));
    ClkMux I__3884 (
            .O(N__17355),
            .I(N__17147));
    ClkMux I__3883 (
            .O(N__17354),
            .I(N__17147));
    ClkMux I__3882 (
            .O(N__17353),
            .I(N__17147));
    ClkMux I__3881 (
            .O(N__17352),
            .I(N__17147));
    ClkMux I__3880 (
            .O(N__17351),
            .I(N__17147));
    ClkMux I__3879 (
            .O(N__17350),
            .I(N__17147));
    ClkMux I__3878 (
            .O(N__17349),
            .I(N__17147));
    ClkMux I__3877 (
            .O(N__17348),
            .I(N__17147));
    ClkMux I__3876 (
            .O(N__17347),
            .I(N__17147));
    ClkMux I__3875 (
            .O(N__17346),
            .I(N__17147));
    ClkMux I__3874 (
            .O(N__17345),
            .I(N__17147));
    ClkMux I__3873 (
            .O(N__17344),
            .I(N__17147));
    ClkMux I__3872 (
            .O(N__17343),
            .I(N__17147));
    ClkMux I__3871 (
            .O(N__17342),
            .I(N__17147));
    ClkMux I__3870 (
            .O(N__17341),
            .I(N__17147));
    ClkMux I__3869 (
            .O(N__17340),
            .I(N__17147));
    ClkMux I__3868 (
            .O(N__17339),
            .I(N__17147));
    ClkMux I__3867 (
            .O(N__17338),
            .I(N__17147));
    ClkMux I__3866 (
            .O(N__17337),
            .I(N__17147));
    ClkMux I__3865 (
            .O(N__17336),
            .I(N__17147));
    ClkMux I__3864 (
            .O(N__17335),
            .I(N__17147));
    ClkMux I__3863 (
            .O(N__17334),
            .I(N__17147));
    ClkMux I__3862 (
            .O(N__17333),
            .I(N__17147));
    ClkMux I__3861 (
            .O(N__17332),
            .I(N__17147));
    ClkMux I__3860 (
            .O(N__17331),
            .I(N__17147));
    ClkMux I__3859 (
            .O(N__17330),
            .I(N__17147));
    ClkMux I__3858 (
            .O(N__17329),
            .I(N__17147));
    ClkMux I__3857 (
            .O(N__17328),
            .I(N__17147));
    ClkMux I__3856 (
            .O(N__17327),
            .I(N__17147));
    ClkMux I__3855 (
            .O(N__17326),
            .I(N__17147));
    ClkMux I__3854 (
            .O(N__17325),
            .I(N__17147));
    ClkMux I__3853 (
            .O(N__17324),
            .I(N__17147));
    ClkMux I__3852 (
            .O(N__17323),
            .I(N__17147));
    ClkMux I__3851 (
            .O(N__17322),
            .I(N__17147));
    ClkMux I__3850 (
            .O(N__17321),
            .I(N__17147));
    ClkMux I__3849 (
            .O(N__17320),
            .I(N__17147));
    ClkMux I__3848 (
            .O(N__17319),
            .I(N__17147));
    ClkMux I__3847 (
            .O(N__17318),
            .I(N__17147));
    ClkMux I__3846 (
            .O(N__17317),
            .I(N__17147));
    ClkMux I__3845 (
            .O(N__17316),
            .I(N__17147));
    ClkMux I__3844 (
            .O(N__17315),
            .I(N__17147));
    ClkMux I__3843 (
            .O(N__17314),
            .I(N__17147));
    ClkMux I__3842 (
            .O(N__17313),
            .I(N__17147));
    ClkMux I__3841 (
            .O(N__17312),
            .I(N__17147));
    ClkMux I__3840 (
            .O(N__17311),
            .I(N__17147));
    ClkMux I__3839 (
            .O(N__17310),
            .I(N__17147));
    ClkMux I__3838 (
            .O(N__17309),
            .I(N__17147));
    ClkMux I__3837 (
            .O(N__17308),
            .I(N__17147));
    ClkMux I__3836 (
            .O(N__17307),
            .I(N__17147));
    ClkMux I__3835 (
            .O(N__17306),
            .I(N__17147));
    ClkMux I__3834 (
            .O(N__17305),
            .I(N__17147));
    ClkMux I__3833 (
            .O(N__17304),
            .I(N__17147));
    ClkMux I__3832 (
            .O(N__17303),
            .I(N__17147));
    ClkMux I__3831 (
            .O(N__17302),
            .I(N__17147));
    GlobalMux I__3830 (
            .O(N__17147),
            .I(N__17144));
    gio2CtrlBuf I__3829 (
            .O(N__17144),
            .I(clk_c_g));
    CascadeMux I__3828 (
            .O(N__17141),
            .I(N__17137));
    InMux I__3827 (
            .O(N__17140),
            .I(N__17131));
    InMux I__3826 (
            .O(N__17137),
            .I(N__17131));
    InMux I__3825 (
            .O(N__17136),
            .I(N__17128));
    LocalMux I__3824 (
            .O(N__17131),
            .I(N__17125));
    LocalMux I__3823 (
            .O(N__17128),
            .I(N__17122));
    Span12Mux_h I__3822 (
            .O(N__17125),
            .I(N__17119));
    Span12Mux_h I__3821 (
            .O(N__17122),
            .I(N__17116));
    Odrv12 I__3820 (
            .O(N__17119),
            .I(port_data_c_0));
    Odrv12 I__3819 (
            .O(N__17116),
            .I(port_data_c_0));
    InMux I__3818 (
            .O(N__17111),
            .I(N__17108));
    LocalMux I__3817 (
            .O(N__17108),
            .I(N__17104));
    InMux I__3816 (
            .O(N__17107),
            .I(N__17101));
    Span4Mux_s2_v I__3815 (
            .O(N__17104),
            .I(N__17095));
    LocalMux I__3814 (
            .O(N__17101),
            .I(N__17095));
    InMux I__3813 (
            .O(N__17100),
            .I(N__17092));
    Span4Mux_v I__3812 (
            .O(N__17095),
            .I(N__17086));
    LocalMux I__3811 (
            .O(N__17092),
            .I(N__17086));
    InMux I__3810 (
            .O(N__17091),
            .I(N__17083));
    Span4Mux_v I__3809 (
            .O(N__17086),
            .I(N__17077));
    LocalMux I__3808 (
            .O(N__17083),
            .I(N__17077));
    InMux I__3807 (
            .O(N__17082),
            .I(N__17074));
    Span4Mux_v I__3806 (
            .O(N__17077),
            .I(N__17067));
    LocalMux I__3805 (
            .O(N__17074),
            .I(N__17067));
    InMux I__3804 (
            .O(N__17073),
            .I(N__17064));
    InMux I__3803 (
            .O(N__17072),
            .I(N__17060));
    Span4Mux_v I__3802 (
            .O(N__17067),
            .I(N__17055));
    LocalMux I__3801 (
            .O(N__17064),
            .I(N__17055));
    InMux I__3800 (
            .O(N__17063),
            .I(N__17052));
    LocalMux I__3799 (
            .O(N__17060),
            .I(N__17049));
    Span4Mux_v I__3798 (
            .O(N__17055),
            .I(N__17044));
    LocalMux I__3797 (
            .O(N__17052),
            .I(N__17044));
    Span4Mux_v I__3796 (
            .O(N__17049),
            .I(N__17039));
    Span4Mux_v I__3795 (
            .O(N__17044),
            .I(N__17039));
    Odrv4 I__3794 (
            .O(N__17039),
            .I(M_this_vram_write_data_0));
    CEMux I__3793 (
            .O(N__17036),
            .I(N__17033));
    LocalMux I__3792 (
            .O(N__17033),
            .I(N__17029));
    CEMux I__3791 (
            .O(N__17032),
            .I(N__17026));
    Span4Mux_v I__3790 (
            .O(N__17029),
            .I(N__17023));
    LocalMux I__3789 (
            .O(N__17026),
            .I(N__17020));
    Odrv4 I__3788 (
            .O(N__17023),
            .I(\this_vram.mem_WE_8 ));
    Odrv12 I__3787 (
            .O(N__17020),
            .I(\this_vram.mem_WE_8 ));
    InMux I__3786 (
            .O(N__17015),
            .I(N__17012));
    LocalMux I__3785 (
            .O(N__17012),
            .I(N__17008));
    InMux I__3784 (
            .O(N__17011),
            .I(N__17005));
    Span4Mux_v I__3783 (
            .O(N__17008),
            .I(N__17000));
    LocalMux I__3782 (
            .O(N__17005),
            .I(N__17000));
    Sp12to4 I__3781 (
            .O(N__17000),
            .I(N__16996));
    InMux I__3780 (
            .O(N__16999),
            .I(N__16993));
    Span12Mux_v I__3779 (
            .O(N__16996),
            .I(N__16988));
    LocalMux I__3778 (
            .O(N__16993),
            .I(N__16988));
    Odrv12 I__3777 (
            .O(N__16988),
            .I(\this_vram.mem_N_91 ));
    InMux I__3776 (
            .O(N__16985),
            .I(N__16981));
    InMux I__3775 (
            .O(N__16984),
            .I(N__16978));
    LocalMux I__3774 (
            .O(N__16981),
            .I(N__16972));
    LocalMux I__3773 (
            .O(N__16978),
            .I(N__16972));
    InMux I__3772 (
            .O(N__16977),
            .I(N__16969));
    Span4Mux_v I__3771 (
            .O(N__16972),
            .I(N__16966));
    LocalMux I__3770 (
            .O(N__16969),
            .I(N__16963));
    Span4Mux_h I__3769 (
            .O(N__16966),
            .I(N__16958));
    Span4Mux_v I__3768 (
            .O(N__16963),
            .I(N__16958));
    Span4Mux_h I__3767 (
            .O(N__16958),
            .I(N__16955));
    Odrv4 I__3766 (
            .O(N__16955),
            .I(\this_vram.mem_N_88 ));
    InMux I__3765 (
            .O(N__16952),
            .I(N__16948));
    CascadeMux I__3764 (
            .O(N__16951),
            .I(N__16945));
    LocalMux I__3763 (
            .O(N__16948),
            .I(N__16942));
    InMux I__3762 (
            .O(N__16945),
            .I(N__16939));
    Span4Mux_h I__3761 (
            .O(N__16942),
            .I(N__16936));
    LocalMux I__3760 (
            .O(N__16939),
            .I(N__16933));
    Span4Mux_h I__3759 (
            .O(N__16936),
            .I(N__16930));
    Span4Mux_h I__3758 (
            .O(N__16933),
            .I(N__16927));
    Odrv4 I__3757 (
            .O(N__16930),
            .I(N_16_0));
    Odrv4 I__3756 (
            .O(N__16927),
            .I(N_16_0));
    InMux I__3755 (
            .O(N__16922),
            .I(N__16919));
    LocalMux I__3754 (
            .O(N__16919),
            .I(N__16916));
    Span12Mux_s9_v I__3753 (
            .O(N__16916),
            .I(N__16913));
    Odrv12 I__3752 (
            .O(N__16913),
            .I(port_address_c_4));
    InMux I__3751 (
            .O(N__16910),
            .I(N__16907));
    LocalMux I__3750 (
            .O(N__16907),
            .I(N__16904));
    Span12Mux_v I__3749 (
            .O(N__16904),
            .I(N__16901));
    Span12Mux_v I__3748 (
            .O(N__16901),
            .I(N__16898));
    Odrv12 I__3747 (
            .O(N__16898),
            .I(port_address_c_7));
    InMux I__3746 (
            .O(N__16895),
            .I(N__16888));
    InMux I__3745 (
            .O(N__16894),
            .I(N__16888));
    CascadeMux I__3744 (
            .O(N__16893),
            .I(N__16884));
    LocalMux I__3743 (
            .O(N__16888),
            .I(N__16881));
    InMux I__3742 (
            .O(N__16887),
            .I(N__16878));
    InMux I__3741 (
            .O(N__16884),
            .I(N__16875));
    Span4Mux_v I__3740 (
            .O(N__16881),
            .I(N__16870));
    LocalMux I__3739 (
            .O(N__16878),
            .I(N__16870));
    LocalMux I__3738 (
            .O(N__16875),
            .I(N__16867));
    Span4Mux_v I__3737 (
            .O(N__16870),
            .I(N__16864));
    Span12Mux_v I__3736 (
            .O(N__16867),
            .I(N__16859));
    Sp12to4 I__3735 (
            .O(N__16864),
            .I(N__16859));
    Span12Mux_h I__3734 (
            .O(N__16859),
            .I(N__16856));
    Odrv12 I__3733 (
            .O(N__16856),
            .I(port_enb_c));
    InMux I__3732 (
            .O(N__16853),
            .I(N__16850));
    LocalMux I__3731 (
            .O(N__16850),
            .I(N__16847));
    Span12Mux_v I__3730 (
            .O(N__16847),
            .I(N__16844));
    Odrv12 I__3729 (
            .O(N__16844),
            .I(port_address_c_2));
    InMux I__3728 (
            .O(N__16841),
            .I(N__16838));
    LocalMux I__3727 (
            .O(N__16838),
            .I(M_state_q_ns_1_0__m7Z0Z_5));
    CascadeMux I__3726 (
            .O(N__16835),
            .I(N__16831));
    CascadeMux I__3725 (
            .O(N__16834),
            .I(N__16827));
    InMux I__3724 (
            .O(N__16831),
            .I(N__16824));
    InMux I__3723 (
            .O(N__16830),
            .I(N__16821));
    InMux I__3722 (
            .O(N__16827),
            .I(N__16818));
    LocalMux I__3721 (
            .O(N__16824),
            .I(N__16815));
    LocalMux I__3720 (
            .O(N__16821),
            .I(N__16810));
    LocalMux I__3719 (
            .O(N__16818),
            .I(N__16810));
    Span4Mux_v I__3718 (
            .O(N__16815),
            .I(N__16807));
    Span4Mux_v I__3717 (
            .O(N__16810),
            .I(N__16804));
    Sp12to4 I__3716 (
            .O(N__16807),
            .I(N__16799));
    Sp12to4 I__3715 (
            .O(N__16804),
            .I(N__16799));
    Span12Mux_h I__3714 (
            .O(N__16799),
            .I(N__16796));
    Odrv12 I__3713 (
            .O(N__16796),
            .I(port_data_c_1));
    InMux I__3712 (
            .O(N__16793),
            .I(N__16790));
    LocalMux I__3711 (
            .O(N__16790),
            .I(N__16786));
    InMux I__3710 (
            .O(N__16789),
            .I(N__16783));
    Span4Mux_h I__3709 (
            .O(N__16786),
            .I(N__16779));
    LocalMux I__3708 (
            .O(N__16783),
            .I(N__16776));
    InMux I__3707 (
            .O(N__16782),
            .I(N__16773));
    Span4Mux_v I__3706 (
            .O(N__16779),
            .I(N__16767));
    Span4Mux_h I__3705 (
            .O(N__16776),
            .I(N__16767));
    LocalMux I__3704 (
            .O(N__16773),
            .I(N__16764));
    InMux I__3703 (
            .O(N__16772),
            .I(N__16761));
    Span4Mux_v I__3702 (
            .O(N__16767),
            .I(N__16755));
    Span4Mux_h I__3701 (
            .O(N__16764),
            .I(N__16755));
    LocalMux I__3700 (
            .O(N__16761),
            .I(N__16752));
    InMux I__3699 (
            .O(N__16760),
            .I(N__16749));
    Span4Mux_v I__3698 (
            .O(N__16755),
            .I(N__16742));
    Span4Mux_h I__3697 (
            .O(N__16752),
            .I(N__16742));
    LocalMux I__3696 (
            .O(N__16749),
            .I(N__16739));
    InMux I__3695 (
            .O(N__16748),
            .I(N__16736));
    InMux I__3694 (
            .O(N__16747),
            .I(N__16733));
    Span4Mux_v I__3693 (
            .O(N__16742),
            .I(N__16727));
    Span4Mux_h I__3692 (
            .O(N__16739),
            .I(N__16727));
    LocalMux I__3691 (
            .O(N__16736),
            .I(N__16724));
    LocalMux I__3690 (
            .O(N__16733),
            .I(N__16721));
    InMux I__3689 (
            .O(N__16732),
            .I(N__16718));
    Span4Mux_v I__3688 (
            .O(N__16727),
            .I(N__16713));
    Span4Mux_h I__3687 (
            .O(N__16724),
            .I(N__16713));
    Span4Mux_v I__3686 (
            .O(N__16721),
            .I(N__16708));
    LocalMux I__3685 (
            .O(N__16718),
            .I(N__16708));
    Odrv4 I__3684 (
            .O(N__16713),
            .I(M_this_vram_write_data_1));
    Odrv4 I__3683 (
            .O(N__16708),
            .I(M_this_vram_write_data_1));
    InMux I__3682 (
            .O(N__16703),
            .I(N__16700));
    LocalMux I__3681 (
            .O(N__16700),
            .I(N__16697));
    Span4Mux_v I__3680 (
            .O(N__16697),
            .I(N__16694));
    Span4Mux_v I__3679 (
            .O(N__16694),
            .I(N__16691));
    Odrv4 I__3678 (
            .O(N__16691),
            .I(\this_vram.mem_out_bus2_1 ));
    InMux I__3677 (
            .O(N__16688),
            .I(N__16685));
    LocalMux I__3676 (
            .O(N__16685),
            .I(N__16682));
    Odrv4 I__3675 (
            .O(N__16682),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_17 ));
    InMux I__3674 (
            .O(N__16679),
            .I(N__16676));
    LocalMux I__3673 (
            .O(N__16676),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_18 ));
    InMux I__3672 (
            .O(N__16673),
            .I(N__16670));
    LocalMux I__3671 (
            .O(N__16670),
            .I(M_this_start_address_delay_out_0));
    CascadeMux I__3670 (
            .O(N__16667),
            .I(M_state_q_ns_1_0__N_24_mux_cascade_));
    CascadeMux I__3669 (
            .O(N__16664),
            .I(M_state_q_ns_1_0__N_10_cascade_));
    CascadeMux I__3668 (
            .O(N__16661),
            .I(N__16658));
    CascadeBuf I__3667 (
            .O(N__16658),
            .I(N__16655));
    CascadeMux I__3666 (
            .O(N__16655),
            .I(N__16652));
    CascadeBuf I__3665 (
            .O(N__16652),
            .I(N__16649));
    CascadeMux I__3664 (
            .O(N__16649),
            .I(N__16646));
    CascadeBuf I__3663 (
            .O(N__16646),
            .I(N__16643));
    CascadeMux I__3662 (
            .O(N__16643),
            .I(N__16640));
    CascadeBuf I__3661 (
            .O(N__16640),
            .I(N__16637));
    CascadeMux I__3660 (
            .O(N__16637),
            .I(N__16634));
    CascadeBuf I__3659 (
            .O(N__16634),
            .I(N__16631));
    CascadeMux I__3658 (
            .O(N__16631),
            .I(N__16628));
    CascadeBuf I__3657 (
            .O(N__16628),
            .I(N__16625));
    CascadeMux I__3656 (
            .O(N__16625),
            .I(N__16622));
    CascadeBuf I__3655 (
            .O(N__16622),
            .I(N__16619));
    CascadeMux I__3654 (
            .O(N__16619),
            .I(N__16616));
    CascadeBuf I__3653 (
            .O(N__16616),
            .I(N__16613));
    CascadeMux I__3652 (
            .O(N__16613),
            .I(N__16610));
    CascadeBuf I__3651 (
            .O(N__16610),
            .I(N__16607));
    CascadeMux I__3650 (
            .O(N__16607),
            .I(N__16604));
    CascadeBuf I__3649 (
            .O(N__16604),
            .I(N__16601));
    CascadeMux I__3648 (
            .O(N__16601),
            .I(N__16598));
    CascadeBuf I__3647 (
            .O(N__16598),
            .I(N__16595));
    CascadeMux I__3646 (
            .O(N__16595),
            .I(N__16592));
    CascadeBuf I__3645 (
            .O(N__16592),
            .I(N__16589));
    CascadeMux I__3644 (
            .O(N__16589),
            .I(N__16586));
    CascadeBuf I__3643 (
            .O(N__16586),
            .I(N__16583));
    CascadeMux I__3642 (
            .O(N__16583),
            .I(N__16580));
    CascadeBuf I__3641 (
            .O(N__16580),
            .I(N__16577));
    CascadeMux I__3640 (
            .O(N__16577),
            .I(N__16574));
    CascadeBuf I__3639 (
            .O(N__16574),
            .I(N__16571));
    CascadeMux I__3638 (
            .O(N__16571),
            .I(N__16568));
    InMux I__3637 (
            .O(N__16568),
            .I(N__16563));
    InMux I__3636 (
            .O(N__16567),
            .I(N__16560));
    InMux I__3635 (
            .O(N__16566),
            .I(N__16557));
    LocalMux I__3634 (
            .O(N__16563),
            .I(N__16554));
    LocalMux I__3633 (
            .O(N__16560),
            .I(N__16551));
    LocalMux I__3632 (
            .O(N__16557),
            .I(N__16546));
    Span12Mux_s7_v I__3631 (
            .O(N__16554),
            .I(N__16546));
    Odrv4 I__3630 (
            .O(N__16551),
            .I(M_current_address_qZ0Z_1));
    Odrv12 I__3629 (
            .O(N__16546),
            .I(M_current_address_qZ0Z_1));
    CascadeMux I__3628 (
            .O(N__16541),
            .I(N__16538));
    InMux I__3627 (
            .O(N__16538),
            .I(N__16535));
    LocalMux I__3626 (
            .O(N__16535),
            .I(N__16532));
    Odrv4 I__3625 (
            .O(N__16532),
            .I(\this_start_data_delay.this_edge_detector.N_211 ));
    CascadeMux I__3624 (
            .O(N__16529),
            .I(N__16526));
    CascadeBuf I__3623 (
            .O(N__16526),
            .I(N__16523));
    CascadeMux I__3622 (
            .O(N__16523),
            .I(N__16520));
    CascadeBuf I__3621 (
            .O(N__16520),
            .I(N__16517));
    CascadeMux I__3620 (
            .O(N__16517),
            .I(N__16514));
    CascadeBuf I__3619 (
            .O(N__16514),
            .I(N__16511));
    CascadeMux I__3618 (
            .O(N__16511),
            .I(N__16508));
    CascadeBuf I__3617 (
            .O(N__16508),
            .I(N__16505));
    CascadeMux I__3616 (
            .O(N__16505),
            .I(N__16502));
    CascadeBuf I__3615 (
            .O(N__16502),
            .I(N__16499));
    CascadeMux I__3614 (
            .O(N__16499),
            .I(N__16496));
    CascadeBuf I__3613 (
            .O(N__16496),
            .I(N__16493));
    CascadeMux I__3612 (
            .O(N__16493),
            .I(N__16490));
    CascadeBuf I__3611 (
            .O(N__16490),
            .I(N__16487));
    CascadeMux I__3610 (
            .O(N__16487),
            .I(N__16484));
    CascadeBuf I__3609 (
            .O(N__16484),
            .I(N__16481));
    CascadeMux I__3608 (
            .O(N__16481),
            .I(N__16478));
    CascadeBuf I__3607 (
            .O(N__16478),
            .I(N__16475));
    CascadeMux I__3606 (
            .O(N__16475),
            .I(N__16472));
    CascadeBuf I__3605 (
            .O(N__16472),
            .I(N__16469));
    CascadeMux I__3604 (
            .O(N__16469),
            .I(N__16466));
    CascadeBuf I__3603 (
            .O(N__16466),
            .I(N__16463));
    CascadeMux I__3602 (
            .O(N__16463),
            .I(N__16460));
    CascadeBuf I__3601 (
            .O(N__16460),
            .I(N__16457));
    CascadeMux I__3600 (
            .O(N__16457),
            .I(N__16454));
    CascadeBuf I__3599 (
            .O(N__16454),
            .I(N__16451));
    CascadeMux I__3598 (
            .O(N__16451),
            .I(N__16448));
    CascadeBuf I__3597 (
            .O(N__16448),
            .I(N__16445));
    CascadeMux I__3596 (
            .O(N__16445),
            .I(N__16442));
    CascadeBuf I__3595 (
            .O(N__16442),
            .I(N__16439));
    CascadeMux I__3594 (
            .O(N__16439),
            .I(N__16436));
    InMux I__3593 (
            .O(N__16436),
            .I(N__16433));
    LocalMux I__3592 (
            .O(N__16433),
            .I(N__16429));
    InMux I__3591 (
            .O(N__16432),
            .I(N__16426));
    Span4Mux_h I__3590 (
            .O(N__16429),
            .I(N__16423));
    LocalMux I__3589 (
            .O(N__16426),
            .I(N__16417));
    Span4Mux_v I__3588 (
            .O(N__16423),
            .I(N__16417));
    InMux I__3587 (
            .O(N__16422),
            .I(N__16414));
    Span4Mux_v I__3586 (
            .O(N__16417),
            .I(N__16411));
    LocalMux I__3585 (
            .O(N__16414),
            .I(M_current_address_qZ0Z_4));
    Odrv4 I__3584 (
            .O(N__16411),
            .I(M_current_address_qZ0Z_4));
    InMux I__3583 (
            .O(N__16406),
            .I(N__16402));
    CascadeMux I__3582 (
            .O(N__16405),
            .I(N__16399));
    LocalMux I__3581 (
            .O(N__16402),
            .I(N__16396));
    InMux I__3580 (
            .O(N__16399),
            .I(N__16393));
    Span4Mux_v I__3579 (
            .O(N__16396),
            .I(N__16390));
    LocalMux I__3578 (
            .O(N__16393),
            .I(N__16387));
    Span4Mux_h I__3577 (
            .O(N__16390),
            .I(N__16384));
    Sp12to4 I__3576 (
            .O(N__16387),
            .I(N__16381));
    Span4Mux_h I__3575 (
            .O(N__16384),
            .I(N__16378));
    Span12Mux_v I__3574 (
            .O(N__16381),
            .I(N__16375));
    Odrv4 I__3573 (
            .O(N__16378),
            .I(port_data_c_4));
    Odrv12 I__3572 (
            .O(N__16375),
            .I(port_data_c_4));
    CascadeMux I__3571 (
            .O(N__16370),
            .I(N__16367));
    InMux I__3570 (
            .O(N__16367),
            .I(N__16364));
    LocalMux I__3569 (
            .O(N__16364),
            .I(N__16361));
    Span4Mux_v I__3568 (
            .O(N__16361),
            .I(N__16358));
    Odrv4 I__3567 (
            .O(N__16358),
            .I(\this_start_data_delay.this_edge_detector.N_214 ));
    InMux I__3566 (
            .O(N__16355),
            .I(N__16352));
    LocalMux I__3565 (
            .O(N__16352),
            .I(N__16348));
    InMux I__3564 (
            .O(N__16351),
            .I(N__16345));
    Span4Mux_h I__3563 (
            .O(N__16348),
            .I(N__16327));
    LocalMux I__3562 (
            .O(N__16345),
            .I(N__16327));
    InMux I__3561 (
            .O(N__16344),
            .I(N__16322));
    InMux I__3560 (
            .O(N__16343),
            .I(N__16322));
    InMux I__3559 (
            .O(N__16342),
            .I(N__16315));
    InMux I__3558 (
            .O(N__16341),
            .I(N__16315));
    InMux I__3557 (
            .O(N__16340),
            .I(N__16315));
    InMux I__3556 (
            .O(N__16339),
            .I(N__16312));
    InMux I__3555 (
            .O(N__16338),
            .I(N__16309));
    InMux I__3554 (
            .O(N__16337),
            .I(N__16302));
    InMux I__3553 (
            .O(N__16336),
            .I(N__16302));
    InMux I__3552 (
            .O(N__16335),
            .I(N__16302));
    InMux I__3551 (
            .O(N__16334),
            .I(N__16297));
    InMux I__3550 (
            .O(N__16333),
            .I(N__16297));
    InMux I__3549 (
            .O(N__16332),
            .I(N__16276));
    Span4Mux_h I__3548 (
            .O(N__16327),
            .I(N__16265));
    LocalMux I__3547 (
            .O(N__16322),
            .I(N__16265));
    LocalMux I__3546 (
            .O(N__16315),
            .I(N__16265));
    LocalMux I__3545 (
            .O(N__16312),
            .I(N__16265));
    LocalMux I__3544 (
            .O(N__16309),
            .I(N__16265));
    LocalMux I__3543 (
            .O(N__16302),
            .I(N__16260));
    LocalMux I__3542 (
            .O(N__16297),
            .I(N__16260));
    InMux I__3541 (
            .O(N__16296),
            .I(N__16257));
    InMux I__3540 (
            .O(N__16295),
            .I(N__16246));
    InMux I__3539 (
            .O(N__16294),
            .I(N__16246));
    InMux I__3538 (
            .O(N__16293),
            .I(N__16246));
    InMux I__3537 (
            .O(N__16292),
            .I(N__16246));
    InMux I__3536 (
            .O(N__16291),
            .I(N__16246));
    InMux I__3535 (
            .O(N__16290),
            .I(N__16243));
    InMux I__3534 (
            .O(N__16289),
            .I(N__16236));
    InMux I__3533 (
            .O(N__16288),
            .I(N__16236));
    InMux I__3532 (
            .O(N__16287),
            .I(N__16236));
    InMux I__3531 (
            .O(N__16286),
            .I(N__16229));
    InMux I__3530 (
            .O(N__16285),
            .I(N__16229));
    InMux I__3529 (
            .O(N__16284),
            .I(N__16229));
    InMux I__3528 (
            .O(N__16283),
            .I(N__16222));
    InMux I__3527 (
            .O(N__16282),
            .I(N__16222));
    InMux I__3526 (
            .O(N__16281),
            .I(N__16222));
    InMux I__3525 (
            .O(N__16280),
            .I(N__16217));
    InMux I__3524 (
            .O(N__16279),
            .I(N__16217));
    LocalMux I__3523 (
            .O(N__16276),
            .I(N__16214));
    Span4Mux_v I__3522 (
            .O(N__16265),
            .I(N__16207));
    Span4Mux_v I__3521 (
            .O(N__16260),
            .I(N__16207));
    LocalMux I__3520 (
            .O(N__16257),
            .I(N__16207));
    LocalMux I__3519 (
            .O(N__16246),
            .I(M_state_qZ0Z_0));
    LocalMux I__3518 (
            .O(N__16243),
            .I(M_state_qZ0Z_0));
    LocalMux I__3517 (
            .O(N__16236),
            .I(M_state_qZ0Z_0));
    LocalMux I__3516 (
            .O(N__16229),
            .I(M_state_qZ0Z_0));
    LocalMux I__3515 (
            .O(N__16222),
            .I(M_state_qZ0Z_0));
    LocalMux I__3514 (
            .O(N__16217),
            .I(M_state_qZ0Z_0));
    Odrv4 I__3513 (
            .O(N__16214),
            .I(M_state_qZ0Z_0));
    Odrv4 I__3512 (
            .O(N__16207),
            .I(M_state_qZ0Z_0));
    InMux I__3511 (
            .O(N__16190),
            .I(N__16187));
    LocalMux I__3510 (
            .O(N__16187),
            .I(N__16184));
    Span12Mux_h I__3509 (
            .O(N__16184),
            .I(N__16181));
    Odrv12 I__3508 (
            .O(N__16181),
            .I(port_address_c_1));
    CascadeMux I__3507 (
            .O(N__16178),
            .I(N__16175));
    InMux I__3506 (
            .O(N__16175),
            .I(N__16172));
    LocalMux I__3505 (
            .O(N__16172),
            .I(M_state_q_ns_1_0__N_24_mux));
    InMux I__3504 (
            .O(N__16169),
            .I(N__16166));
    LocalMux I__3503 (
            .O(N__16166),
            .I(N__16162));
    InMux I__3502 (
            .O(N__16165),
            .I(N__16159));
    Span4Mux_v I__3501 (
            .O(N__16162),
            .I(N__16154));
    LocalMux I__3500 (
            .O(N__16159),
            .I(N__16154));
    Sp12to4 I__3499 (
            .O(N__16154),
            .I(N__16151));
    Span12Mux_h I__3498 (
            .O(N__16151),
            .I(N__16148));
    Odrv12 I__3497 (
            .O(N__16148),
            .I(port_address_c_0));
    CascadeMux I__3496 (
            .O(N__16145),
            .I(N__16142));
    CascadeBuf I__3495 (
            .O(N__16142),
            .I(N__16139));
    CascadeMux I__3494 (
            .O(N__16139),
            .I(N__16136));
    CascadeBuf I__3493 (
            .O(N__16136),
            .I(N__16133));
    CascadeMux I__3492 (
            .O(N__16133),
            .I(N__16130));
    CascadeBuf I__3491 (
            .O(N__16130),
            .I(N__16127));
    CascadeMux I__3490 (
            .O(N__16127),
            .I(N__16124));
    CascadeBuf I__3489 (
            .O(N__16124),
            .I(N__16121));
    CascadeMux I__3488 (
            .O(N__16121),
            .I(N__16118));
    CascadeBuf I__3487 (
            .O(N__16118),
            .I(N__16115));
    CascadeMux I__3486 (
            .O(N__16115),
            .I(N__16112));
    CascadeBuf I__3485 (
            .O(N__16112),
            .I(N__16109));
    CascadeMux I__3484 (
            .O(N__16109),
            .I(N__16106));
    CascadeBuf I__3483 (
            .O(N__16106),
            .I(N__16103));
    CascadeMux I__3482 (
            .O(N__16103),
            .I(N__16100));
    CascadeBuf I__3481 (
            .O(N__16100),
            .I(N__16097));
    CascadeMux I__3480 (
            .O(N__16097),
            .I(N__16094));
    CascadeBuf I__3479 (
            .O(N__16094),
            .I(N__16091));
    CascadeMux I__3478 (
            .O(N__16091),
            .I(N__16088));
    CascadeBuf I__3477 (
            .O(N__16088),
            .I(N__16085));
    CascadeMux I__3476 (
            .O(N__16085),
            .I(N__16082));
    CascadeBuf I__3475 (
            .O(N__16082),
            .I(N__16079));
    CascadeMux I__3474 (
            .O(N__16079),
            .I(N__16076));
    CascadeBuf I__3473 (
            .O(N__16076),
            .I(N__16073));
    CascadeMux I__3472 (
            .O(N__16073),
            .I(N__16070));
    CascadeBuf I__3471 (
            .O(N__16070),
            .I(N__16067));
    CascadeMux I__3470 (
            .O(N__16067),
            .I(N__16064));
    CascadeBuf I__3469 (
            .O(N__16064),
            .I(N__16061));
    CascadeMux I__3468 (
            .O(N__16061),
            .I(N__16058));
    CascadeBuf I__3467 (
            .O(N__16058),
            .I(N__16055));
    CascadeMux I__3466 (
            .O(N__16055),
            .I(N__16052));
    InMux I__3465 (
            .O(N__16052),
            .I(N__16049));
    LocalMux I__3464 (
            .O(N__16049),
            .I(N__16046));
    Span4Mux_v I__3463 (
            .O(N__16046),
            .I(N__16042));
    InMux I__3462 (
            .O(N__16045),
            .I(N__16038));
    Span4Mux_h I__3461 (
            .O(N__16042),
            .I(N__16035));
    InMux I__3460 (
            .O(N__16041),
            .I(N__16032));
    LocalMux I__3459 (
            .O(N__16038),
            .I(N__16027));
    Span4Mux_v I__3458 (
            .O(N__16035),
            .I(N__16027));
    LocalMux I__3457 (
            .O(N__16032),
            .I(M_current_address_qZ0Z_8));
    Odrv4 I__3456 (
            .O(N__16027),
            .I(M_current_address_qZ0Z_8));
    InMux I__3455 (
            .O(N__16022),
            .I(N__16019));
    LocalMux I__3454 (
            .O(N__16019),
            .I(N__16016));
    Odrv4 I__3453 (
            .O(N__16016),
            .I(\this_start_data_delay.this_edge_detector.N_218 ));
    CascadeMux I__3452 (
            .O(N__16013),
            .I(N__16010));
    CascadeBuf I__3451 (
            .O(N__16010),
            .I(N__16007));
    CascadeMux I__3450 (
            .O(N__16007),
            .I(N__16004));
    CascadeBuf I__3449 (
            .O(N__16004),
            .I(N__16001));
    CascadeMux I__3448 (
            .O(N__16001),
            .I(N__15998));
    CascadeBuf I__3447 (
            .O(N__15998),
            .I(N__15995));
    CascadeMux I__3446 (
            .O(N__15995),
            .I(N__15992));
    CascadeBuf I__3445 (
            .O(N__15992),
            .I(N__15989));
    CascadeMux I__3444 (
            .O(N__15989),
            .I(N__15986));
    CascadeBuf I__3443 (
            .O(N__15986),
            .I(N__15983));
    CascadeMux I__3442 (
            .O(N__15983),
            .I(N__15980));
    CascadeBuf I__3441 (
            .O(N__15980),
            .I(N__15977));
    CascadeMux I__3440 (
            .O(N__15977),
            .I(N__15974));
    CascadeBuf I__3439 (
            .O(N__15974),
            .I(N__15971));
    CascadeMux I__3438 (
            .O(N__15971),
            .I(N__15968));
    CascadeBuf I__3437 (
            .O(N__15968),
            .I(N__15965));
    CascadeMux I__3436 (
            .O(N__15965),
            .I(N__15962));
    CascadeBuf I__3435 (
            .O(N__15962),
            .I(N__15959));
    CascadeMux I__3434 (
            .O(N__15959),
            .I(N__15956));
    CascadeBuf I__3433 (
            .O(N__15956),
            .I(N__15953));
    CascadeMux I__3432 (
            .O(N__15953),
            .I(N__15950));
    CascadeBuf I__3431 (
            .O(N__15950),
            .I(N__15947));
    CascadeMux I__3430 (
            .O(N__15947),
            .I(N__15944));
    CascadeBuf I__3429 (
            .O(N__15944),
            .I(N__15941));
    CascadeMux I__3428 (
            .O(N__15941),
            .I(N__15938));
    CascadeBuf I__3427 (
            .O(N__15938),
            .I(N__15935));
    CascadeMux I__3426 (
            .O(N__15935),
            .I(N__15932));
    CascadeBuf I__3425 (
            .O(N__15932),
            .I(N__15929));
    CascadeMux I__3424 (
            .O(N__15929),
            .I(N__15926));
    CascadeBuf I__3423 (
            .O(N__15926),
            .I(N__15923));
    CascadeMux I__3422 (
            .O(N__15923),
            .I(N__15920));
    InMux I__3421 (
            .O(N__15920),
            .I(N__15917));
    LocalMux I__3420 (
            .O(N__15917),
            .I(N__15914));
    Span4Mux_s3_v I__3419 (
            .O(N__15914),
            .I(N__15910));
    InMux I__3418 (
            .O(N__15913),
            .I(N__15906));
    Span4Mux_h I__3417 (
            .O(N__15910),
            .I(N__15903));
    InMux I__3416 (
            .O(N__15909),
            .I(N__15900));
    LocalMux I__3415 (
            .O(N__15906),
            .I(N__15895));
    Span4Mux_v I__3414 (
            .O(N__15903),
            .I(N__15895));
    LocalMux I__3413 (
            .O(N__15900),
            .I(M_current_address_qZ0Z_10));
    Odrv4 I__3412 (
            .O(N__15895),
            .I(M_current_address_qZ0Z_10));
    CascadeMux I__3411 (
            .O(N__15890),
            .I(N__15887));
    InMux I__3410 (
            .O(N__15887),
            .I(N__15884));
    LocalMux I__3409 (
            .O(N__15884),
            .I(\this_start_data_delay.this_edge_detector.N_220 ));
    CascadeMux I__3408 (
            .O(N__15881),
            .I(N__15878));
    InMux I__3407 (
            .O(N__15878),
            .I(N__15875));
    LocalMux I__3406 (
            .O(N__15875),
            .I(N__15872));
    Odrv4 I__3405 (
            .O(N__15872),
            .I(\this_start_data_delay.this_edge_detector.N_221 ));
    CascadeMux I__3404 (
            .O(N__15869),
            .I(N__15865));
    InMux I__3403 (
            .O(N__15868),
            .I(N__15862));
    InMux I__3402 (
            .O(N__15865),
            .I(N__15859));
    LocalMux I__3401 (
            .O(N__15862),
            .I(N__15854));
    LocalMux I__3400 (
            .O(N__15859),
            .I(N__15854));
    Span12Mux_s9_v I__3399 (
            .O(N__15854),
            .I(N__15851));
    Span12Mux_v I__3398 (
            .O(N__15851),
            .I(N__15848));
    Span12Mux_h I__3397 (
            .O(N__15848),
            .I(N__15845));
    Odrv12 I__3396 (
            .O(N__15845),
            .I(port_data_c_6));
    CascadeMux I__3395 (
            .O(N__15842),
            .I(N__15839));
    InMux I__3394 (
            .O(N__15839),
            .I(N__15836));
    LocalMux I__3393 (
            .O(N__15836),
            .I(\this_start_data_delay.this_edge_detector.N_223 ));
    InMux I__3392 (
            .O(N__15833),
            .I(N__15830));
    LocalMux I__3391 (
            .O(N__15830),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_15 ));
    InMux I__3390 (
            .O(N__15827),
            .I(N__15824));
    LocalMux I__3389 (
            .O(N__15824),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_16 ));
    CascadeMux I__3388 (
            .O(N__15821),
            .I(N__15818));
    CascadeBuf I__3387 (
            .O(N__15818),
            .I(N__15815));
    CascadeMux I__3386 (
            .O(N__15815),
            .I(N__15812));
    CascadeBuf I__3385 (
            .O(N__15812),
            .I(N__15809));
    CascadeMux I__3384 (
            .O(N__15809),
            .I(N__15806));
    CascadeBuf I__3383 (
            .O(N__15806),
            .I(N__15803));
    CascadeMux I__3382 (
            .O(N__15803),
            .I(N__15800));
    CascadeBuf I__3381 (
            .O(N__15800),
            .I(N__15797));
    CascadeMux I__3380 (
            .O(N__15797),
            .I(N__15794));
    CascadeBuf I__3379 (
            .O(N__15794),
            .I(N__15791));
    CascadeMux I__3378 (
            .O(N__15791),
            .I(N__15788));
    CascadeBuf I__3377 (
            .O(N__15788),
            .I(N__15785));
    CascadeMux I__3376 (
            .O(N__15785),
            .I(N__15782));
    CascadeBuf I__3375 (
            .O(N__15782),
            .I(N__15779));
    CascadeMux I__3374 (
            .O(N__15779),
            .I(N__15776));
    CascadeBuf I__3373 (
            .O(N__15776),
            .I(N__15773));
    CascadeMux I__3372 (
            .O(N__15773),
            .I(N__15770));
    CascadeBuf I__3371 (
            .O(N__15770),
            .I(N__15767));
    CascadeMux I__3370 (
            .O(N__15767),
            .I(N__15764));
    CascadeBuf I__3369 (
            .O(N__15764),
            .I(N__15761));
    CascadeMux I__3368 (
            .O(N__15761),
            .I(N__15758));
    CascadeBuf I__3367 (
            .O(N__15758),
            .I(N__15755));
    CascadeMux I__3366 (
            .O(N__15755),
            .I(N__15752));
    CascadeBuf I__3365 (
            .O(N__15752),
            .I(N__15749));
    CascadeMux I__3364 (
            .O(N__15749),
            .I(N__15746));
    CascadeBuf I__3363 (
            .O(N__15746),
            .I(N__15743));
    CascadeMux I__3362 (
            .O(N__15743),
            .I(N__15740));
    CascadeBuf I__3361 (
            .O(N__15740),
            .I(N__15737));
    CascadeMux I__3360 (
            .O(N__15737),
            .I(N__15734));
    CascadeBuf I__3359 (
            .O(N__15734),
            .I(N__15731));
    CascadeMux I__3358 (
            .O(N__15731),
            .I(N__15728));
    InMux I__3357 (
            .O(N__15728),
            .I(N__15725));
    LocalMux I__3356 (
            .O(N__15725),
            .I(N__15722));
    Span4Mux_s2_v I__3355 (
            .O(N__15722),
            .I(N__15718));
    CascadeMux I__3354 (
            .O(N__15721),
            .I(N__15715));
    Span4Mux_h I__3353 (
            .O(N__15718),
            .I(N__15711));
    InMux I__3352 (
            .O(N__15715),
            .I(N__15708));
    InMux I__3351 (
            .O(N__15714),
            .I(N__15705));
    Span4Mux_v I__3350 (
            .O(N__15711),
            .I(N__15702));
    LocalMux I__3349 (
            .O(N__15708),
            .I(M_current_address_qZ0Z_7));
    LocalMux I__3348 (
            .O(N__15705),
            .I(M_current_address_qZ0Z_7));
    Odrv4 I__3347 (
            .O(N__15702),
            .I(M_current_address_qZ0Z_7));
    CascadeMux I__3346 (
            .O(N__15695),
            .I(N__15692));
    InMux I__3345 (
            .O(N__15692),
            .I(N__15689));
    LocalMux I__3344 (
            .O(N__15689),
            .I(\this_start_data_delay.this_edge_detector.N_217 ));
    CascadeMux I__3343 (
            .O(N__15686),
            .I(N__15683));
    CascadeBuf I__3342 (
            .O(N__15683),
            .I(N__15680));
    CascadeMux I__3341 (
            .O(N__15680),
            .I(N__15677));
    CascadeBuf I__3340 (
            .O(N__15677),
            .I(N__15674));
    CascadeMux I__3339 (
            .O(N__15674),
            .I(N__15671));
    CascadeBuf I__3338 (
            .O(N__15671),
            .I(N__15668));
    CascadeMux I__3337 (
            .O(N__15668),
            .I(N__15665));
    CascadeBuf I__3336 (
            .O(N__15665),
            .I(N__15662));
    CascadeMux I__3335 (
            .O(N__15662),
            .I(N__15659));
    CascadeBuf I__3334 (
            .O(N__15659),
            .I(N__15656));
    CascadeMux I__3333 (
            .O(N__15656),
            .I(N__15653));
    CascadeBuf I__3332 (
            .O(N__15653),
            .I(N__15650));
    CascadeMux I__3331 (
            .O(N__15650),
            .I(N__15647));
    CascadeBuf I__3330 (
            .O(N__15647),
            .I(N__15644));
    CascadeMux I__3329 (
            .O(N__15644),
            .I(N__15641));
    CascadeBuf I__3328 (
            .O(N__15641),
            .I(N__15638));
    CascadeMux I__3327 (
            .O(N__15638),
            .I(N__15635));
    CascadeBuf I__3326 (
            .O(N__15635),
            .I(N__15632));
    CascadeMux I__3325 (
            .O(N__15632),
            .I(N__15629));
    CascadeBuf I__3324 (
            .O(N__15629),
            .I(N__15626));
    CascadeMux I__3323 (
            .O(N__15626),
            .I(N__15623));
    CascadeBuf I__3322 (
            .O(N__15623),
            .I(N__15620));
    CascadeMux I__3321 (
            .O(N__15620),
            .I(N__15617));
    CascadeBuf I__3320 (
            .O(N__15617),
            .I(N__15614));
    CascadeMux I__3319 (
            .O(N__15614),
            .I(N__15611));
    CascadeBuf I__3318 (
            .O(N__15611),
            .I(N__15608));
    CascadeMux I__3317 (
            .O(N__15608),
            .I(N__15605));
    CascadeBuf I__3316 (
            .O(N__15605),
            .I(N__15602));
    CascadeMux I__3315 (
            .O(N__15602),
            .I(N__15599));
    CascadeBuf I__3314 (
            .O(N__15599),
            .I(N__15596));
    CascadeMux I__3313 (
            .O(N__15596),
            .I(N__15593));
    InMux I__3312 (
            .O(N__15593),
            .I(N__15590));
    LocalMux I__3311 (
            .O(N__15590),
            .I(N__15587));
    Span4Mux_s3_v I__3310 (
            .O(N__15587),
            .I(N__15584));
    Span4Mux_h I__3309 (
            .O(N__15584),
            .I(N__15579));
    InMux I__3308 (
            .O(N__15583),
            .I(N__15576));
    InMux I__3307 (
            .O(N__15582),
            .I(N__15573));
    Span4Mux_v I__3306 (
            .O(N__15579),
            .I(N__15570));
    LocalMux I__3305 (
            .O(N__15576),
            .I(M_current_address_qZ0Z_0));
    LocalMux I__3304 (
            .O(N__15573),
            .I(M_current_address_qZ0Z_0));
    Odrv4 I__3303 (
            .O(N__15570),
            .I(M_current_address_qZ0Z_0));
    CascadeMux I__3302 (
            .O(N__15563),
            .I(N__15560));
    InMux I__3301 (
            .O(N__15560),
            .I(N__15557));
    LocalMux I__3300 (
            .O(N__15557),
            .I(\this_start_data_delay.this_edge_detector.N_210 ));
    InMux I__3299 (
            .O(N__15554),
            .I(N__15551));
    LocalMux I__3298 (
            .O(N__15551),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_13 ));
    InMux I__3297 (
            .O(N__15548),
            .I(N__15545));
    LocalMux I__3296 (
            .O(N__15545),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_14 ));
    InMux I__3295 (
            .O(N__15542),
            .I(N__15539));
    LocalMux I__3294 (
            .O(N__15539),
            .I(M_current_address_q_RNIHDTUZ0Z_0));
    InMux I__3293 (
            .O(N__15536),
            .I(N__15533));
    LocalMux I__3292 (
            .O(N__15533),
            .I(un1_M_current_address_q_cry_5_c_RNIC9GNZ0));
    InMux I__3291 (
            .O(N__15530),
            .I(N__15527));
    LocalMux I__3290 (
            .O(N__15527),
            .I(un1_M_current_address_q_cry_6_c_RNIECHNZ0));
    InMux I__3289 (
            .O(N__15524),
            .I(N__15521));
    LocalMux I__3288 (
            .O(N__15521),
            .I(un1_M_current_address_q_cry_10_c_RNI4KKHZ0));
    InMux I__3287 (
            .O(N__15518),
            .I(N__15515));
    LocalMux I__3286 (
            .O(N__15515),
            .I(un1_M_current_address_q_cry_2_c_RNI60DNZ0));
    InMux I__3285 (
            .O(N__15512),
            .I(N__15500));
    InMux I__3284 (
            .O(N__15511),
            .I(N__15497));
    InMux I__3283 (
            .O(N__15510),
            .I(N__15494));
    InMux I__3282 (
            .O(N__15509),
            .I(N__15491));
    InMux I__3281 (
            .O(N__15508),
            .I(N__15488));
    InMux I__3280 (
            .O(N__15507),
            .I(N__15485));
    InMux I__3279 (
            .O(N__15506),
            .I(N__15480));
    InMux I__3278 (
            .O(N__15505),
            .I(N__15480));
    InMux I__3277 (
            .O(N__15504),
            .I(N__15477));
    InMux I__3276 (
            .O(N__15503),
            .I(N__15474));
    LocalMux I__3275 (
            .O(N__15500),
            .I(N__15459));
    LocalMux I__3274 (
            .O(N__15497),
            .I(N__15456));
    LocalMux I__3273 (
            .O(N__15494),
            .I(N__15453));
    LocalMux I__3272 (
            .O(N__15491),
            .I(N__15450));
    LocalMux I__3271 (
            .O(N__15488),
            .I(N__15447));
    LocalMux I__3270 (
            .O(N__15485),
            .I(N__15444));
    LocalMux I__3269 (
            .O(N__15480),
            .I(N__15441));
    LocalMux I__3268 (
            .O(N__15477),
            .I(N__15438));
    LocalMux I__3267 (
            .O(N__15474),
            .I(N__15435));
    SRMux I__3266 (
            .O(N__15473),
            .I(N__15392));
    SRMux I__3265 (
            .O(N__15472),
            .I(N__15392));
    SRMux I__3264 (
            .O(N__15471),
            .I(N__15392));
    SRMux I__3263 (
            .O(N__15470),
            .I(N__15392));
    SRMux I__3262 (
            .O(N__15469),
            .I(N__15392));
    SRMux I__3261 (
            .O(N__15468),
            .I(N__15392));
    SRMux I__3260 (
            .O(N__15467),
            .I(N__15392));
    SRMux I__3259 (
            .O(N__15466),
            .I(N__15392));
    SRMux I__3258 (
            .O(N__15465),
            .I(N__15392));
    SRMux I__3257 (
            .O(N__15464),
            .I(N__15392));
    SRMux I__3256 (
            .O(N__15463),
            .I(N__15392));
    SRMux I__3255 (
            .O(N__15462),
            .I(N__15392));
    Glb2LocalMux I__3254 (
            .O(N__15459),
            .I(N__15392));
    Glb2LocalMux I__3253 (
            .O(N__15456),
            .I(N__15392));
    Glb2LocalMux I__3252 (
            .O(N__15453),
            .I(N__15392));
    Glb2LocalMux I__3251 (
            .O(N__15450),
            .I(N__15392));
    Glb2LocalMux I__3250 (
            .O(N__15447),
            .I(N__15392));
    Glb2LocalMux I__3249 (
            .O(N__15444),
            .I(N__15392));
    Glb2LocalMux I__3248 (
            .O(N__15441),
            .I(N__15392));
    Glb2LocalMux I__3247 (
            .O(N__15438),
            .I(N__15392));
    Glb2LocalMux I__3246 (
            .O(N__15435),
            .I(N__15392));
    GlobalMux I__3245 (
            .O(N__15392),
            .I(N__15389));
    gio2CtrlBuf I__3244 (
            .O(N__15389),
            .I(N_339_g));
    CascadeMux I__3243 (
            .O(N__15386),
            .I(N__15383));
    CascadeBuf I__3242 (
            .O(N__15383),
            .I(N__15380));
    CascadeMux I__3241 (
            .O(N__15380),
            .I(N__15377));
    CascadeBuf I__3240 (
            .O(N__15377),
            .I(N__15374));
    CascadeMux I__3239 (
            .O(N__15374),
            .I(N__15371));
    CascadeBuf I__3238 (
            .O(N__15371),
            .I(N__15368));
    CascadeMux I__3237 (
            .O(N__15368),
            .I(N__15365));
    CascadeBuf I__3236 (
            .O(N__15365),
            .I(N__15362));
    CascadeMux I__3235 (
            .O(N__15362),
            .I(N__15359));
    CascadeBuf I__3234 (
            .O(N__15359),
            .I(N__15356));
    CascadeMux I__3233 (
            .O(N__15356),
            .I(N__15353));
    CascadeBuf I__3232 (
            .O(N__15353),
            .I(N__15350));
    CascadeMux I__3231 (
            .O(N__15350),
            .I(N__15347));
    CascadeBuf I__3230 (
            .O(N__15347),
            .I(N__15344));
    CascadeMux I__3229 (
            .O(N__15344),
            .I(N__15341));
    CascadeBuf I__3228 (
            .O(N__15341),
            .I(N__15338));
    CascadeMux I__3227 (
            .O(N__15338),
            .I(N__15335));
    CascadeBuf I__3226 (
            .O(N__15335),
            .I(N__15332));
    CascadeMux I__3225 (
            .O(N__15332),
            .I(N__15329));
    CascadeBuf I__3224 (
            .O(N__15329),
            .I(N__15326));
    CascadeMux I__3223 (
            .O(N__15326),
            .I(N__15323));
    CascadeBuf I__3222 (
            .O(N__15323),
            .I(N__15320));
    CascadeMux I__3221 (
            .O(N__15320),
            .I(N__15317));
    CascadeBuf I__3220 (
            .O(N__15317),
            .I(N__15314));
    CascadeMux I__3219 (
            .O(N__15314),
            .I(N__15311));
    CascadeBuf I__3218 (
            .O(N__15311),
            .I(N__15308));
    CascadeMux I__3217 (
            .O(N__15308),
            .I(N__15305));
    CascadeBuf I__3216 (
            .O(N__15305),
            .I(N__15302));
    CascadeMux I__3215 (
            .O(N__15302),
            .I(N__15299));
    CascadeBuf I__3214 (
            .O(N__15299),
            .I(N__15296));
    CascadeMux I__3213 (
            .O(N__15296),
            .I(N__15293));
    InMux I__3212 (
            .O(N__15293),
            .I(N__15290));
    LocalMux I__3211 (
            .O(N__15290),
            .I(N__15285));
    InMux I__3210 (
            .O(N__15289),
            .I(N__15282));
    InMux I__3209 (
            .O(N__15288),
            .I(N__15279));
    Span12Mux_h I__3208 (
            .O(N__15285),
            .I(N__15276));
    LocalMux I__3207 (
            .O(N__15282),
            .I(M_current_address_qZ0Z_6));
    LocalMux I__3206 (
            .O(N__15279),
            .I(M_current_address_qZ0Z_6));
    Odrv12 I__3205 (
            .O(N__15276),
            .I(M_current_address_qZ0Z_6));
    InMux I__3204 (
            .O(N__15269),
            .I(N__15266));
    LocalMux I__3203 (
            .O(N__15266),
            .I(\this_start_data_delay.this_edge_detector.N_216 ));
    CascadeMux I__3202 (
            .O(N__15263),
            .I(N__15260));
    CascadeBuf I__3201 (
            .O(N__15260),
            .I(N__15257));
    CascadeMux I__3200 (
            .O(N__15257),
            .I(N__15254));
    CascadeBuf I__3199 (
            .O(N__15254),
            .I(N__15251));
    CascadeMux I__3198 (
            .O(N__15251),
            .I(N__15248));
    CascadeBuf I__3197 (
            .O(N__15248),
            .I(N__15245));
    CascadeMux I__3196 (
            .O(N__15245),
            .I(N__15242));
    CascadeBuf I__3195 (
            .O(N__15242),
            .I(N__15239));
    CascadeMux I__3194 (
            .O(N__15239),
            .I(N__15236));
    CascadeBuf I__3193 (
            .O(N__15236),
            .I(N__15233));
    CascadeMux I__3192 (
            .O(N__15233),
            .I(N__15230));
    CascadeBuf I__3191 (
            .O(N__15230),
            .I(N__15227));
    CascadeMux I__3190 (
            .O(N__15227),
            .I(N__15224));
    CascadeBuf I__3189 (
            .O(N__15224),
            .I(N__15221));
    CascadeMux I__3188 (
            .O(N__15221),
            .I(N__15218));
    CascadeBuf I__3187 (
            .O(N__15218),
            .I(N__15215));
    CascadeMux I__3186 (
            .O(N__15215),
            .I(N__15212));
    CascadeBuf I__3185 (
            .O(N__15212),
            .I(N__15209));
    CascadeMux I__3184 (
            .O(N__15209),
            .I(N__15206));
    CascadeBuf I__3183 (
            .O(N__15206),
            .I(N__15203));
    CascadeMux I__3182 (
            .O(N__15203),
            .I(N__15200));
    CascadeBuf I__3181 (
            .O(N__15200),
            .I(N__15197));
    CascadeMux I__3180 (
            .O(N__15197),
            .I(N__15194));
    CascadeBuf I__3179 (
            .O(N__15194),
            .I(N__15191));
    CascadeMux I__3178 (
            .O(N__15191),
            .I(N__15188));
    CascadeBuf I__3177 (
            .O(N__15188),
            .I(N__15185));
    CascadeMux I__3176 (
            .O(N__15185),
            .I(N__15182));
    CascadeBuf I__3175 (
            .O(N__15182),
            .I(N__15179));
    CascadeMux I__3174 (
            .O(N__15179),
            .I(N__15176));
    CascadeBuf I__3173 (
            .O(N__15176),
            .I(N__15173));
    CascadeMux I__3172 (
            .O(N__15173),
            .I(N__15170));
    InMux I__3171 (
            .O(N__15170),
            .I(N__15167));
    LocalMux I__3170 (
            .O(N__15167),
            .I(N__15164));
    Span4Mux_s2_v I__3169 (
            .O(N__15164),
            .I(N__15161));
    Span4Mux_h I__3168 (
            .O(N__15161),
            .I(N__15156));
    InMux I__3167 (
            .O(N__15160),
            .I(N__15153));
    InMux I__3166 (
            .O(N__15159),
            .I(N__15150));
    Span4Mux_v I__3165 (
            .O(N__15156),
            .I(N__15147));
    LocalMux I__3164 (
            .O(N__15153),
            .I(M_current_address_qZ0Z_3));
    LocalMux I__3163 (
            .O(N__15150),
            .I(M_current_address_qZ0Z_3));
    Odrv4 I__3162 (
            .O(N__15147),
            .I(M_current_address_qZ0Z_3));
    CascadeMux I__3161 (
            .O(N__15140),
            .I(N__15137));
    InMux I__3160 (
            .O(N__15137),
            .I(N__15134));
    LocalMux I__3159 (
            .O(N__15134),
            .I(\this_start_data_delay.this_edge_detector.N_213 ));
    InMux I__3158 (
            .O(N__15131),
            .I(N__15128));
    LocalMux I__3157 (
            .O(N__15128),
            .I(N__15125));
    Odrv12 I__3156 (
            .O(N__15125),
            .I(un1_M_current_address_q_cry_11_c_RNI6NLHZ0));
    InMux I__3155 (
            .O(N__15122),
            .I(un1_M_current_address_q_cry_11));
    InMux I__3154 (
            .O(N__15119),
            .I(un1_M_current_address_q_cry_12));
    CascadeMux I__3153 (
            .O(N__15116),
            .I(N__15112));
    InMux I__3152 (
            .O(N__15115),
            .I(N__15109));
    InMux I__3151 (
            .O(N__15112),
            .I(N__15106));
    LocalMux I__3150 (
            .O(N__15109),
            .I(N_177_0));
    LocalMux I__3149 (
            .O(N__15106),
            .I(N_177_0));
    InMux I__3148 (
            .O(N__15101),
            .I(N__15098));
    LocalMux I__3147 (
            .O(N__15098),
            .I(un1_M_current_address_q_cry_9_c_RNIRDIMZ0));
    InMux I__3146 (
            .O(N__15095),
            .I(N__15092));
    LocalMux I__3145 (
            .O(N__15092),
            .I(N__15089));
    Odrv4 I__3144 (
            .O(N__15089),
            .I(un1_M_current_address_q_cry_0_c_RNI2QANZ0));
    InMux I__3143 (
            .O(N__15086),
            .I(N__15083));
    LocalMux I__3142 (
            .O(N__15083),
            .I(un1_M_current_address_q_cry_12_c_RNI8QMHZ0));
    InMux I__3141 (
            .O(N__15080),
            .I(N__15077));
    LocalMux I__3140 (
            .O(N__15077),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_12 ));
    InMux I__3139 (
            .O(N__15074),
            .I(N__15071));
    LocalMux I__3138 (
            .O(N__15071),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_10 ));
    InMux I__3137 (
            .O(N__15068),
            .I(N__15065));
    LocalMux I__3136 (
            .O(N__15065),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_11 ));
    InMux I__3135 (
            .O(N__15062),
            .I(un1_M_current_address_q_cry_2));
    InMux I__3134 (
            .O(N__15059),
            .I(N__15056));
    LocalMux I__3133 (
            .O(N__15056),
            .I(un1_M_current_address_q_cry_3_c_RNI83ENZ0));
    InMux I__3132 (
            .O(N__15053),
            .I(un1_M_current_address_q_cry_3));
    CascadeMux I__3131 (
            .O(N__15050),
            .I(N__15047));
    CascadeBuf I__3130 (
            .O(N__15047),
            .I(N__15044));
    CascadeMux I__3129 (
            .O(N__15044),
            .I(N__15041));
    CascadeBuf I__3128 (
            .O(N__15041),
            .I(N__15038));
    CascadeMux I__3127 (
            .O(N__15038),
            .I(N__15035));
    CascadeBuf I__3126 (
            .O(N__15035),
            .I(N__15032));
    CascadeMux I__3125 (
            .O(N__15032),
            .I(N__15029));
    CascadeBuf I__3124 (
            .O(N__15029),
            .I(N__15026));
    CascadeMux I__3123 (
            .O(N__15026),
            .I(N__15023));
    CascadeBuf I__3122 (
            .O(N__15023),
            .I(N__15020));
    CascadeMux I__3121 (
            .O(N__15020),
            .I(N__15017));
    CascadeBuf I__3120 (
            .O(N__15017),
            .I(N__15014));
    CascadeMux I__3119 (
            .O(N__15014),
            .I(N__15011));
    CascadeBuf I__3118 (
            .O(N__15011),
            .I(N__15008));
    CascadeMux I__3117 (
            .O(N__15008),
            .I(N__15005));
    CascadeBuf I__3116 (
            .O(N__15005),
            .I(N__15002));
    CascadeMux I__3115 (
            .O(N__15002),
            .I(N__14999));
    CascadeBuf I__3114 (
            .O(N__14999),
            .I(N__14996));
    CascadeMux I__3113 (
            .O(N__14996),
            .I(N__14993));
    CascadeBuf I__3112 (
            .O(N__14993),
            .I(N__14990));
    CascadeMux I__3111 (
            .O(N__14990),
            .I(N__14987));
    CascadeBuf I__3110 (
            .O(N__14987),
            .I(N__14984));
    CascadeMux I__3109 (
            .O(N__14984),
            .I(N__14981));
    CascadeBuf I__3108 (
            .O(N__14981),
            .I(N__14978));
    CascadeMux I__3107 (
            .O(N__14978),
            .I(N__14975));
    CascadeBuf I__3106 (
            .O(N__14975),
            .I(N__14972));
    CascadeMux I__3105 (
            .O(N__14972),
            .I(N__14969));
    CascadeBuf I__3104 (
            .O(N__14969),
            .I(N__14966));
    CascadeMux I__3103 (
            .O(N__14966),
            .I(N__14963));
    CascadeBuf I__3102 (
            .O(N__14963),
            .I(N__14960));
    CascadeMux I__3101 (
            .O(N__14960),
            .I(N__14957));
    InMux I__3100 (
            .O(N__14957),
            .I(N__14954));
    LocalMux I__3099 (
            .O(N__14954),
            .I(N__14951));
    Span4Mux_s3_v I__3098 (
            .O(N__14951),
            .I(N__14946));
    InMux I__3097 (
            .O(N__14950),
            .I(N__14943));
    InMux I__3096 (
            .O(N__14949),
            .I(N__14940));
    Sp12to4 I__3095 (
            .O(N__14946),
            .I(N__14937));
    LocalMux I__3094 (
            .O(N__14943),
            .I(N__14934));
    LocalMux I__3093 (
            .O(N__14940),
            .I(N__14929));
    Span12Mux_h I__3092 (
            .O(N__14937),
            .I(N__14929));
    Odrv4 I__3091 (
            .O(N__14934),
            .I(M_current_address_qZ0Z_5));
    Odrv12 I__3090 (
            .O(N__14929),
            .I(M_current_address_qZ0Z_5));
    InMux I__3089 (
            .O(N__14924),
            .I(N__14921));
    LocalMux I__3088 (
            .O(N__14921),
            .I(un1_M_current_address_q_cry_4_c_RNIA6FNZ0));
    InMux I__3087 (
            .O(N__14918),
            .I(un1_M_current_address_q_cry_4));
    InMux I__3086 (
            .O(N__14915),
            .I(un1_M_current_address_q_cry_5));
    InMux I__3085 (
            .O(N__14912),
            .I(un1_M_current_address_q_cry_6));
    InMux I__3084 (
            .O(N__14909),
            .I(N__14906));
    LocalMux I__3083 (
            .O(N__14906),
            .I(un1_M_current_address_q_cry_7_c_RNIGFINZ0));
    InMux I__3082 (
            .O(N__14903),
            .I(bfn_19_24_0_));
    CascadeMux I__3081 (
            .O(N__14900),
            .I(N__14897));
    CascadeBuf I__3080 (
            .O(N__14897),
            .I(N__14894));
    CascadeMux I__3079 (
            .O(N__14894),
            .I(N__14891));
    CascadeBuf I__3078 (
            .O(N__14891),
            .I(N__14888));
    CascadeMux I__3077 (
            .O(N__14888),
            .I(N__14885));
    CascadeBuf I__3076 (
            .O(N__14885),
            .I(N__14882));
    CascadeMux I__3075 (
            .O(N__14882),
            .I(N__14879));
    CascadeBuf I__3074 (
            .O(N__14879),
            .I(N__14876));
    CascadeMux I__3073 (
            .O(N__14876),
            .I(N__14873));
    CascadeBuf I__3072 (
            .O(N__14873),
            .I(N__14870));
    CascadeMux I__3071 (
            .O(N__14870),
            .I(N__14867));
    CascadeBuf I__3070 (
            .O(N__14867),
            .I(N__14864));
    CascadeMux I__3069 (
            .O(N__14864),
            .I(N__14861));
    CascadeBuf I__3068 (
            .O(N__14861),
            .I(N__14858));
    CascadeMux I__3067 (
            .O(N__14858),
            .I(N__14855));
    CascadeBuf I__3066 (
            .O(N__14855),
            .I(N__14852));
    CascadeMux I__3065 (
            .O(N__14852),
            .I(N__14849));
    CascadeBuf I__3064 (
            .O(N__14849),
            .I(N__14846));
    CascadeMux I__3063 (
            .O(N__14846),
            .I(N__14843));
    CascadeBuf I__3062 (
            .O(N__14843),
            .I(N__14840));
    CascadeMux I__3061 (
            .O(N__14840),
            .I(N__14837));
    CascadeBuf I__3060 (
            .O(N__14837),
            .I(N__14834));
    CascadeMux I__3059 (
            .O(N__14834),
            .I(N__14831));
    CascadeBuf I__3058 (
            .O(N__14831),
            .I(N__14828));
    CascadeMux I__3057 (
            .O(N__14828),
            .I(N__14825));
    CascadeBuf I__3056 (
            .O(N__14825),
            .I(N__14822));
    CascadeMux I__3055 (
            .O(N__14822),
            .I(N__14819));
    CascadeBuf I__3054 (
            .O(N__14819),
            .I(N__14816));
    CascadeMux I__3053 (
            .O(N__14816),
            .I(N__14813));
    CascadeBuf I__3052 (
            .O(N__14813),
            .I(N__14810));
    CascadeMux I__3051 (
            .O(N__14810),
            .I(N__14807));
    InMux I__3050 (
            .O(N__14807),
            .I(N__14804));
    LocalMux I__3049 (
            .O(N__14804),
            .I(N__14801));
    Span4Mux_v I__3048 (
            .O(N__14801),
            .I(N__14796));
    InMux I__3047 (
            .O(N__14800),
            .I(N__14793));
    InMux I__3046 (
            .O(N__14799),
            .I(N__14790));
    Span4Mux_h I__3045 (
            .O(N__14796),
            .I(N__14787));
    LocalMux I__3044 (
            .O(N__14793),
            .I(N__14784));
    LocalMux I__3043 (
            .O(N__14790),
            .I(N__14779));
    Span4Mux_v I__3042 (
            .O(N__14787),
            .I(N__14779));
    Odrv4 I__3041 (
            .O(N__14784),
            .I(M_current_address_qZ0Z_9));
    Odrv4 I__3040 (
            .O(N__14779),
            .I(M_current_address_qZ0Z_9));
    InMux I__3039 (
            .O(N__14774),
            .I(N__14771));
    LocalMux I__3038 (
            .O(N__14771),
            .I(un1_M_current_address_q_cry_8_c_RNIIIJNZ0));
    InMux I__3037 (
            .O(N__14768),
            .I(un1_M_current_address_q_cry_8));
    InMux I__3036 (
            .O(N__14765),
            .I(un1_M_current_address_q_cry_9));
    InMux I__3035 (
            .O(N__14762),
            .I(un1_M_current_address_q_cry_10));
    InMux I__3034 (
            .O(N__14759),
            .I(N__14756));
    LocalMux I__3033 (
            .O(N__14756),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_8 ));
    CascadeMux I__3032 (
            .O(N__14753),
            .I(N__14749));
    CascadeMux I__3031 (
            .O(N__14752),
            .I(N__14746));
    InMux I__3030 (
            .O(N__14749),
            .I(N__14743));
    InMux I__3029 (
            .O(N__14746),
            .I(N__14740));
    LocalMux I__3028 (
            .O(N__14743),
            .I(N__14735));
    LocalMux I__3027 (
            .O(N__14740),
            .I(N__14735));
    Span4Mux_v I__3026 (
            .O(N__14735),
            .I(N__14732));
    Sp12to4 I__3025 (
            .O(N__14732),
            .I(N__14729));
    Span12Mux_h I__3024 (
            .O(N__14729),
            .I(N__14726));
    Odrv12 I__3023 (
            .O(N__14726),
            .I(port_data_c_5));
    CascadeMux I__3022 (
            .O(N__14723),
            .I(N__14720));
    InMux I__3021 (
            .O(N__14720),
            .I(N__14717));
    LocalMux I__3020 (
            .O(N__14717),
            .I(\this_start_data_delay.this_edge_detector.N_222 ));
    InMux I__3019 (
            .O(N__14714),
            .I(N__14711));
    LocalMux I__3018 (
            .O(N__14711),
            .I(N__14708));
    Span4Mux_h I__3017 (
            .O(N__14708),
            .I(N__14705));
    Odrv4 I__3016 (
            .O(N__14705),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_6 ));
    InMux I__3015 (
            .O(N__14702),
            .I(N__14699));
    LocalMux I__3014 (
            .O(N__14699),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_7 ));
    InMux I__3013 (
            .O(N__14696),
            .I(N__14693));
    LocalMux I__3012 (
            .O(N__14693),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_9 ));
    InMux I__3011 (
            .O(N__14690),
            .I(un1_M_current_address_q_cry_0));
    CascadeMux I__3010 (
            .O(N__14687),
            .I(N__14684));
    CascadeBuf I__3009 (
            .O(N__14684),
            .I(N__14681));
    CascadeMux I__3008 (
            .O(N__14681),
            .I(N__14678));
    CascadeBuf I__3007 (
            .O(N__14678),
            .I(N__14675));
    CascadeMux I__3006 (
            .O(N__14675),
            .I(N__14672));
    CascadeBuf I__3005 (
            .O(N__14672),
            .I(N__14669));
    CascadeMux I__3004 (
            .O(N__14669),
            .I(N__14666));
    CascadeBuf I__3003 (
            .O(N__14666),
            .I(N__14663));
    CascadeMux I__3002 (
            .O(N__14663),
            .I(N__14660));
    CascadeBuf I__3001 (
            .O(N__14660),
            .I(N__14657));
    CascadeMux I__3000 (
            .O(N__14657),
            .I(N__14654));
    CascadeBuf I__2999 (
            .O(N__14654),
            .I(N__14651));
    CascadeMux I__2998 (
            .O(N__14651),
            .I(N__14648));
    CascadeBuf I__2997 (
            .O(N__14648),
            .I(N__14645));
    CascadeMux I__2996 (
            .O(N__14645),
            .I(N__14642));
    CascadeBuf I__2995 (
            .O(N__14642),
            .I(N__14639));
    CascadeMux I__2994 (
            .O(N__14639),
            .I(N__14636));
    CascadeBuf I__2993 (
            .O(N__14636),
            .I(N__14633));
    CascadeMux I__2992 (
            .O(N__14633),
            .I(N__14630));
    CascadeBuf I__2991 (
            .O(N__14630),
            .I(N__14627));
    CascadeMux I__2990 (
            .O(N__14627),
            .I(N__14624));
    CascadeBuf I__2989 (
            .O(N__14624),
            .I(N__14621));
    CascadeMux I__2988 (
            .O(N__14621),
            .I(N__14618));
    CascadeBuf I__2987 (
            .O(N__14618),
            .I(N__14615));
    CascadeMux I__2986 (
            .O(N__14615),
            .I(N__14612));
    CascadeBuf I__2985 (
            .O(N__14612),
            .I(N__14609));
    CascadeMux I__2984 (
            .O(N__14609),
            .I(N__14606));
    CascadeBuf I__2983 (
            .O(N__14606),
            .I(N__14603));
    CascadeMux I__2982 (
            .O(N__14603),
            .I(N__14600));
    CascadeBuf I__2981 (
            .O(N__14600),
            .I(N__14597));
    CascadeMux I__2980 (
            .O(N__14597),
            .I(N__14594));
    InMux I__2979 (
            .O(N__14594),
            .I(N__14590));
    InMux I__2978 (
            .O(N__14593),
            .I(N__14586));
    LocalMux I__2977 (
            .O(N__14590),
            .I(N__14583));
    InMux I__2976 (
            .O(N__14589),
            .I(N__14580));
    LocalMux I__2975 (
            .O(N__14586),
            .I(N__14577));
    Span12Mux_s9_v I__2974 (
            .O(N__14583),
            .I(N__14574));
    LocalMux I__2973 (
            .O(N__14580),
            .I(M_current_address_qZ0Z_2));
    Odrv4 I__2972 (
            .O(N__14577),
            .I(M_current_address_qZ0Z_2));
    Odrv12 I__2971 (
            .O(N__14574),
            .I(M_current_address_qZ0Z_2));
    InMux I__2970 (
            .O(N__14567),
            .I(N__14564));
    LocalMux I__2969 (
            .O(N__14564),
            .I(un1_M_current_address_q_cry_1_c_RNI4TBNZ0));
    InMux I__2968 (
            .O(N__14561),
            .I(un1_M_current_address_q_cry_1));
    InMux I__2967 (
            .O(N__14558),
            .I(N__14555));
    LocalMux I__2966 (
            .O(N__14555),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_17 ));
    InMux I__2965 (
            .O(N__14552),
            .I(N__14549));
    LocalMux I__2964 (
            .O(N__14549),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_18 ));
    InMux I__2963 (
            .O(N__14546),
            .I(N__14543));
    LocalMux I__2962 (
            .O(N__14543),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_7 ));
    InMux I__2961 (
            .O(N__14540),
            .I(N__14537));
    LocalMux I__2960 (
            .O(N__14537),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_8 ));
    CascadeMux I__2959 (
            .O(N__14534),
            .I(N__14531));
    InMux I__2958 (
            .O(N__14531),
            .I(N__14528));
    LocalMux I__2957 (
            .O(N__14528),
            .I(N__14525));
    Odrv4 I__2956 (
            .O(N__14525),
            .I(\this_start_data_delay.this_edge_detector.N_215 ));
    CascadeMux I__2955 (
            .O(N__14522),
            .I(N__14519));
    InMux I__2954 (
            .O(N__14519),
            .I(N__14516));
    LocalMux I__2953 (
            .O(N__14516),
            .I(N__14513));
    Odrv4 I__2952 (
            .O(N__14513),
            .I(\this_start_data_delay.this_edge_detector.N_212 ));
    CascadeMux I__2951 (
            .O(N__14510),
            .I(N__14507));
    InMux I__2950 (
            .O(N__14507),
            .I(N__14504));
    LocalMux I__2949 (
            .O(N__14504),
            .I(\this_start_data_delay.this_edge_detector.N_219 ));
    CascadeMux I__2948 (
            .O(N__14501),
            .I(N__14497));
    CascadeMux I__2947 (
            .O(N__14500),
            .I(N__14494));
    InMux I__2946 (
            .O(N__14497),
            .I(N__14491));
    InMux I__2945 (
            .O(N__14494),
            .I(N__14488));
    LocalMux I__2944 (
            .O(N__14491),
            .I(N__14485));
    LocalMux I__2943 (
            .O(N__14488),
            .I(N__14482));
    Span4Mux_h I__2942 (
            .O(N__14485),
            .I(N__14479));
    Span4Mux_h I__2941 (
            .O(N__14482),
            .I(N__14476));
    Span4Mux_v I__2940 (
            .O(N__14479),
            .I(N__14473));
    Span4Mux_h I__2939 (
            .O(N__14476),
            .I(N__14470));
    Odrv4 I__2938 (
            .O(N__14473),
            .I(\this_vram.N_17_0 ));
    Odrv4 I__2937 (
            .O(N__14470),
            .I(\this_vram.N_17_0 ));
    InMux I__2936 (
            .O(N__14465),
            .I(N__14462));
    LocalMux I__2935 (
            .O(N__14462),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_11 ));
    InMux I__2934 (
            .O(N__14459),
            .I(N__14456));
    LocalMux I__2933 (
            .O(N__14456),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_12 ));
    IoInMux I__2932 (
            .O(N__14453),
            .I(N__14450));
    LocalMux I__2931 (
            .O(N__14450),
            .I(N__14447));
    Span12Mux_s7_v I__2930 (
            .O(N__14447),
            .I(N__14444));
    Span12Mux_h I__2929 (
            .O(N__14444),
            .I(N__14441));
    Span12Mux_v I__2928 (
            .O(N__14441),
            .I(N__14438));
    Odrv12 I__2927 (
            .O(N__14438),
            .I(debug_d));
    InMux I__2926 (
            .O(N__14435),
            .I(N__14432));
    LocalMux I__2925 (
            .O(N__14432),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_13 ));
    InMux I__2924 (
            .O(N__14429),
            .I(N__14426));
    LocalMux I__2923 (
            .O(N__14426),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_14 ));
    InMux I__2922 (
            .O(N__14423),
            .I(N__14420));
    LocalMux I__2921 (
            .O(N__14420),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_15 ));
    InMux I__2920 (
            .O(N__14417),
            .I(N__14414));
    LocalMux I__2919 (
            .O(N__14414),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_16 ));
    InMux I__2918 (
            .O(N__14411),
            .I(N__14408));
    LocalMux I__2917 (
            .O(N__14408),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_3 ));
    InMux I__2916 (
            .O(N__14405),
            .I(N__14402));
    LocalMux I__2915 (
            .O(N__14402),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_4 ));
    InMux I__2914 (
            .O(N__14399),
            .I(N__14396));
    LocalMux I__2913 (
            .O(N__14396),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_10 ));
    InMux I__2912 (
            .O(N__14393),
            .I(N__14390));
    LocalMux I__2911 (
            .O(N__14390),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_9 ));
    InMux I__2910 (
            .O(N__14387),
            .I(N__14384));
    LocalMux I__2909 (
            .O(N__14384),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_6 ));
    InMux I__2908 (
            .O(N__14381),
            .I(N__14378));
    LocalMux I__2907 (
            .O(N__14378),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_4 ));
    InMux I__2906 (
            .O(N__14375),
            .I(N__14372));
    LocalMux I__2905 (
            .O(N__14372),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_5 ));
    InMux I__2904 (
            .O(N__14369),
            .I(N__14365));
    InMux I__2903 (
            .O(N__14368),
            .I(N__14362));
    LocalMux I__2902 (
            .O(N__14365),
            .I(N__14359));
    LocalMux I__2901 (
            .O(N__14362),
            .I(N__14354));
    Span4Mux_h I__2900 (
            .O(N__14359),
            .I(N__14345));
    InMux I__2899 (
            .O(N__14358),
            .I(N__14342));
    InMux I__2898 (
            .O(N__14357),
            .I(N__14339));
    Span4Mux_h I__2897 (
            .O(N__14354),
            .I(N__14336));
    InMux I__2896 (
            .O(N__14353),
            .I(N__14333));
    InMux I__2895 (
            .O(N__14352),
            .I(N__14330));
    InMux I__2894 (
            .O(N__14351),
            .I(N__14327));
    InMux I__2893 (
            .O(N__14350),
            .I(N__14322));
    InMux I__2892 (
            .O(N__14349),
            .I(N__14322));
    InMux I__2891 (
            .O(N__14348),
            .I(N__14319));
    Odrv4 I__2890 (
            .O(N__14345),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__2889 (
            .O(N__14342),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__2888 (
            .O(N__14339),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    Odrv4 I__2887 (
            .O(N__14336),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__2886 (
            .O(N__14333),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__2885 (
            .O(N__14330),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__2884 (
            .O(N__14327),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__2883 (
            .O(N__14322),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__2882 (
            .O(N__14319),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    InMux I__2881 (
            .O(N__14300),
            .I(N__14296));
    InMux I__2880 (
            .O(N__14299),
            .I(N__14293));
    LocalMux I__2879 (
            .O(N__14296),
            .I(N__14290));
    LocalMux I__2878 (
            .O(N__14293),
            .I(N__14281));
    Span4Mux_h I__2877 (
            .O(N__14290),
            .I(N__14278));
    InMux I__2876 (
            .O(N__14289),
            .I(N__14275));
    InMux I__2875 (
            .O(N__14288),
            .I(N__14268));
    InMux I__2874 (
            .O(N__14287),
            .I(N__14268));
    InMux I__2873 (
            .O(N__14286),
            .I(N__14268));
    InMux I__2872 (
            .O(N__14285),
            .I(N__14263));
    InMux I__2871 (
            .O(N__14284),
            .I(N__14263));
    Odrv12 I__2870 (
            .O(N__14281),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1 ));
    Odrv4 I__2869 (
            .O(N__14278),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1 ));
    LocalMux I__2868 (
            .O(N__14275),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1 ));
    LocalMux I__2867 (
            .O(N__14268),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1 ));
    LocalMux I__2866 (
            .O(N__14263),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1 ));
    CascadeMux I__2865 (
            .O(N__14252),
            .I(N__14249));
    CascadeBuf I__2864 (
            .O(N__14249),
            .I(N__14246));
    CascadeMux I__2863 (
            .O(N__14246),
            .I(N__14243));
    CascadeBuf I__2862 (
            .O(N__14243),
            .I(N__14240));
    CascadeMux I__2861 (
            .O(N__14240),
            .I(N__14237));
    CascadeBuf I__2860 (
            .O(N__14237),
            .I(N__14234));
    CascadeMux I__2859 (
            .O(N__14234),
            .I(N__14231));
    CascadeBuf I__2858 (
            .O(N__14231),
            .I(N__14228));
    CascadeMux I__2857 (
            .O(N__14228),
            .I(N__14225));
    CascadeBuf I__2856 (
            .O(N__14225),
            .I(N__14222));
    CascadeMux I__2855 (
            .O(N__14222),
            .I(N__14219));
    CascadeBuf I__2854 (
            .O(N__14219),
            .I(N__14216));
    CascadeMux I__2853 (
            .O(N__14216),
            .I(N__14213));
    CascadeBuf I__2852 (
            .O(N__14213),
            .I(N__14210));
    CascadeMux I__2851 (
            .O(N__14210),
            .I(N__14207));
    CascadeBuf I__2850 (
            .O(N__14207),
            .I(N__14204));
    CascadeMux I__2849 (
            .O(N__14204),
            .I(N__14201));
    CascadeBuf I__2848 (
            .O(N__14201),
            .I(N__14198));
    CascadeMux I__2847 (
            .O(N__14198),
            .I(N__14195));
    CascadeBuf I__2846 (
            .O(N__14195),
            .I(N__14192));
    CascadeMux I__2845 (
            .O(N__14192),
            .I(N__14189));
    CascadeBuf I__2844 (
            .O(N__14189),
            .I(N__14186));
    CascadeMux I__2843 (
            .O(N__14186),
            .I(N__14183));
    CascadeBuf I__2842 (
            .O(N__14183),
            .I(N__14180));
    CascadeMux I__2841 (
            .O(N__14180),
            .I(N__14177));
    CascadeBuf I__2840 (
            .O(N__14177),
            .I(N__14174));
    CascadeMux I__2839 (
            .O(N__14174),
            .I(N__14171));
    CascadeBuf I__2838 (
            .O(N__14171),
            .I(N__14168));
    CascadeMux I__2837 (
            .O(N__14168),
            .I(N__14165));
    CascadeBuf I__2836 (
            .O(N__14165),
            .I(N__14162));
    CascadeMux I__2835 (
            .O(N__14162),
            .I(N__14159));
    InMux I__2834 (
            .O(N__14159),
            .I(N__14156));
    LocalMux I__2833 (
            .O(N__14156),
            .I(N__14153));
    Span4Mux_v I__2832 (
            .O(N__14153),
            .I(N__14150));
    Span4Mux_h I__2831 (
            .O(N__14150),
            .I(N__14147));
    Span4Mux_v I__2830 (
            .O(N__14147),
            .I(N__14144));
    Odrv4 I__2829 (
            .O(N__14144),
            .I(M_this_vga_signals_address_10));
    InMux I__2828 (
            .O(N__14141),
            .I(N__14138));
    LocalMux I__2827 (
            .O(N__14138),
            .I(N__14135));
    Odrv4 I__2826 (
            .O(N__14135),
            .I(\this_vram.M_this_vram_read_data_0 ));
    InMux I__2825 (
            .O(N__14132),
            .I(N__14126));
    InMux I__2824 (
            .O(N__14131),
            .I(N__14126));
    LocalMux I__2823 (
            .O(N__14126),
            .I(N__14123));
    Span4Mux_v I__2822 (
            .O(N__14123),
            .I(N__14119));
    InMux I__2821 (
            .O(N__14122),
            .I(N__14116));
    Sp12to4 I__2820 (
            .O(N__14119),
            .I(N__14111));
    LocalMux I__2819 (
            .O(N__14116),
            .I(N__14111));
    Span12Mux_h I__2818 (
            .O(N__14111),
            .I(N__14108));
    Odrv12 I__2817 (
            .O(N__14108),
            .I(port_clk_c));
    InMux I__2816 (
            .O(N__14105),
            .I(N__14101));
    InMux I__2815 (
            .O(N__14104),
            .I(N__14098));
    LocalMux I__2814 (
            .O(N__14101),
            .I(this_start_data_delay_this_edge_detector_M_last_q));
    LocalMux I__2813 (
            .O(N__14098),
            .I(this_start_data_delay_this_edge_detector_M_last_q));
    InMux I__2812 (
            .O(N__14093),
            .I(N__14090));
    LocalMux I__2811 (
            .O(N__14090),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_0 ));
    InMux I__2810 (
            .O(N__14087),
            .I(N__14084));
    LocalMux I__2809 (
            .O(N__14084),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_3 ));
    InMux I__2808 (
            .O(N__14081),
            .I(N__14078));
    LocalMux I__2807 (
            .O(N__14078),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_1 ));
    InMux I__2806 (
            .O(N__14075),
            .I(N__14072));
    LocalMux I__2805 (
            .O(N__14072),
            .I(\this_start_data_delay.this_delay.M_pipe_qZ0Z_2 ));
    InMux I__2804 (
            .O(N__14069),
            .I(N__14066));
    LocalMux I__2803 (
            .O(N__14066),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_5 ));
    InMux I__2802 (
            .O(N__14063),
            .I(N__14060));
    LocalMux I__2801 (
            .O(N__14060),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_1 ));
    InMux I__2800 (
            .O(N__14057),
            .I(N__14054));
    LocalMux I__2799 (
            .O(N__14054),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_2 ));
    InMux I__2798 (
            .O(N__14051),
            .I(N__14043));
    InMux I__2797 (
            .O(N__14050),
            .I(N__14043));
    InMux I__2796 (
            .O(N__14049),
            .I(N__14039));
    InMux I__2795 (
            .O(N__14048),
            .I(N__14036));
    LocalMux I__2794 (
            .O(N__14043),
            .I(N__14033));
    InMux I__2793 (
            .O(N__14042),
            .I(N__14030));
    LocalMux I__2792 (
            .O(N__14039),
            .I(N__14025));
    LocalMux I__2791 (
            .O(N__14036),
            .I(N__14025));
    Span4Mux_h I__2790 (
            .O(N__14033),
            .I(N__14022));
    LocalMux I__2789 (
            .O(N__14030),
            .I(N__14017));
    Span12Mux_v I__2788 (
            .O(N__14025),
            .I(N__14017));
    Odrv4 I__2787 (
            .O(N__14022),
            .I(\this_vga_signals.un12_address_cry_2_c_RNIPIBB ));
    Odrv12 I__2786 (
            .O(N__14017),
            .I(\this_vga_signals.un12_address_cry_2_c_RNIPIBB ));
    InMux I__2785 (
            .O(N__14012),
            .I(N__14009));
    LocalMux I__2784 (
            .O(N__14009),
            .I(N__14005));
    InMux I__2783 (
            .O(N__14008),
            .I(N__14002));
    Span12Mux_s10_h I__2782 (
            .O(N__14005),
            .I(N__13997));
    LocalMux I__2781 (
            .O(N__14002),
            .I(N__13997));
    Span12Mux_h I__2780 (
            .O(N__13997),
            .I(N__13994));
    Odrv12 I__2779 (
            .O(N__13994),
            .I(\this_vga_signals.un12_address_cry_1_c_RNINFAB ));
    CascadeMux I__2778 (
            .O(N__13991),
            .I(\this_vga_signals.mult1_un96_sum_c5_0_1_0_1_cascade_ ));
    InMux I__2777 (
            .O(N__13988),
            .I(N__13985));
    LocalMux I__2776 (
            .O(N__13985),
            .I(\this_vga_signals.N_3_1_2 ));
    InMux I__2775 (
            .O(N__13982),
            .I(N__13979));
    LocalMux I__2774 (
            .O(N__13979),
            .I(\this_vga_signals.g1_0_0_0_1 ));
    CascadeMux I__2773 (
            .O(N__13976),
            .I(\this_vga_signals.mult1_un96_sum_c5_cascade_ ));
    InMux I__2772 (
            .O(N__13973),
            .I(N__13970));
    LocalMux I__2771 (
            .O(N__13970),
            .I(N__13967));
    Odrv4 I__2770 (
            .O(N__13967),
            .I(\this_vga_signals.g2_0 ));
    InMux I__2769 (
            .O(N__13964),
            .I(N__13961));
    LocalMux I__2768 (
            .O(N__13961),
            .I(\this_vga_signals.mult1_un96_sum_axbxc5_2 ));
    CascadeMux I__2767 (
            .O(N__13958),
            .I(\this_vga_signals.g1_0_3_cascade_ ));
    InMux I__2766 (
            .O(N__13955),
            .I(N__13952));
    LocalMux I__2765 (
            .O(N__13952),
            .I(\this_vga_signals.mult1_un89_sum_c5_0_0_0_0 ));
    CascadeMux I__2764 (
            .O(N__13949),
            .I(N__13946));
    CascadeBuf I__2763 (
            .O(N__13946),
            .I(N__13943));
    CascadeMux I__2762 (
            .O(N__13943),
            .I(N__13940));
    CascadeBuf I__2761 (
            .O(N__13940),
            .I(N__13937));
    CascadeMux I__2760 (
            .O(N__13937),
            .I(N__13934));
    CascadeBuf I__2759 (
            .O(N__13934),
            .I(N__13931));
    CascadeMux I__2758 (
            .O(N__13931),
            .I(N__13928));
    CascadeBuf I__2757 (
            .O(N__13928),
            .I(N__13925));
    CascadeMux I__2756 (
            .O(N__13925),
            .I(N__13922));
    CascadeBuf I__2755 (
            .O(N__13922),
            .I(N__13919));
    CascadeMux I__2754 (
            .O(N__13919),
            .I(N__13916));
    CascadeBuf I__2753 (
            .O(N__13916),
            .I(N__13913));
    CascadeMux I__2752 (
            .O(N__13913),
            .I(N__13910));
    CascadeBuf I__2751 (
            .O(N__13910),
            .I(N__13907));
    CascadeMux I__2750 (
            .O(N__13907),
            .I(N__13904));
    CascadeBuf I__2749 (
            .O(N__13904),
            .I(N__13901));
    CascadeMux I__2748 (
            .O(N__13901),
            .I(N__13898));
    CascadeBuf I__2747 (
            .O(N__13898),
            .I(N__13895));
    CascadeMux I__2746 (
            .O(N__13895),
            .I(N__13892));
    CascadeBuf I__2745 (
            .O(N__13892),
            .I(N__13889));
    CascadeMux I__2744 (
            .O(N__13889),
            .I(N__13886));
    CascadeBuf I__2743 (
            .O(N__13886),
            .I(N__13883));
    CascadeMux I__2742 (
            .O(N__13883),
            .I(N__13880));
    CascadeBuf I__2741 (
            .O(N__13880),
            .I(N__13877));
    CascadeMux I__2740 (
            .O(N__13877),
            .I(N__13874));
    CascadeBuf I__2739 (
            .O(N__13874),
            .I(N__13871));
    CascadeMux I__2738 (
            .O(N__13871),
            .I(N__13868));
    CascadeBuf I__2737 (
            .O(N__13868),
            .I(N__13865));
    CascadeMux I__2736 (
            .O(N__13865),
            .I(N__13862));
    CascadeBuf I__2735 (
            .O(N__13862),
            .I(N__13859));
    CascadeMux I__2734 (
            .O(N__13859),
            .I(N__13856));
    InMux I__2733 (
            .O(N__13856),
            .I(N__13853));
    LocalMux I__2732 (
            .O(N__13853),
            .I(N__13850));
    Span12Mux_h I__2731 (
            .O(N__13850),
            .I(N__13847));
    Span12Mux_v I__2730 (
            .O(N__13847),
            .I(N__13844));
    Odrv12 I__2729 (
            .O(N__13844),
            .I(M_this_vga_signals_address_0));
    InMux I__2728 (
            .O(N__13841),
            .I(N__13838));
    LocalMux I__2727 (
            .O(N__13838),
            .I(N__13835));
    Span4Mux_h I__2726 (
            .O(N__13835),
            .I(N__13832));
    Odrv4 I__2725 (
            .O(N__13832),
            .I(\this_vga_signals.g1_0_0 ));
    InMux I__2724 (
            .O(N__13829),
            .I(N__13826));
    LocalMux I__2723 (
            .O(N__13826),
            .I(\this_vga_signals.if_N_3_2_i_1 ));
    CascadeMux I__2722 (
            .O(N__13823),
            .I(N__13810));
    CascadeMux I__2721 (
            .O(N__13822),
            .I(N__13807));
    CascadeMux I__2720 (
            .O(N__13821),
            .I(N__13803));
    CascadeMux I__2719 (
            .O(N__13820),
            .I(N__13799));
    CascadeMux I__2718 (
            .O(N__13819),
            .I(N__13795));
    CascadeMux I__2717 (
            .O(N__13818),
            .I(N__13792));
    CascadeMux I__2716 (
            .O(N__13817),
            .I(N__13789));
    CascadeMux I__2715 (
            .O(N__13816),
            .I(N__13786));
    InMux I__2714 (
            .O(N__13815),
            .I(N__13781));
    CascadeMux I__2713 (
            .O(N__13814),
            .I(N__13778));
    InMux I__2712 (
            .O(N__13813),
            .I(N__13766));
    InMux I__2711 (
            .O(N__13810),
            .I(N__13763));
    InMux I__2710 (
            .O(N__13807),
            .I(N__13757));
    InMux I__2709 (
            .O(N__13806),
            .I(N__13752));
    InMux I__2708 (
            .O(N__13803),
            .I(N__13752));
    CascadeMux I__2707 (
            .O(N__13802),
            .I(N__13749));
    InMux I__2706 (
            .O(N__13799),
            .I(N__13739));
    InMux I__2705 (
            .O(N__13798),
            .I(N__13739));
    InMux I__2704 (
            .O(N__13795),
            .I(N__13739));
    InMux I__2703 (
            .O(N__13792),
            .I(N__13739));
    InMux I__2702 (
            .O(N__13789),
            .I(N__13734));
    InMux I__2701 (
            .O(N__13786),
            .I(N__13734));
    CascadeMux I__2700 (
            .O(N__13785),
            .I(N__13730));
    CascadeMux I__2699 (
            .O(N__13784),
            .I(N__13726));
    LocalMux I__2698 (
            .O(N__13781),
            .I(N__13723));
    InMux I__2697 (
            .O(N__13778),
            .I(N__13720));
    InMux I__2696 (
            .O(N__13777),
            .I(N__13717));
    InMux I__2695 (
            .O(N__13776),
            .I(N__13710));
    InMux I__2694 (
            .O(N__13775),
            .I(N__13710));
    InMux I__2693 (
            .O(N__13774),
            .I(N__13710));
    InMux I__2692 (
            .O(N__13773),
            .I(N__13706));
    InMux I__2691 (
            .O(N__13772),
            .I(N__13703));
    InMux I__2690 (
            .O(N__13771),
            .I(N__13698));
    InMux I__2689 (
            .O(N__13770),
            .I(N__13698));
    InMux I__2688 (
            .O(N__13769),
            .I(N__13695));
    LocalMux I__2687 (
            .O(N__13766),
            .I(N__13690));
    LocalMux I__2686 (
            .O(N__13763),
            .I(N__13690));
    InMux I__2685 (
            .O(N__13762),
            .I(N__13687));
    InMux I__2684 (
            .O(N__13761),
            .I(N__13682));
    InMux I__2683 (
            .O(N__13760),
            .I(N__13682));
    LocalMux I__2682 (
            .O(N__13757),
            .I(N__13677));
    LocalMux I__2681 (
            .O(N__13752),
            .I(N__13677));
    InMux I__2680 (
            .O(N__13749),
            .I(N__13674));
    InMux I__2679 (
            .O(N__13748),
            .I(N__13671));
    LocalMux I__2678 (
            .O(N__13739),
            .I(N__13666));
    LocalMux I__2677 (
            .O(N__13734),
            .I(N__13666));
    InMux I__2676 (
            .O(N__13733),
            .I(N__13657));
    InMux I__2675 (
            .O(N__13730),
            .I(N__13657));
    InMux I__2674 (
            .O(N__13729),
            .I(N__13657));
    InMux I__2673 (
            .O(N__13726),
            .I(N__13657));
    Span4Mux_v I__2672 (
            .O(N__13723),
            .I(N__13654));
    LocalMux I__2671 (
            .O(N__13720),
            .I(N__13649));
    LocalMux I__2670 (
            .O(N__13717),
            .I(N__13649));
    LocalMux I__2669 (
            .O(N__13710),
            .I(N__13646));
    InMux I__2668 (
            .O(N__13709),
            .I(N__13643));
    LocalMux I__2667 (
            .O(N__13706),
            .I(N__13640));
    LocalMux I__2666 (
            .O(N__13703),
            .I(N__13633));
    LocalMux I__2665 (
            .O(N__13698),
            .I(N__13633));
    LocalMux I__2664 (
            .O(N__13695),
            .I(N__13633));
    Span4Mux_v I__2663 (
            .O(N__13690),
            .I(N__13630));
    LocalMux I__2662 (
            .O(N__13687),
            .I(N__13625));
    LocalMux I__2661 (
            .O(N__13682),
            .I(N__13625));
    Span4Mux_h I__2660 (
            .O(N__13677),
            .I(N__13614));
    LocalMux I__2659 (
            .O(N__13674),
            .I(N__13614));
    LocalMux I__2658 (
            .O(N__13671),
            .I(N__13614));
    Span4Mux_v I__2657 (
            .O(N__13666),
            .I(N__13614));
    LocalMux I__2656 (
            .O(N__13657),
            .I(N__13614));
    Span4Mux_h I__2655 (
            .O(N__13654),
            .I(N__13611));
    Span4Mux_h I__2654 (
            .O(N__13649),
            .I(N__13604));
    Span4Mux_v I__2653 (
            .O(N__13646),
            .I(N__13604));
    LocalMux I__2652 (
            .O(N__13643),
            .I(N__13604));
    Span4Mux_h I__2651 (
            .O(N__13640),
            .I(N__13599));
    Span4Mux_h I__2650 (
            .O(N__13633),
            .I(N__13599));
    Span4Mux_h I__2649 (
            .O(N__13630),
            .I(N__13592));
    Span4Mux_h I__2648 (
            .O(N__13625),
            .I(N__13592));
    Span4Mux_h I__2647 (
            .O(N__13614),
            .I(N__13592));
    Odrv4 I__2646 (
            .O(N__13611),
            .I(\this_vga_signals.un12_address_cry_4_c_RNITODB ));
    Odrv4 I__2645 (
            .O(N__13604),
            .I(\this_vga_signals.un12_address_cry_4_c_RNITODB ));
    Odrv4 I__2644 (
            .O(N__13599),
            .I(\this_vga_signals.un12_address_cry_4_c_RNITODB ));
    Odrv4 I__2643 (
            .O(N__13592),
            .I(\this_vga_signals.un12_address_cry_4_c_RNITODB ));
    InMux I__2642 (
            .O(N__13583),
            .I(N__13580));
    LocalMux I__2641 (
            .O(N__13580),
            .I(N__13571));
    InMux I__2640 (
            .O(N__13579),
            .I(N__13566));
    InMux I__2639 (
            .O(N__13578),
            .I(N__13566));
    CascadeMux I__2638 (
            .O(N__13577),
            .I(N__13560));
    CascadeMux I__2637 (
            .O(N__13576),
            .I(N__13557));
    InMux I__2636 (
            .O(N__13575),
            .I(N__13549));
    InMux I__2635 (
            .O(N__13574),
            .I(N__13546));
    Span4Mux_v I__2634 (
            .O(N__13571),
            .I(N__13541));
    LocalMux I__2633 (
            .O(N__13566),
            .I(N__13541));
    InMux I__2632 (
            .O(N__13565),
            .I(N__13532));
    InMux I__2631 (
            .O(N__13564),
            .I(N__13532));
    InMux I__2630 (
            .O(N__13563),
            .I(N__13532));
    InMux I__2629 (
            .O(N__13560),
            .I(N__13532));
    InMux I__2628 (
            .O(N__13557),
            .I(N__13529));
    InMux I__2627 (
            .O(N__13556),
            .I(N__13524));
    InMux I__2626 (
            .O(N__13555),
            .I(N__13524));
    InMux I__2625 (
            .O(N__13554),
            .I(N__13519));
    InMux I__2624 (
            .O(N__13553),
            .I(N__13519));
    InMux I__2623 (
            .O(N__13552),
            .I(N__13516));
    LocalMux I__2622 (
            .O(N__13549),
            .I(N__13513));
    LocalMux I__2621 (
            .O(N__13546),
            .I(\this_vga_signals.mult1_un75_sum_axbxc5 ));
    Odrv4 I__2620 (
            .O(N__13541),
            .I(\this_vga_signals.mult1_un75_sum_axbxc5 ));
    LocalMux I__2619 (
            .O(N__13532),
            .I(\this_vga_signals.mult1_un75_sum_axbxc5 ));
    LocalMux I__2618 (
            .O(N__13529),
            .I(\this_vga_signals.mult1_un75_sum_axbxc5 ));
    LocalMux I__2617 (
            .O(N__13524),
            .I(\this_vga_signals.mult1_un75_sum_axbxc5 ));
    LocalMux I__2616 (
            .O(N__13519),
            .I(\this_vga_signals.mult1_un75_sum_axbxc5 ));
    LocalMux I__2615 (
            .O(N__13516),
            .I(\this_vga_signals.mult1_un75_sum_axbxc5 ));
    Odrv4 I__2614 (
            .O(N__13513),
            .I(\this_vga_signals.mult1_un75_sum_axbxc5 ));
    InMux I__2613 (
            .O(N__13496),
            .I(N__13493));
    LocalMux I__2612 (
            .O(N__13493),
            .I(\this_vga_signals.mult1_un82_sum_ac0_7_0_1_3 ));
    CascadeMux I__2611 (
            .O(N__13490),
            .I(N__13483));
    CascadeMux I__2610 (
            .O(N__13489),
            .I(N__13479));
    CascadeMux I__2609 (
            .O(N__13488),
            .I(N__13475));
    InMux I__2608 (
            .O(N__13487),
            .I(N__13472));
    InMux I__2607 (
            .O(N__13486),
            .I(N__13467));
    InMux I__2606 (
            .O(N__13483),
            .I(N__13458));
    InMux I__2605 (
            .O(N__13482),
            .I(N__13458));
    InMux I__2604 (
            .O(N__13479),
            .I(N__13455));
    InMux I__2603 (
            .O(N__13478),
            .I(N__13444));
    InMux I__2602 (
            .O(N__13475),
            .I(N__13441));
    LocalMux I__2601 (
            .O(N__13472),
            .I(N__13438));
    InMux I__2600 (
            .O(N__13471),
            .I(N__13433));
    InMux I__2599 (
            .O(N__13470),
            .I(N__13433));
    LocalMux I__2598 (
            .O(N__13467),
            .I(N__13430));
    InMux I__2597 (
            .O(N__13466),
            .I(N__13425));
    InMux I__2596 (
            .O(N__13465),
            .I(N__13425));
    InMux I__2595 (
            .O(N__13464),
            .I(N__13422));
    InMux I__2594 (
            .O(N__13463),
            .I(N__13419));
    LocalMux I__2593 (
            .O(N__13458),
            .I(N__13414));
    LocalMux I__2592 (
            .O(N__13455),
            .I(N__13414));
    InMux I__2591 (
            .O(N__13454),
            .I(N__13409));
    InMux I__2590 (
            .O(N__13453),
            .I(N__13409));
    CascadeMux I__2589 (
            .O(N__13452),
            .I(N__13406));
    CascadeMux I__2588 (
            .O(N__13451),
            .I(N__13403));
    InMux I__2587 (
            .O(N__13450),
            .I(N__13396));
    InMux I__2586 (
            .O(N__13449),
            .I(N__13393));
    InMux I__2585 (
            .O(N__13448),
            .I(N__13390));
    InMux I__2584 (
            .O(N__13447),
            .I(N__13387));
    LocalMux I__2583 (
            .O(N__13444),
            .I(N__13378));
    LocalMux I__2582 (
            .O(N__13441),
            .I(N__13378));
    Span4Mux_v I__2581 (
            .O(N__13438),
            .I(N__13378));
    LocalMux I__2580 (
            .O(N__13433),
            .I(N__13378));
    Span4Mux_v I__2579 (
            .O(N__13430),
            .I(N__13373));
    LocalMux I__2578 (
            .O(N__13425),
            .I(N__13373));
    LocalMux I__2577 (
            .O(N__13422),
            .I(N__13368));
    LocalMux I__2576 (
            .O(N__13419),
            .I(N__13368));
    Span4Mux_v I__2575 (
            .O(N__13414),
            .I(N__13363));
    LocalMux I__2574 (
            .O(N__13409),
            .I(N__13363));
    InMux I__2573 (
            .O(N__13406),
            .I(N__13360));
    InMux I__2572 (
            .O(N__13403),
            .I(N__13355));
    InMux I__2571 (
            .O(N__13402),
            .I(N__13355));
    InMux I__2570 (
            .O(N__13401),
            .I(N__13350));
    InMux I__2569 (
            .O(N__13400),
            .I(N__13350));
    InMux I__2568 (
            .O(N__13399),
            .I(N__13346));
    LocalMux I__2567 (
            .O(N__13396),
            .I(N__13337));
    LocalMux I__2566 (
            .O(N__13393),
            .I(N__13337));
    LocalMux I__2565 (
            .O(N__13390),
            .I(N__13337));
    LocalMux I__2564 (
            .O(N__13387),
            .I(N__13337));
    Span4Mux_h I__2563 (
            .O(N__13378),
            .I(N__13334));
    Span4Mux_h I__2562 (
            .O(N__13373),
            .I(N__13329));
    Span4Mux_h I__2561 (
            .O(N__13368),
            .I(N__13329));
    Span4Mux_h I__2560 (
            .O(N__13363),
            .I(N__13324));
    LocalMux I__2559 (
            .O(N__13360),
            .I(N__13324));
    LocalMux I__2558 (
            .O(N__13355),
            .I(N__13319));
    LocalMux I__2557 (
            .O(N__13350),
            .I(N__13319));
    InMux I__2556 (
            .O(N__13349),
            .I(N__13316));
    LocalMux I__2555 (
            .O(N__13346),
            .I(\this_vga_signals.un12_address_cry_5_c_RNIVREB ));
    Odrv12 I__2554 (
            .O(N__13337),
            .I(\this_vga_signals.un12_address_cry_5_c_RNIVREB ));
    Odrv4 I__2553 (
            .O(N__13334),
            .I(\this_vga_signals.un12_address_cry_5_c_RNIVREB ));
    Odrv4 I__2552 (
            .O(N__13329),
            .I(\this_vga_signals.un12_address_cry_5_c_RNIVREB ));
    Odrv4 I__2551 (
            .O(N__13324),
            .I(\this_vga_signals.un12_address_cry_5_c_RNIVREB ));
    Odrv4 I__2550 (
            .O(N__13319),
            .I(\this_vga_signals.un12_address_cry_5_c_RNIVREB ));
    LocalMux I__2549 (
            .O(N__13316),
            .I(\this_vga_signals.un12_address_cry_5_c_RNIVREB ));
    InMux I__2548 (
            .O(N__13301),
            .I(N__13295));
    InMux I__2547 (
            .O(N__13300),
            .I(N__13292));
    InMux I__2546 (
            .O(N__13299),
            .I(N__13289));
    InMux I__2545 (
            .O(N__13298),
            .I(N__13284));
    LocalMux I__2544 (
            .O(N__13295),
            .I(N__13275));
    LocalMux I__2543 (
            .O(N__13292),
            .I(N__13272));
    LocalMux I__2542 (
            .O(N__13289),
            .I(N__13268));
    InMux I__2541 (
            .O(N__13288),
            .I(N__13265));
    InMux I__2540 (
            .O(N__13287),
            .I(N__13262));
    LocalMux I__2539 (
            .O(N__13284),
            .I(N__13259));
    InMux I__2538 (
            .O(N__13283),
            .I(N__13256));
    InMux I__2537 (
            .O(N__13282),
            .I(N__13253));
    InMux I__2536 (
            .O(N__13281),
            .I(N__13250));
    InMux I__2535 (
            .O(N__13280),
            .I(N__13245));
    InMux I__2534 (
            .O(N__13279),
            .I(N__13245));
    InMux I__2533 (
            .O(N__13278),
            .I(N__13242));
    Span4Mux_h I__2532 (
            .O(N__13275),
            .I(N__13237));
    Span4Mux_h I__2531 (
            .O(N__13272),
            .I(N__13237));
    InMux I__2530 (
            .O(N__13271),
            .I(N__13234));
    Odrv12 I__2529 (
            .O(N__13268),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    LocalMux I__2528 (
            .O(N__13265),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    LocalMux I__2527 (
            .O(N__13262),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    Odrv4 I__2526 (
            .O(N__13259),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    LocalMux I__2525 (
            .O(N__13256),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    LocalMux I__2524 (
            .O(N__13253),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    LocalMux I__2523 (
            .O(N__13250),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    LocalMux I__2522 (
            .O(N__13245),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    LocalMux I__2521 (
            .O(N__13242),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    Odrv4 I__2520 (
            .O(N__13237),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    LocalMux I__2519 (
            .O(N__13234),
            .I(this_vga_signals_un17_address_if_m2_2_0));
    CascadeMux I__2518 (
            .O(N__13211),
            .I(N__13207));
    CascadeMux I__2517 (
            .O(N__13210),
            .I(N__13204));
    InMux I__2516 (
            .O(N__13207),
            .I(N__13201));
    InMux I__2515 (
            .O(N__13204),
            .I(N__13198));
    LocalMux I__2514 (
            .O(N__13201),
            .I(N__13193));
    LocalMux I__2513 (
            .O(N__13198),
            .I(N__13193));
    Odrv12 I__2512 (
            .O(N__13193),
            .I(\this_vga_signals.g0_38 ));
    InMux I__2511 (
            .O(N__13190),
            .I(N__13186));
    InMux I__2510 (
            .O(N__13189),
            .I(N__13183));
    LocalMux I__2509 (
            .O(N__13186),
            .I(N__13180));
    LocalMux I__2508 (
            .O(N__13183),
            .I(\this_vga_signals.N_4_0_1 ));
    Odrv4 I__2507 (
            .O(N__13180),
            .I(\this_vga_signals.N_4_0_1 ));
    InMux I__2506 (
            .O(N__13175),
            .I(N__13172));
    LocalMux I__2505 (
            .O(N__13172),
            .I(\this_vga_signals.if_N_3_2_i_2_0 ));
    InMux I__2504 (
            .O(N__13169),
            .I(N__13166));
    LocalMux I__2503 (
            .O(N__13166),
            .I(\this_start_address_delay.this_delay.M_pipe_qZ0Z_0 ));
    InMux I__2502 (
            .O(N__13163),
            .I(N__13160));
    LocalMux I__2501 (
            .O(N__13160),
            .I(\this_vga_signals.g1_0_0_0_0 ));
    CascadeMux I__2500 (
            .O(N__13157),
            .I(\this_vga_signals.g0_0_3_cascade_ ));
    InMux I__2499 (
            .O(N__13154),
            .I(N__13151));
    LocalMux I__2498 (
            .O(N__13151),
            .I(\this_vga_signals.mult1_un82_sum_ac0_7_0_1_4 ));
    InMux I__2497 (
            .O(N__13148),
            .I(N__13145));
    LocalMux I__2496 (
            .O(N__13145),
            .I(\this_vga_signals.g0_6 ));
    InMux I__2495 (
            .O(N__13142),
            .I(N__13139));
    LocalMux I__2494 (
            .O(N__13139),
            .I(\this_vga_signals.g0_13 ));
    InMux I__2493 (
            .O(N__13136),
            .I(N__13132));
    InMux I__2492 (
            .O(N__13135),
            .I(N__13129));
    LocalMux I__2491 (
            .O(N__13132),
            .I(\this_vga_signals.if_N_3_2_i_0 ));
    LocalMux I__2490 (
            .O(N__13129),
            .I(\this_vga_signals.if_N_3_2_i_0 ));
    InMux I__2489 (
            .O(N__13124),
            .I(N__13121));
    LocalMux I__2488 (
            .O(N__13121),
            .I(N__13118));
    Odrv4 I__2487 (
            .O(N__13118),
            .I(\this_vga_signals.g0_0_0_a2_1 ));
    InMux I__2486 (
            .O(N__13115),
            .I(N__13112));
    LocalMux I__2485 (
            .O(N__13112),
            .I(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_0 ));
    CascadeMux I__2484 (
            .O(N__13109),
            .I(\this_vga_signals.g1_2_cascade_ ));
    CascadeMux I__2483 (
            .O(N__13106),
            .I(\this_vga_signals.r_N_2_0_0_2_cascade_ ));
    InMux I__2482 (
            .O(N__13103),
            .I(N__13100));
    LocalMux I__2481 (
            .O(N__13100),
            .I(\this_vga_signals.N_3_1_1 ));
    CascadeMux I__2480 (
            .O(N__13097),
            .I(N__13094));
    InMux I__2479 (
            .O(N__13094),
            .I(N__13091));
    LocalMux I__2478 (
            .O(N__13091),
            .I(N__13088));
    Odrv4 I__2477 (
            .O(N__13088),
            .I(\this_vga_signals.g0_3_1 ));
    InMux I__2476 (
            .O(N__13085),
            .I(N__13078));
    InMux I__2475 (
            .O(N__13084),
            .I(N__13073));
    InMux I__2474 (
            .O(N__13083),
            .I(N__13068));
    InMux I__2473 (
            .O(N__13082),
            .I(N__13063));
    InMux I__2472 (
            .O(N__13081),
            .I(N__13063));
    LocalMux I__2471 (
            .O(N__13078),
            .I(N__13059));
    InMux I__2470 (
            .O(N__13077),
            .I(N__13054));
    InMux I__2469 (
            .O(N__13076),
            .I(N__13054));
    LocalMux I__2468 (
            .O(N__13073),
            .I(N__13051));
    InMux I__2467 (
            .O(N__13072),
            .I(N__13046));
    InMux I__2466 (
            .O(N__13071),
            .I(N__13046));
    LocalMux I__2465 (
            .O(N__13068),
            .I(N__13036));
    LocalMux I__2464 (
            .O(N__13063),
            .I(N__13036));
    InMux I__2463 (
            .O(N__13062),
            .I(N__13032));
    Span4Mux_h I__2462 (
            .O(N__13059),
            .I(N__13027));
    LocalMux I__2461 (
            .O(N__13054),
            .I(N__13027));
    Span4Mux_v I__2460 (
            .O(N__13051),
            .I(N__13022));
    LocalMux I__2459 (
            .O(N__13046),
            .I(N__13022));
    InMux I__2458 (
            .O(N__13045),
            .I(N__13017));
    InMux I__2457 (
            .O(N__13044),
            .I(N__13017));
    InMux I__2456 (
            .O(N__13043),
            .I(N__13010));
    InMux I__2455 (
            .O(N__13042),
            .I(N__13010));
    InMux I__2454 (
            .O(N__13041),
            .I(N__13010));
    Span4Mux_h I__2453 (
            .O(N__13036),
            .I(N__13007));
    InMux I__2452 (
            .O(N__13035),
            .I(N__13004));
    LocalMux I__2451 (
            .O(N__13032),
            .I(\this_vga_signals.mult1_un68_sum_c5 ));
    Odrv4 I__2450 (
            .O(N__13027),
            .I(\this_vga_signals.mult1_un68_sum_c5 ));
    Odrv4 I__2449 (
            .O(N__13022),
            .I(\this_vga_signals.mult1_un68_sum_c5 ));
    LocalMux I__2448 (
            .O(N__13017),
            .I(\this_vga_signals.mult1_un68_sum_c5 ));
    LocalMux I__2447 (
            .O(N__13010),
            .I(\this_vga_signals.mult1_un68_sum_c5 ));
    Odrv4 I__2446 (
            .O(N__13007),
            .I(\this_vga_signals.mult1_un68_sum_c5 ));
    LocalMux I__2445 (
            .O(N__13004),
            .I(\this_vga_signals.mult1_un68_sum_c5 ));
    CascadeMux I__2444 (
            .O(N__12989),
            .I(N__12983));
    CascadeMux I__2443 (
            .O(N__12988),
            .I(N__12972));
    CascadeMux I__2442 (
            .O(N__12987),
            .I(N__12969));
    InMux I__2441 (
            .O(N__12986),
            .I(N__12964));
    InMux I__2440 (
            .O(N__12983),
            .I(N__12964));
    InMux I__2439 (
            .O(N__12982),
            .I(N__12961));
    InMux I__2438 (
            .O(N__12981),
            .I(N__12958));
    InMux I__2437 (
            .O(N__12980),
            .I(N__12954));
    InMux I__2436 (
            .O(N__12979),
            .I(N__12951));
    CascadeMux I__2435 (
            .O(N__12978),
            .I(N__12946));
    InMux I__2434 (
            .O(N__12977),
            .I(N__12942));
    InMux I__2433 (
            .O(N__12976),
            .I(N__12933));
    InMux I__2432 (
            .O(N__12975),
            .I(N__12933));
    InMux I__2431 (
            .O(N__12972),
            .I(N__12933));
    InMux I__2430 (
            .O(N__12969),
            .I(N__12933));
    LocalMux I__2429 (
            .O(N__12964),
            .I(N__12930));
    LocalMux I__2428 (
            .O(N__12961),
            .I(N__12925));
    LocalMux I__2427 (
            .O(N__12958),
            .I(N__12925));
    InMux I__2426 (
            .O(N__12957),
            .I(N__12922));
    LocalMux I__2425 (
            .O(N__12954),
            .I(N__12919));
    LocalMux I__2424 (
            .O(N__12951),
            .I(N__12916));
    InMux I__2423 (
            .O(N__12950),
            .I(N__12913));
    InMux I__2422 (
            .O(N__12949),
            .I(N__12908));
    InMux I__2421 (
            .O(N__12946),
            .I(N__12908));
    CascadeMux I__2420 (
            .O(N__12945),
            .I(N__12904));
    LocalMux I__2419 (
            .O(N__12942),
            .I(N__12901));
    LocalMux I__2418 (
            .O(N__12933),
            .I(N__12898));
    Span4Mux_v I__2417 (
            .O(N__12930),
            .I(N__12891));
    Span4Mux_v I__2416 (
            .O(N__12925),
            .I(N__12891));
    LocalMux I__2415 (
            .O(N__12922),
            .I(N__12891));
    Span4Mux_v I__2414 (
            .O(N__12919),
            .I(N__12888));
    Span4Mux_h I__2413 (
            .O(N__12916),
            .I(N__12881));
    LocalMux I__2412 (
            .O(N__12913),
            .I(N__12881));
    LocalMux I__2411 (
            .O(N__12908),
            .I(N__12881));
    InMux I__2410 (
            .O(N__12907),
            .I(N__12876));
    InMux I__2409 (
            .O(N__12904),
            .I(N__12876));
    Span4Mux_h I__2408 (
            .O(N__12901),
            .I(N__12873));
    Span12Mux_v I__2407 (
            .O(N__12898),
            .I(N__12870));
    Span4Mux_h I__2406 (
            .O(N__12891),
            .I(N__12867));
    Span4Mux_h I__2405 (
            .O(N__12888),
            .I(N__12862));
    Span4Mux_h I__2404 (
            .O(N__12881),
            .I(N__12862));
    LocalMux I__2403 (
            .O(N__12876),
            .I(N__12859));
    Odrv4 I__2402 (
            .O(N__12873),
            .I(\this_vga_signals.un12_address_cry_3_c_RNIRLCB ));
    Odrv12 I__2401 (
            .O(N__12870),
            .I(\this_vga_signals.un12_address_cry_3_c_RNIRLCB ));
    Odrv4 I__2400 (
            .O(N__12867),
            .I(\this_vga_signals.un12_address_cry_3_c_RNIRLCB ));
    Odrv4 I__2399 (
            .O(N__12862),
            .I(\this_vga_signals.un12_address_cry_3_c_RNIRLCB ));
    Odrv4 I__2398 (
            .O(N__12859),
            .I(\this_vga_signals.un12_address_cry_3_c_RNIRLCB ));
    CascadeMux I__2397 (
            .O(N__12848),
            .I(\this_vga_signals.g0_5_3_cascade_ ));
    CascadeMux I__2396 (
            .O(N__12845),
            .I(\this_vga_signals.g0_3_0_a2_1_cascade_ ));
    InMux I__2395 (
            .O(N__12842),
            .I(N__12839));
    LocalMux I__2394 (
            .O(N__12839),
            .I(\this_vga_signals.mult1_un82_sum_ac0_7_0_1_2 ));
    InMux I__2393 (
            .O(N__12836),
            .I(N__12833));
    LocalMux I__2392 (
            .O(N__12833),
            .I(N__12829));
    InMux I__2391 (
            .O(N__12832),
            .I(N__12826));
    Span4Mux_h I__2390 (
            .O(N__12829),
            .I(N__12823));
    LocalMux I__2389 (
            .O(N__12826),
            .I(N__12820));
    Odrv4 I__2388 (
            .O(N__12823),
            .I(\this_vga_signals.if_N_8_mux_2_0 ));
    Odrv4 I__2387 (
            .O(N__12820),
            .I(\this_vga_signals.if_N_8_mux_2_0 ));
    InMux I__2386 (
            .O(N__12815),
            .I(N__12809));
    CascadeMux I__2385 (
            .O(N__12814),
            .I(N__12791));
    CascadeMux I__2384 (
            .O(N__12813),
            .I(N__12787));
    InMux I__2383 (
            .O(N__12812),
            .I(N__12783));
    LocalMux I__2382 (
            .O(N__12809),
            .I(N__12780));
    InMux I__2381 (
            .O(N__12808),
            .I(N__12775));
    InMux I__2380 (
            .O(N__12807),
            .I(N__12775));
    InMux I__2379 (
            .O(N__12806),
            .I(N__12772));
    InMux I__2378 (
            .O(N__12805),
            .I(N__12767));
    InMux I__2377 (
            .O(N__12804),
            .I(N__12767));
    InMux I__2376 (
            .O(N__12803),
            .I(N__12760));
    InMux I__2375 (
            .O(N__12802),
            .I(N__12760));
    InMux I__2374 (
            .O(N__12801),
            .I(N__12760));
    InMux I__2373 (
            .O(N__12800),
            .I(N__12751));
    InMux I__2372 (
            .O(N__12799),
            .I(N__12751));
    InMux I__2371 (
            .O(N__12798),
            .I(N__12751));
    InMux I__2370 (
            .O(N__12797),
            .I(N__12751));
    InMux I__2369 (
            .O(N__12796),
            .I(N__12744));
    InMux I__2368 (
            .O(N__12795),
            .I(N__12744));
    InMux I__2367 (
            .O(N__12794),
            .I(N__12744));
    InMux I__2366 (
            .O(N__12791),
            .I(N__12741));
    InMux I__2365 (
            .O(N__12790),
            .I(N__12734));
    InMux I__2364 (
            .O(N__12787),
            .I(N__12734));
    InMux I__2363 (
            .O(N__12786),
            .I(N__12734));
    LocalMux I__2362 (
            .O(N__12783),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5));
    Odrv4 I__2361 (
            .O(N__12780),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5));
    LocalMux I__2360 (
            .O(N__12775),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5));
    LocalMux I__2359 (
            .O(N__12772),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5));
    LocalMux I__2358 (
            .O(N__12767),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5));
    LocalMux I__2357 (
            .O(N__12760),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5));
    LocalMux I__2356 (
            .O(N__12751),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5));
    LocalMux I__2355 (
            .O(N__12744),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5));
    LocalMux I__2354 (
            .O(N__12741),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5));
    LocalMux I__2353 (
            .O(N__12734),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5));
    InMux I__2352 (
            .O(N__12713),
            .I(N__12707));
    InMux I__2351 (
            .O(N__12712),
            .I(N__12704));
    InMux I__2350 (
            .O(N__12711),
            .I(N__12701));
    InMux I__2349 (
            .O(N__12710),
            .I(N__12698));
    LocalMux I__2348 (
            .O(N__12707),
            .I(\this_vga_signals.if_N_3_2_i ));
    LocalMux I__2347 (
            .O(N__12704),
            .I(\this_vga_signals.if_N_3_2_i ));
    LocalMux I__2346 (
            .O(N__12701),
            .I(\this_vga_signals.if_N_3_2_i ));
    LocalMux I__2345 (
            .O(N__12698),
            .I(\this_vga_signals.if_N_3_2_i ));
    InMux I__2344 (
            .O(N__12689),
            .I(N__12686));
    LocalMux I__2343 (
            .O(N__12686),
            .I(N__12683));
    Span4Mux_h I__2342 (
            .O(N__12683),
            .I(N__12680));
    Odrv4 I__2341 (
            .O(N__12680),
            .I(\this_vga_signals.g1_0_0_0 ));
    CascadeMux I__2340 (
            .O(N__12677),
            .I(N__12668));
    InMux I__2339 (
            .O(N__12676),
            .I(N__12664));
    InMux I__2338 (
            .O(N__12675),
            .I(N__12656));
    CascadeMux I__2337 (
            .O(N__12674),
            .I(N__12653));
    InMux I__2336 (
            .O(N__12673),
            .I(N__12643));
    InMux I__2335 (
            .O(N__12672),
            .I(N__12643));
    InMux I__2334 (
            .O(N__12671),
            .I(N__12643));
    InMux I__2333 (
            .O(N__12668),
            .I(N__12638));
    InMux I__2332 (
            .O(N__12667),
            .I(N__12638));
    LocalMux I__2331 (
            .O(N__12664),
            .I(N__12634));
    InMux I__2330 (
            .O(N__12663),
            .I(N__12629));
    InMux I__2329 (
            .O(N__12662),
            .I(N__12629));
    CascadeMux I__2328 (
            .O(N__12661),
            .I(N__12621));
    InMux I__2327 (
            .O(N__12660),
            .I(N__12615));
    InMux I__2326 (
            .O(N__12659),
            .I(N__12615));
    LocalMux I__2325 (
            .O(N__12656),
            .I(N__12612));
    InMux I__2324 (
            .O(N__12653),
            .I(N__12607));
    InMux I__2323 (
            .O(N__12652),
            .I(N__12607));
    InMux I__2322 (
            .O(N__12651),
            .I(N__12604));
    CascadeMux I__2321 (
            .O(N__12650),
            .I(N__12596));
    LocalMux I__2320 (
            .O(N__12643),
            .I(N__12593));
    LocalMux I__2319 (
            .O(N__12638),
            .I(N__12590));
    InMux I__2318 (
            .O(N__12637),
            .I(N__12586));
    Span4Mux_v I__2317 (
            .O(N__12634),
            .I(N__12581));
    LocalMux I__2316 (
            .O(N__12629),
            .I(N__12581));
    InMux I__2315 (
            .O(N__12628),
            .I(N__12578));
    InMux I__2314 (
            .O(N__12627),
            .I(N__12569));
    InMux I__2313 (
            .O(N__12626),
            .I(N__12569));
    InMux I__2312 (
            .O(N__12625),
            .I(N__12569));
    InMux I__2311 (
            .O(N__12624),
            .I(N__12569));
    InMux I__2310 (
            .O(N__12621),
            .I(N__12564));
    InMux I__2309 (
            .O(N__12620),
            .I(N__12564));
    LocalMux I__2308 (
            .O(N__12615),
            .I(N__12561));
    Span4Mux_h I__2307 (
            .O(N__12612),
            .I(N__12554));
    LocalMux I__2306 (
            .O(N__12607),
            .I(N__12554));
    LocalMux I__2305 (
            .O(N__12604),
            .I(N__12554));
    InMux I__2304 (
            .O(N__12603),
            .I(N__12547));
    InMux I__2303 (
            .O(N__12602),
            .I(N__12547));
    InMux I__2302 (
            .O(N__12601),
            .I(N__12547));
    InMux I__2301 (
            .O(N__12600),
            .I(N__12540));
    InMux I__2300 (
            .O(N__12599),
            .I(N__12540));
    InMux I__2299 (
            .O(N__12596),
            .I(N__12540));
    Span4Mux_h I__2298 (
            .O(N__12593),
            .I(N__12535));
    Span4Mux_h I__2297 (
            .O(N__12590),
            .I(N__12535));
    InMux I__2296 (
            .O(N__12589),
            .I(N__12532));
    LocalMux I__2295 (
            .O(N__12586),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    Odrv4 I__2294 (
            .O(N__12581),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__2293 (
            .O(N__12578),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__2292 (
            .O(N__12569),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__2291 (
            .O(N__12564),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    Odrv4 I__2290 (
            .O(N__12561),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    Odrv4 I__2289 (
            .O(N__12554),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__2288 (
            .O(N__12547),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__2287 (
            .O(N__12540),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    Odrv4 I__2286 (
            .O(N__12535),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__2285 (
            .O(N__12532),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0));
    InMux I__2284 (
            .O(N__12509),
            .I(N__12506));
    LocalMux I__2283 (
            .O(N__12506),
            .I(N__12503));
    Odrv4 I__2282 (
            .O(N__12503),
            .I(\this_vga_signals.g0_6_0 ));
    CascadeMux I__2281 (
            .O(N__12500),
            .I(\this_vga_signals.g1_2_0_cascade_ ));
    InMux I__2280 (
            .O(N__12497),
            .I(N__12494));
    LocalMux I__2279 (
            .O(N__12494),
            .I(N__12491));
    Odrv4 I__2278 (
            .O(N__12491),
            .I(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5 ));
    CascadeMux I__2277 (
            .O(N__12488),
            .I(\this_vga_signals.g1_5_cascade_ ));
    InMux I__2276 (
            .O(N__12485),
            .I(N__12478));
    InMux I__2275 (
            .O(N__12484),
            .I(N__12473));
    InMux I__2274 (
            .O(N__12483),
            .I(N__12473));
    InMux I__2273 (
            .O(N__12482),
            .I(N__12470));
    InMux I__2272 (
            .O(N__12481),
            .I(N__12467));
    LocalMux I__2271 (
            .O(N__12478),
            .I(N__12462));
    LocalMux I__2270 (
            .O(N__12473),
            .I(N__12459));
    LocalMux I__2269 (
            .O(N__12470),
            .I(N__12456));
    LocalMux I__2268 (
            .O(N__12467),
            .I(N__12453));
    InMux I__2267 (
            .O(N__12466),
            .I(N__12448));
    InMux I__2266 (
            .O(N__12465),
            .I(N__12448));
    Span4Mux_v I__2265 (
            .O(N__12462),
            .I(N__12437));
    Span4Mux_v I__2264 (
            .O(N__12459),
            .I(N__12437));
    Span4Mux_h I__2263 (
            .O(N__12456),
            .I(N__12437));
    Span4Mux_v I__2262 (
            .O(N__12453),
            .I(N__12437));
    LocalMux I__2261 (
            .O(N__12448),
            .I(N__12437));
    Odrv4 I__2260 (
            .O(N__12437),
            .I(\this_vga_signals.mult1_un75_sum_axb3 ));
    InMux I__2259 (
            .O(N__12434),
            .I(N__12431));
    LocalMux I__2258 (
            .O(N__12431),
            .I(N__12428));
    Odrv12 I__2257 (
            .O(N__12428),
            .I(\this_vga_signals.g0_0_1_1 ));
    CascadeMux I__2256 (
            .O(N__12425),
            .I(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_2_cascade_ ));
    InMux I__2255 (
            .O(N__12422),
            .I(N__12419));
    LocalMux I__2254 (
            .O(N__12419),
            .I(\this_vga_signals.g0_3 ));
    InMux I__2253 (
            .O(N__12416),
            .I(N__12413));
    LocalMux I__2252 (
            .O(N__12413),
            .I(\this_vga_signals.N_20_i_i_0 ));
    InMux I__2251 (
            .O(N__12410),
            .I(N__12407));
    LocalMux I__2250 (
            .O(N__12407),
            .I(N__12404));
    Odrv4 I__2249 (
            .O(N__12404),
            .I(\this_vga_signals.g0_0_a3_3 ));
    InMux I__2248 (
            .O(N__12401),
            .I(N__12397));
    InMux I__2247 (
            .O(N__12400),
            .I(N__12394));
    LocalMux I__2246 (
            .O(N__12397),
            .I(\this_vga_signals.mult1_un82_sum_ac0_7_0_1_0 ));
    LocalMux I__2245 (
            .O(N__12394),
            .I(\this_vga_signals.mult1_un82_sum_ac0_7_0_1_0 ));
    CascadeMux I__2244 (
            .O(N__12389),
            .I(\this_vga_signals.N_11_cascade_ ));
    InMux I__2243 (
            .O(N__12386),
            .I(N__12383));
    LocalMux I__2242 (
            .O(N__12383),
            .I(\this_vga_signals.g0_0_a3_2 ));
    CascadeMux I__2241 (
            .O(N__12380),
            .I(\this_vga_signals.g0_0_a3_5_cascade_ ));
    InMux I__2240 (
            .O(N__12377),
            .I(N__12374));
    LocalMux I__2239 (
            .O(N__12374),
            .I(\this_vga_signals.g0_i_x4_4_a3 ));
    InMux I__2238 (
            .O(N__12371),
            .I(N__12368));
    LocalMux I__2237 (
            .O(N__12368),
            .I(\this_vga_signals.N_3_3_0 ));
    InMux I__2236 (
            .O(N__12365),
            .I(N__12362));
    LocalMux I__2235 (
            .O(N__12362),
            .I(N__12359));
    Odrv12 I__2234 (
            .O(N__12359),
            .I(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_1 ));
    InMux I__2233 (
            .O(N__12356),
            .I(N__12353));
    LocalMux I__2232 (
            .O(N__12353),
            .I(\this_vga_signals.g0_0_1_0 ));
    CascadeMux I__2231 (
            .O(N__12350),
            .I(\this_vga_signals.g1_5_0_0_cascade_ ));
    InMux I__2230 (
            .O(N__12347),
            .I(N__12344));
    LocalMux I__2229 (
            .O(N__12344),
            .I(\this_vga_signals.r_N_2_0_0_0 ));
    CascadeMux I__2228 (
            .O(N__12341),
            .I(N__12338));
    InMux I__2227 (
            .O(N__12338),
            .I(N__12335));
    LocalMux I__2226 (
            .O(N__12335),
            .I(N__12332));
    Span4Mux_h I__2225 (
            .O(N__12332),
            .I(N__12329));
    Odrv4 I__2224 (
            .O(N__12329),
            .I(\this_vga_signals.g0_1_0 ));
    CascadeMux I__2223 (
            .O(N__12326),
            .I(\this_vga_signals.g0_1_2_cascade_ ));
    InMux I__2222 (
            .O(N__12323),
            .I(N__12320));
    LocalMux I__2221 (
            .O(N__12320),
            .I(N__12310));
    InMux I__2220 (
            .O(N__12319),
            .I(N__12303));
    InMux I__2219 (
            .O(N__12318),
            .I(N__12303));
    InMux I__2218 (
            .O(N__12317),
            .I(N__12295));
    InMux I__2217 (
            .O(N__12316),
            .I(N__12292));
    InMux I__2216 (
            .O(N__12315),
            .I(N__12289));
    InMux I__2215 (
            .O(N__12314),
            .I(N__12284));
    InMux I__2214 (
            .O(N__12313),
            .I(N__12284));
    Span4Mux_h I__2213 (
            .O(N__12310),
            .I(N__12281));
    InMux I__2212 (
            .O(N__12309),
            .I(N__12276));
    InMux I__2211 (
            .O(N__12308),
            .I(N__12276));
    LocalMux I__2210 (
            .O(N__12303),
            .I(N__12273));
    InMux I__2209 (
            .O(N__12302),
            .I(N__12266));
    InMux I__2208 (
            .O(N__12301),
            .I(N__12266));
    InMux I__2207 (
            .O(N__12300),
            .I(N__12266));
    InMux I__2206 (
            .O(N__12299),
            .I(N__12261));
    InMux I__2205 (
            .O(N__12298),
            .I(N__12261));
    LocalMux I__2204 (
            .O(N__12295),
            .I(this_vga_signals_un17_address_if_N_8_mux));
    LocalMux I__2203 (
            .O(N__12292),
            .I(this_vga_signals_un17_address_if_N_8_mux));
    LocalMux I__2202 (
            .O(N__12289),
            .I(this_vga_signals_un17_address_if_N_8_mux));
    LocalMux I__2201 (
            .O(N__12284),
            .I(this_vga_signals_un17_address_if_N_8_mux));
    Odrv4 I__2200 (
            .O(N__12281),
            .I(this_vga_signals_un17_address_if_N_8_mux));
    LocalMux I__2199 (
            .O(N__12276),
            .I(this_vga_signals_un17_address_if_N_8_mux));
    Odrv4 I__2198 (
            .O(N__12273),
            .I(this_vga_signals_un17_address_if_N_8_mux));
    LocalMux I__2197 (
            .O(N__12266),
            .I(this_vga_signals_un17_address_if_N_8_mux));
    LocalMux I__2196 (
            .O(N__12261),
            .I(this_vga_signals_un17_address_if_N_8_mux));
    InMux I__2195 (
            .O(N__12242),
            .I(N__12239));
    LocalMux I__2194 (
            .O(N__12239),
            .I(N__12236));
    Span4Mux_h I__2193 (
            .O(N__12236),
            .I(N__12233));
    Span4Mux_v I__2192 (
            .O(N__12233),
            .I(N__12228));
    InMux I__2191 (
            .O(N__12232),
            .I(N__12223));
    InMux I__2190 (
            .O(N__12231),
            .I(N__12223));
    Odrv4 I__2189 (
            .O(N__12228),
            .I(\this_vga_signals.mult1_un54_sum_ac0_8 ));
    LocalMux I__2188 (
            .O(N__12223),
            .I(\this_vga_signals.mult1_un54_sum_ac0_8 ));
    CascadeMux I__2187 (
            .O(N__12218),
            .I(N__12215));
    CascadeBuf I__2186 (
            .O(N__12215),
            .I(N__12212));
    CascadeMux I__2185 (
            .O(N__12212),
            .I(N__12209));
    CascadeBuf I__2184 (
            .O(N__12209),
            .I(N__12206));
    CascadeMux I__2183 (
            .O(N__12206),
            .I(N__12203));
    CascadeBuf I__2182 (
            .O(N__12203),
            .I(N__12200));
    CascadeMux I__2181 (
            .O(N__12200),
            .I(N__12197));
    CascadeBuf I__2180 (
            .O(N__12197),
            .I(N__12194));
    CascadeMux I__2179 (
            .O(N__12194),
            .I(N__12191));
    CascadeBuf I__2178 (
            .O(N__12191),
            .I(N__12188));
    CascadeMux I__2177 (
            .O(N__12188),
            .I(N__12185));
    CascadeBuf I__2176 (
            .O(N__12185),
            .I(N__12182));
    CascadeMux I__2175 (
            .O(N__12182),
            .I(N__12179));
    CascadeBuf I__2174 (
            .O(N__12179),
            .I(N__12176));
    CascadeMux I__2173 (
            .O(N__12176),
            .I(N__12173));
    CascadeBuf I__2172 (
            .O(N__12173),
            .I(N__12170));
    CascadeMux I__2171 (
            .O(N__12170),
            .I(N__12167));
    CascadeBuf I__2170 (
            .O(N__12167),
            .I(N__12164));
    CascadeMux I__2169 (
            .O(N__12164),
            .I(N__12161));
    CascadeBuf I__2168 (
            .O(N__12161),
            .I(N__12158));
    CascadeMux I__2167 (
            .O(N__12158),
            .I(N__12155));
    CascadeBuf I__2166 (
            .O(N__12155),
            .I(N__12152));
    CascadeMux I__2165 (
            .O(N__12152),
            .I(N__12149));
    CascadeBuf I__2164 (
            .O(N__12149),
            .I(N__12146));
    CascadeMux I__2163 (
            .O(N__12146),
            .I(N__12143));
    CascadeBuf I__2162 (
            .O(N__12143),
            .I(N__12140));
    CascadeMux I__2161 (
            .O(N__12140),
            .I(N__12137));
    CascadeBuf I__2160 (
            .O(N__12137),
            .I(N__12134));
    CascadeMux I__2159 (
            .O(N__12134),
            .I(N__12131));
    CascadeBuf I__2158 (
            .O(N__12131),
            .I(N__12128));
    CascadeMux I__2157 (
            .O(N__12128),
            .I(N__12125));
    InMux I__2156 (
            .O(N__12125),
            .I(N__12122));
    LocalMux I__2155 (
            .O(N__12122),
            .I(N__12119));
    Sp12to4 I__2154 (
            .O(N__12119),
            .I(N__12116));
    Span12Mux_s11_v I__2153 (
            .O(N__12116),
            .I(N__12113));
    Span12Mux_h I__2152 (
            .O(N__12113),
            .I(N__12110));
    Odrv12 I__2151 (
            .O(N__12110),
            .I(M_this_vga_signals_address_6));
    InMux I__2150 (
            .O(N__12107),
            .I(N__12104));
    LocalMux I__2149 (
            .O(N__12104),
            .I(\this_vga_signals.N_4 ));
    CascadeMux I__2148 (
            .O(N__12101),
            .I(\this_vram.M_this_vram_read_data_1_cascade_ ));
    IoInMux I__2147 (
            .O(N__12098),
            .I(N__12095));
    LocalMux I__2146 (
            .O(N__12095),
            .I(N__12092));
    IoSpan4Mux I__2145 (
            .O(N__12092),
            .I(N__12089));
    IoSpan4Mux I__2144 (
            .O(N__12089),
            .I(N__12085));
    IoInMux I__2143 (
            .O(N__12088),
            .I(N__12082));
    Sp12to4 I__2142 (
            .O(N__12085),
            .I(N__12077));
    LocalMux I__2141 (
            .O(N__12082),
            .I(N__12077));
    Span12Mux_s6_h I__2140 (
            .O(N__12077),
            .I(N__12074));
    Odrv12 I__2139 (
            .O(N__12074),
            .I(rgb_c_2));
    CascadeMux I__2138 (
            .O(N__12071),
            .I(N__12068));
    InMux I__2137 (
            .O(N__12068),
            .I(N__12065));
    LocalMux I__2136 (
            .O(N__12065),
            .I(N__12062));
    Odrv4 I__2135 (
            .O(N__12062),
            .I(\this_vga_signals.g0_4 ));
    InMux I__2134 (
            .O(N__12059),
            .I(N__12056));
    LocalMux I__2133 (
            .O(N__12056),
            .I(N__12053));
    Odrv4 I__2132 (
            .O(N__12053),
            .I(\this_vga_signals.if_N_8_mux_2_2_1 ));
    CascadeMux I__2131 (
            .O(N__12050),
            .I(\this_vga_signals.N_3_1_0_1_cascade_ ));
    InMux I__2130 (
            .O(N__12047),
            .I(N__12044));
    LocalMux I__2129 (
            .O(N__12044),
            .I(\this_vga_signals.g1_2_0_0 ));
    InMux I__2128 (
            .O(N__12041),
            .I(N__12038));
    LocalMux I__2127 (
            .O(N__12038),
            .I(\this_vga_signals.g0_0_0_0 ));
    CascadeMux I__2126 (
            .O(N__12035),
            .I(N__12026));
    CascadeMux I__2125 (
            .O(N__12034),
            .I(N__12018));
    InMux I__2124 (
            .O(N__12033),
            .I(N__12014));
    InMux I__2123 (
            .O(N__12032),
            .I(N__12009));
    InMux I__2122 (
            .O(N__12031),
            .I(N__12004));
    InMux I__2121 (
            .O(N__12030),
            .I(N__12004));
    CascadeMux I__2120 (
            .O(N__12029),
            .I(N__12001));
    InMux I__2119 (
            .O(N__12026),
            .I(N__11997));
    CascadeMux I__2118 (
            .O(N__12025),
            .I(N__11990));
    InMux I__2117 (
            .O(N__12024),
            .I(N__11986));
    InMux I__2116 (
            .O(N__12023),
            .I(N__11983));
    InMux I__2115 (
            .O(N__12022),
            .I(N__11978));
    InMux I__2114 (
            .O(N__12021),
            .I(N__11978));
    InMux I__2113 (
            .O(N__12018),
            .I(N__11973));
    InMux I__2112 (
            .O(N__12017),
            .I(N__11973));
    LocalMux I__2111 (
            .O(N__12014),
            .I(N__11970));
    InMux I__2110 (
            .O(N__12013),
            .I(N__11965));
    InMux I__2109 (
            .O(N__12012),
            .I(N__11965));
    LocalMux I__2108 (
            .O(N__12009),
            .I(N__11960));
    LocalMux I__2107 (
            .O(N__12004),
            .I(N__11960));
    InMux I__2106 (
            .O(N__12001),
            .I(N__11955));
    InMux I__2105 (
            .O(N__12000),
            .I(N__11955));
    LocalMux I__2104 (
            .O(N__11997),
            .I(N__11950));
    InMux I__2103 (
            .O(N__11996),
            .I(N__11943));
    InMux I__2102 (
            .O(N__11995),
            .I(N__11943));
    InMux I__2101 (
            .O(N__11994),
            .I(N__11943));
    InMux I__2100 (
            .O(N__11993),
            .I(N__11940));
    InMux I__2099 (
            .O(N__11990),
            .I(N__11935));
    InMux I__2098 (
            .O(N__11989),
            .I(N__11935));
    LocalMux I__2097 (
            .O(N__11986),
            .I(N__11930));
    LocalMux I__2096 (
            .O(N__11983),
            .I(N__11930));
    LocalMux I__2095 (
            .O(N__11978),
            .I(N__11925));
    LocalMux I__2094 (
            .O(N__11973),
            .I(N__11925));
    Span4Mux_h I__2093 (
            .O(N__11970),
            .I(N__11916));
    LocalMux I__2092 (
            .O(N__11965),
            .I(N__11916));
    Span4Mux_v I__2091 (
            .O(N__11960),
            .I(N__11916));
    LocalMux I__2090 (
            .O(N__11955),
            .I(N__11916));
    InMux I__2089 (
            .O(N__11954),
            .I(N__11913));
    InMux I__2088 (
            .O(N__11953),
            .I(N__11910));
    Span4Mux_h I__2087 (
            .O(N__11950),
            .I(N__11901));
    LocalMux I__2086 (
            .O(N__11943),
            .I(N__11901));
    LocalMux I__2085 (
            .O(N__11940),
            .I(N__11901));
    LocalMux I__2084 (
            .O(N__11935),
            .I(N__11901));
    Span4Mux_h I__2083 (
            .O(N__11930),
            .I(N__11896));
    Span4Mux_v I__2082 (
            .O(N__11925),
            .I(N__11896));
    Span4Mux_h I__2081 (
            .O(N__11916),
            .I(N__11893));
    LocalMux I__2080 (
            .O(N__11913),
            .I(\this_vga_signals.if_m1_0_0 ));
    LocalMux I__2079 (
            .O(N__11910),
            .I(\this_vga_signals.if_m1_0_0 ));
    Odrv4 I__2078 (
            .O(N__11901),
            .I(\this_vga_signals.if_m1_0_0 ));
    Odrv4 I__2077 (
            .O(N__11896),
            .I(\this_vga_signals.if_m1_0_0 ));
    Odrv4 I__2076 (
            .O(N__11893),
            .I(\this_vga_signals.if_m1_0_0 ));
    InMux I__2075 (
            .O(N__11882),
            .I(N__11878));
    InMux I__2074 (
            .O(N__11881),
            .I(N__11875));
    LocalMux I__2073 (
            .O(N__11878),
            .I(\this_vga_signals.N_21 ));
    LocalMux I__2072 (
            .O(N__11875),
            .I(\this_vga_signals.N_21 ));
    CascadeMux I__2071 (
            .O(N__11870),
            .I(N__11866));
    InMux I__2070 (
            .O(N__11869),
            .I(N__11861));
    InMux I__2069 (
            .O(N__11866),
            .I(N__11856));
    InMux I__2068 (
            .O(N__11865),
            .I(N__11856));
    InMux I__2067 (
            .O(N__11864),
            .I(N__11853));
    LocalMux I__2066 (
            .O(N__11861),
            .I(N__11848));
    LocalMux I__2065 (
            .O(N__11856),
            .I(N__11841));
    LocalMux I__2064 (
            .O(N__11853),
            .I(N__11828));
    InMux I__2063 (
            .O(N__11852),
            .I(N__11823));
    InMux I__2062 (
            .O(N__11851),
            .I(N__11823));
    Span4Mux_h I__2061 (
            .O(N__11848),
            .I(N__11820));
    InMux I__2060 (
            .O(N__11847),
            .I(N__11817));
    InMux I__2059 (
            .O(N__11846),
            .I(N__11810));
    InMux I__2058 (
            .O(N__11845),
            .I(N__11810));
    InMux I__2057 (
            .O(N__11844),
            .I(N__11810));
    Span4Mux_h I__2056 (
            .O(N__11841),
            .I(N__11807));
    InMux I__2055 (
            .O(N__11840),
            .I(N__11802));
    InMux I__2054 (
            .O(N__11839),
            .I(N__11802));
    InMux I__2053 (
            .O(N__11838),
            .I(N__11795));
    InMux I__2052 (
            .O(N__11837),
            .I(N__11795));
    InMux I__2051 (
            .O(N__11836),
            .I(N__11795));
    InMux I__2050 (
            .O(N__11835),
            .I(N__11792));
    InMux I__2049 (
            .O(N__11834),
            .I(N__11783));
    InMux I__2048 (
            .O(N__11833),
            .I(N__11783));
    InMux I__2047 (
            .O(N__11832),
            .I(N__11783));
    InMux I__2046 (
            .O(N__11831),
            .I(N__11783));
    Odrv4 I__2045 (
            .O(N__11828),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ));
    LocalMux I__2044 (
            .O(N__11823),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ));
    Odrv4 I__2043 (
            .O(N__11820),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ));
    LocalMux I__2042 (
            .O(N__11817),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ));
    LocalMux I__2041 (
            .O(N__11810),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ));
    Odrv4 I__2040 (
            .O(N__11807),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ));
    LocalMux I__2039 (
            .O(N__11802),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ));
    LocalMux I__2038 (
            .O(N__11795),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ));
    LocalMux I__2037 (
            .O(N__11792),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ));
    LocalMux I__2036 (
            .O(N__11783),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ));
    CascadeMux I__2035 (
            .O(N__11762),
            .I(N__11757));
    CascadeMux I__2034 (
            .O(N__11761),
            .I(N__11752));
    InMux I__2033 (
            .O(N__11760),
            .I(N__11749));
    InMux I__2032 (
            .O(N__11757),
            .I(N__11744));
    InMux I__2031 (
            .O(N__11756),
            .I(N__11735));
    InMux I__2030 (
            .O(N__11755),
            .I(N__11735));
    InMux I__2029 (
            .O(N__11752),
            .I(N__11735));
    LocalMux I__2028 (
            .O(N__11749),
            .I(N__11732));
    CascadeMux I__2027 (
            .O(N__11748),
            .I(N__11729));
    CascadeMux I__2026 (
            .O(N__11747),
            .I(N__11725));
    LocalMux I__2025 (
            .O(N__11744),
            .I(N__11719));
    InMux I__2024 (
            .O(N__11743),
            .I(N__11714));
    InMux I__2023 (
            .O(N__11742),
            .I(N__11714));
    LocalMux I__2022 (
            .O(N__11735),
            .I(N__11711));
    Span4Mux_h I__2021 (
            .O(N__11732),
            .I(N__11708));
    InMux I__2020 (
            .O(N__11729),
            .I(N__11701));
    InMux I__2019 (
            .O(N__11728),
            .I(N__11701));
    InMux I__2018 (
            .O(N__11725),
            .I(N__11701));
    InMux I__2017 (
            .O(N__11724),
            .I(N__11698));
    InMux I__2016 (
            .O(N__11723),
            .I(N__11693));
    InMux I__2015 (
            .O(N__11722),
            .I(N__11693));
    Odrv4 I__2014 (
            .O(N__11719),
            .I(\this_vga_signals.mult1_un61_sum_ac0_5 ));
    LocalMux I__2013 (
            .O(N__11714),
            .I(\this_vga_signals.mult1_un61_sum_ac0_5 ));
    Odrv4 I__2012 (
            .O(N__11711),
            .I(\this_vga_signals.mult1_un61_sum_ac0_5 ));
    Odrv4 I__2011 (
            .O(N__11708),
            .I(\this_vga_signals.mult1_un61_sum_ac0_5 ));
    LocalMux I__2010 (
            .O(N__11701),
            .I(\this_vga_signals.mult1_un61_sum_ac0_5 ));
    LocalMux I__2009 (
            .O(N__11698),
            .I(\this_vga_signals.mult1_un61_sum_ac0_5 ));
    LocalMux I__2008 (
            .O(N__11693),
            .I(\this_vga_signals.mult1_un61_sum_ac0_5 ));
    InMux I__2007 (
            .O(N__11678),
            .I(N__11673));
    InMux I__2006 (
            .O(N__11677),
            .I(N__11670));
    InMux I__2005 (
            .O(N__11676),
            .I(N__11667));
    LocalMux I__2004 (
            .O(N__11673),
            .I(\this_vga_signals.N_12 ));
    LocalMux I__2003 (
            .O(N__11670),
            .I(\this_vga_signals.N_12 ));
    LocalMux I__2002 (
            .O(N__11667),
            .I(\this_vga_signals.N_12 ));
    CascadeMux I__2001 (
            .O(N__11660),
            .I(\this_vga_signals.g0_0_0_a2_1_0_cascade_ ));
    CascadeMux I__2000 (
            .O(N__11657),
            .I(\this_vga_signals.if_N_3_2_i_3_1_cascade_ ));
    CascadeMux I__1999 (
            .O(N__11654),
            .I(N__11651));
    InMux I__1998 (
            .O(N__11651),
            .I(N__11648));
    LocalMux I__1997 (
            .O(N__11648),
            .I(\this_vga_signals.N_31 ));
    InMux I__1996 (
            .O(N__11645),
            .I(N__11642));
    LocalMux I__1995 (
            .O(N__11642),
            .I(\this_vga_signals.N_20_i_i ));
    CascadeMux I__1994 (
            .O(N__11639),
            .I(\this_vga_signals.N_20_i_i_cascade_ ));
    InMux I__1993 (
            .O(N__11636),
            .I(N__11633));
    LocalMux I__1992 (
            .O(N__11633),
            .I(N__11630));
    Odrv4 I__1991 (
            .O(N__11630),
            .I(\this_vga_signals.N_26_i_i ));
    InMux I__1990 (
            .O(N__11627),
            .I(N__11624));
    LocalMux I__1989 (
            .O(N__11624),
            .I(N__11619));
    InMux I__1988 (
            .O(N__11623),
            .I(N__11616));
    InMux I__1987 (
            .O(N__11622),
            .I(N__11608));
    Span4Mux_h I__1986 (
            .O(N__11619),
            .I(N__11603));
    LocalMux I__1985 (
            .O(N__11616),
            .I(N__11603));
    InMux I__1984 (
            .O(N__11615),
            .I(N__11600));
    InMux I__1983 (
            .O(N__11614),
            .I(N__11595));
    InMux I__1982 (
            .O(N__11613),
            .I(N__11595));
    InMux I__1981 (
            .O(N__11612),
            .I(N__11592));
    InMux I__1980 (
            .O(N__11611),
            .I(N__11589));
    LocalMux I__1979 (
            .O(N__11608),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    Odrv4 I__1978 (
            .O(N__11603),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1977 (
            .O(N__11600),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1976 (
            .O(N__11595),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1975 (
            .O(N__11592),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1974 (
            .O(N__11589),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    InMux I__1973 (
            .O(N__11576),
            .I(N__11573));
    LocalMux I__1972 (
            .O(N__11573),
            .I(N__11569));
    InMux I__1971 (
            .O(N__11572),
            .I(N__11566));
    Span4Mux_h I__1970 (
            .O(N__11569),
            .I(N__11557));
    LocalMux I__1969 (
            .O(N__11566),
            .I(N__11557));
    InMux I__1968 (
            .O(N__11565),
            .I(N__11554));
    InMux I__1967 (
            .O(N__11564),
            .I(N__11547));
    InMux I__1966 (
            .O(N__11563),
            .I(N__11547));
    InMux I__1965 (
            .O(N__11562),
            .I(N__11547));
    Odrv4 I__1964 (
            .O(N__11557),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1 ));
    LocalMux I__1963 (
            .O(N__11554),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1 ));
    LocalMux I__1962 (
            .O(N__11547),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1 ));
    InMux I__1961 (
            .O(N__11540),
            .I(N__11536));
    InMux I__1960 (
            .O(N__11539),
            .I(N__11533));
    LocalMux I__1959 (
            .O(N__11536),
            .I(N__11530));
    LocalMux I__1958 (
            .O(N__11533),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    Odrv4 I__1957 (
            .O(N__11530),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    InMux I__1956 (
            .O(N__11525),
            .I(N__11521));
    InMux I__1955 (
            .O(N__11524),
            .I(N__11518));
    LocalMux I__1954 (
            .O(N__11521),
            .I(N__11515));
    LocalMux I__1953 (
            .O(N__11518),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    Odrv4 I__1952 (
            .O(N__11515),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    CascadeMux I__1951 (
            .O(N__11510),
            .I(N__11507));
    CascadeBuf I__1950 (
            .O(N__11507),
            .I(N__11504));
    CascadeMux I__1949 (
            .O(N__11504),
            .I(N__11501));
    CascadeBuf I__1948 (
            .O(N__11501),
            .I(N__11498));
    CascadeMux I__1947 (
            .O(N__11498),
            .I(N__11495));
    CascadeBuf I__1946 (
            .O(N__11495),
            .I(N__11492));
    CascadeMux I__1945 (
            .O(N__11492),
            .I(N__11489));
    CascadeBuf I__1944 (
            .O(N__11489),
            .I(N__11486));
    CascadeMux I__1943 (
            .O(N__11486),
            .I(N__11483));
    CascadeBuf I__1942 (
            .O(N__11483),
            .I(N__11480));
    CascadeMux I__1941 (
            .O(N__11480),
            .I(N__11477));
    CascadeBuf I__1940 (
            .O(N__11477),
            .I(N__11474));
    CascadeMux I__1939 (
            .O(N__11474),
            .I(N__11471));
    CascadeBuf I__1938 (
            .O(N__11471),
            .I(N__11468));
    CascadeMux I__1937 (
            .O(N__11468),
            .I(N__11465));
    CascadeBuf I__1936 (
            .O(N__11465),
            .I(N__11462));
    CascadeMux I__1935 (
            .O(N__11462),
            .I(N__11459));
    CascadeBuf I__1934 (
            .O(N__11459),
            .I(N__11456));
    CascadeMux I__1933 (
            .O(N__11456),
            .I(N__11453));
    CascadeBuf I__1932 (
            .O(N__11453),
            .I(N__11450));
    CascadeMux I__1931 (
            .O(N__11450),
            .I(N__11447));
    CascadeBuf I__1930 (
            .O(N__11447),
            .I(N__11444));
    CascadeMux I__1929 (
            .O(N__11444),
            .I(N__11441));
    CascadeBuf I__1928 (
            .O(N__11441),
            .I(N__11438));
    CascadeMux I__1927 (
            .O(N__11438),
            .I(N__11435));
    CascadeBuf I__1926 (
            .O(N__11435),
            .I(N__11432));
    CascadeMux I__1925 (
            .O(N__11432),
            .I(N__11429));
    CascadeBuf I__1924 (
            .O(N__11429),
            .I(N__11426));
    CascadeMux I__1923 (
            .O(N__11426),
            .I(N__11423));
    CascadeBuf I__1922 (
            .O(N__11423),
            .I(N__11420));
    CascadeMux I__1921 (
            .O(N__11420),
            .I(N__11417));
    InMux I__1920 (
            .O(N__11417),
            .I(N__11414));
    LocalMux I__1919 (
            .O(N__11414),
            .I(N__11411));
    Span12Mux_h I__1918 (
            .O(N__11411),
            .I(N__11408));
    Odrv12 I__1917 (
            .O(N__11408),
            .I(M_this_vga_signals_address_9));
    InMux I__1916 (
            .O(N__11405),
            .I(N__11402));
    LocalMux I__1915 (
            .O(N__11402),
            .I(N__11398));
    InMux I__1914 (
            .O(N__11401),
            .I(N__11395));
    Span4Mux_v I__1913 (
            .O(N__11398),
            .I(N__11390));
    LocalMux I__1912 (
            .O(N__11395),
            .I(N__11387));
    InMux I__1911 (
            .O(N__11394),
            .I(N__11382));
    InMux I__1910 (
            .O(N__11393),
            .I(N__11382));
    Odrv4 I__1909 (
            .O(N__11390),
            .I(\this_vga_signals.mult1_un54_sum_ac0_7 ));
    Odrv4 I__1908 (
            .O(N__11387),
            .I(\this_vga_signals.mult1_un54_sum_ac0_7 ));
    LocalMux I__1907 (
            .O(N__11382),
            .I(\this_vga_signals.mult1_un54_sum_ac0_7 ));
    InMux I__1906 (
            .O(N__11375),
            .I(N__11372));
    LocalMux I__1905 (
            .O(N__11372),
            .I(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_4 ));
    InMux I__1904 (
            .O(N__11369),
            .I(N__11366));
    LocalMux I__1903 (
            .O(N__11366),
            .I(\this_vga_signals.g0_i_x4_4_a3_1 ));
    InMux I__1902 (
            .O(N__11363),
            .I(N__11360));
    LocalMux I__1901 (
            .O(N__11360),
            .I(N__11357));
    Odrv4 I__1900 (
            .O(N__11357),
            .I(\this_vga_signals.if_m1_0 ));
    InMux I__1899 (
            .O(N__11354),
            .I(N__11351));
    LocalMux I__1898 (
            .O(N__11351),
            .I(\this_vga_signals.if_N_3_3_i ));
    CascadeMux I__1897 (
            .O(N__11348),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5_cascade_));
    CascadeMux I__1896 (
            .O(N__11345),
            .I(\this_vga_signals.if_N_3_2_i_cascade_ ));
    CascadeMux I__1895 (
            .O(N__11342),
            .I(N__11339));
    CascadeBuf I__1894 (
            .O(N__11339),
            .I(N__11336));
    CascadeMux I__1893 (
            .O(N__11336),
            .I(N__11333));
    CascadeBuf I__1892 (
            .O(N__11333),
            .I(N__11330));
    CascadeMux I__1891 (
            .O(N__11330),
            .I(N__11327));
    CascadeBuf I__1890 (
            .O(N__11327),
            .I(N__11324));
    CascadeMux I__1889 (
            .O(N__11324),
            .I(N__11321));
    CascadeBuf I__1888 (
            .O(N__11321),
            .I(N__11318));
    CascadeMux I__1887 (
            .O(N__11318),
            .I(N__11315));
    CascadeBuf I__1886 (
            .O(N__11315),
            .I(N__11312));
    CascadeMux I__1885 (
            .O(N__11312),
            .I(N__11309));
    CascadeBuf I__1884 (
            .O(N__11309),
            .I(N__11306));
    CascadeMux I__1883 (
            .O(N__11306),
            .I(N__11303));
    CascadeBuf I__1882 (
            .O(N__11303),
            .I(N__11300));
    CascadeMux I__1881 (
            .O(N__11300),
            .I(N__11297));
    CascadeBuf I__1880 (
            .O(N__11297),
            .I(N__11294));
    CascadeMux I__1879 (
            .O(N__11294),
            .I(N__11291));
    CascadeBuf I__1878 (
            .O(N__11291),
            .I(N__11288));
    CascadeMux I__1877 (
            .O(N__11288),
            .I(N__11285));
    CascadeBuf I__1876 (
            .O(N__11285),
            .I(N__11282));
    CascadeMux I__1875 (
            .O(N__11282),
            .I(N__11279));
    CascadeBuf I__1874 (
            .O(N__11279),
            .I(N__11276));
    CascadeMux I__1873 (
            .O(N__11276),
            .I(N__11273));
    CascadeBuf I__1872 (
            .O(N__11273),
            .I(N__11270));
    CascadeMux I__1871 (
            .O(N__11270),
            .I(N__11267));
    CascadeBuf I__1870 (
            .O(N__11267),
            .I(N__11264));
    CascadeMux I__1869 (
            .O(N__11264),
            .I(N__11261));
    CascadeBuf I__1868 (
            .O(N__11261),
            .I(N__11258));
    CascadeMux I__1867 (
            .O(N__11258),
            .I(N__11255));
    CascadeBuf I__1866 (
            .O(N__11255),
            .I(N__11252));
    CascadeMux I__1865 (
            .O(N__11252),
            .I(N__11249));
    InMux I__1864 (
            .O(N__11249),
            .I(N__11246));
    LocalMux I__1863 (
            .O(N__11246),
            .I(N__11243));
    Span12Mux_s9_h I__1862 (
            .O(N__11243),
            .I(N__11240));
    Span12Mux_v I__1861 (
            .O(N__11240),
            .I(N__11237));
    Odrv12 I__1860 (
            .O(N__11237),
            .I(M_this_vga_signals_address_3));
    CascadeMux I__1859 (
            .O(N__11234),
            .I(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_3L3_cascade_ ));
    InMux I__1858 (
            .O(N__11231),
            .I(N__11228));
    LocalMux I__1857 (
            .O(N__11228),
            .I(N__11225));
    Span4Mux_v I__1856 (
            .O(N__11225),
            .I(N__11222));
    Odrv4 I__1855 (
            .O(N__11222),
            .I(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_2L1 ));
    CascadeMux I__1854 (
            .O(N__11219),
            .I(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5_cascade_ ));
    InMux I__1853 (
            .O(N__11216),
            .I(N__11213));
    LocalMux I__1852 (
            .O(N__11213),
            .I(\this_vga_signals.N_21_0 ));
    CascadeMux I__1851 (
            .O(N__11210),
            .I(N__11207));
    InMux I__1850 (
            .O(N__11207),
            .I(N__11204));
    LocalMux I__1849 (
            .O(N__11204),
            .I(N__11201));
    Odrv4 I__1848 (
            .O(N__11201),
            .I(\this_vga_signals.g0_6_0_0_2 ));
    InMux I__1847 (
            .O(N__11198),
            .I(N__11195));
    LocalMux I__1846 (
            .O(N__11195),
            .I(\this_vga_signals.if_N_8_mux_2_2 ));
    CascadeMux I__1845 (
            .O(N__11192),
            .I(\this_vga_signals.mult1_un82_sum_axb3_cascade_ ));
    CascadeMux I__1844 (
            .O(N__11189),
            .I(\this_vga_signals.address_i2_mux_cascade_ ));
    InMux I__1843 (
            .O(N__11186),
            .I(N__11183));
    LocalMux I__1842 (
            .O(N__11183),
            .I(\this_vga_signals.address_N_11 ));
    InMux I__1841 (
            .O(N__11180),
            .I(N__11177));
    LocalMux I__1840 (
            .O(N__11177),
            .I(\this_vga_signals.address_i2_mux_0 ));
    CascadeMux I__1839 (
            .O(N__11174),
            .I(\this_vga_signals.address_m21_ns_1_cascade_ ));
    InMux I__1838 (
            .O(N__11171),
            .I(N__11168));
    LocalMux I__1837 (
            .O(N__11168),
            .I(\this_vga_signals.address_i2_mux_1 ));
    CascadeMux I__1836 (
            .O(N__11165),
            .I(\this_vga_signals.address_N_22_cascade_ ));
    InMux I__1835 (
            .O(N__11162),
            .I(N__11159));
    LocalMux I__1834 (
            .O(N__11159),
            .I(\this_vga_signals.address_N_36 ));
    CascadeMux I__1833 (
            .O(N__11156),
            .I(N__11153));
    CascadeBuf I__1832 (
            .O(N__11153),
            .I(N__11150));
    CascadeMux I__1831 (
            .O(N__11150),
            .I(N__11147));
    CascadeBuf I__1830 (
            .O(N__11147),
            .I(N__11144));
    CascadeMux I__1829 (
            .O(N__11144),
            .I(N__11141));
    CascadeBuf I__1828 (
            .O(N__11141),
            .I(N__11138));
    CascadeMux I__1827 (
            .O(N__11138),
            .I(N__11135));
    CascadeBuf I__1826 (
            .O(N__11135),
            .I(N__11132));
    CascadeMux I__1825 (
            .O(N__11132),
            .I(N__11129));
    CascadeBuf I__1824 (
            .O(N__11129),
            .I(N__11126));
    CascadeMux I__1823 (
            .O(N__11126),
            .I(N__11123));
    CascadeBuf I__1822 (
            .O(N__11123),
            .I(N__11120));
    CascadeMux I__1821 (
            .O(N__11120),
            .I(N__11117));
    CascadeBuf I__1820 (
            .O(N__11117),
            .I(N__11114));
    CascadeMux I__1819 (
            .O(N__11114),
            .I(N__11111));
    CascadeBuf I__1818 (
            .O(N__11111),
            .I(N__11108));
    CascadeMux I__1817 (
            .O(N__11108),
            .I(N__11105));
    CascadeBuf I__1816 (
            .O(N__11105),
            .I(N__11102));
    CascadeMux I__1815 (
            .O(N__11102),
            .I(N__11099));
    CascadeBuf I__1814 (
            .O(N__11099),
            .I(N__11096));
    CascadeMux I__1813 (
            .O(N__11096),
            .I(N__11093));
    CascadeBuf I__1812 (
            .O(N__11093),
            .I(N__11090));
    CascadeMux I__1811 (
            .O(N__11090),
            .I(N__11087));
    CascadeBuf I__1810 (
            .O(N__11087),
            .I(N__11084));
    CascadeMux I__1809 (
            .O(N__11084),
            .I(N__11081));
    CascadeBuf I__1808 (
            .O(N__11081),
            .I(N__11078));
    CascadeMux I__1807 (
            .O(N__11078),
            .I(N__11075));
    CascadeBuf I__1806 (
            .O(N__11075),
            .I(N__11072));
    CascadeMux I__1805 (
            .O(N__11072),
            .I(N__11069));
    CascadeBuf I__1804 (
            .O(N__11069),
            .I(N__11066));
    CascadeMux I__1803 (
            .O(N__11066),
            .I(N__11063));
    InMux I__1802 (
            .O(N__11063),
            .I(N__11060));
    LocalMux I__1801 (
            .O(N__11060),
            .I(N__11057));
    Sp12to4 I__1800 (
            .O(N__11057),
            .I(N__11054));
    Span12Mux_s9_v I__1799 (
            .O(N__11054),
            .I(N__11051));
    Odrv12 I__1798 (
            .O(N__11051),
            .I(M_this_vga_signals_address_7));
    InMux I__1797 (
            .O(N__11048),
            .I(N__11043));
    InMux I__1796 (
            .O(N__11047),
            .I(N__11038));
    InMux I__1795 (
            .O(N__11046),
            .I(N__11038));
    LocalMux I__1794 (
            .O(N__11043),
            .I(N__11035));
    LocalMux I__1793 (
            .O(N__11038),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    Odrv4 I__1792 (
            .O(N__11035),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    InMux I__1791 (
            .O(N__11030),
            .I(N__11020));
    InMux I__1790 (
            .O(N__11029),
            .I(N__11017));
    InMux I__1789 (
            .O(N__11028),
            .I(N__11011));
    InMux I__1788 (
            .O(N__11027),
            .I(N__11011));
    InMux I__1787 (
            .O(N__11026),
            .I(N__11008));
    InMux I__1786 (
            .O(N__11025),
            .I(N__11005));
    CascadeMux I__1785 (
            .O(N__11024),
            .I(N__10999));
    InMux I__1784 (
            .O(N__11023),
            .I(N__10994));
    LocalMux I__1783 (
            .O(N__11020),
            .I(N__10987));
    LocalMux I__1782 (
            .O(N__11017),
            .I(N__10987));
    CascadeMux I__1781 (
            .O(N__11016),
            .I(N__10983));
    LocalMux I__1780 (
            .O(N__11011),
            .I(N__10978));
    LocalMux I__1779 (
            .O(N__11008),
            .I(N__10978));
    LocalMux I__1778 (
            .O(N__11005),
            .I(N__10975));
    InMux I__1777 (
            .O(N__11004),
            .I(N__10972));
    InMux I__1776 (
            .O(N__11003),
            .I(N__10969));
    InMux I__1775 (
            .O(N__11002),
            .I(N__10966));
    InMux I__1774 (
            .O(N__10999),
            .I(N__10959));
    InMux I__1773 (
            .O(N__10998),
            .I(N__10959));
    InMux I__1772 (
            .O(N__10997),
            .I(N__10959));
    LocalMux I__1771 (
            .O(N__10994),
            .I(N__10956));
    InMux I__1770 (
            .O(N__10993),
            .I(N__10951));
    InMux I__1769 (
            .O(N__10992),
            .I(N__10951));
    Span4Mux_h I__1768 (
            .O(N__10987),
            .I(N__10948));
    InMux I__1767 (
            .O(N__10986),
            .I(N__10943));
    InMux I__1766 (
            .O(N__10983),
            .I(N__10943));
    Odrv4 I__1765 (
            .O(N__10978),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__1764 (
            .O(N__10975),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__1763 (
            .O(N__10972),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__1762 (
            .O(N__10969),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__1761 (
            .O(N__10966),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__1760 (
            .O(N__10959),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__1759 (
            .O(N__10956),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__1758 (
            .O(N__10951),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__1757 (
            .O(N__10948),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__1756 (
            .O(N__10943),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    InMux I__1755 (
            .O(N__10922),
            .I(N__10918));
    CascadeMux I__1754 (
            .O(N__10921),
            .I(N__10914));
    LocalMux I__1753 (
            .O(N__10918),
            .I(N__10910));
    InMux I__1752 (
            .O(N__10917),
            .I(N__10905));
    InMux I__1751 (
            .O(N__10914),
            .I(N__10905));
    CascadeMux I__1750 (
            .O(N__10913),
            .I(N__10900));
    Span4Mux_h I__1749 (
            .O(N__10910),
            .I(N__10895));
    LocalMux I__1748 (
            .O(N__10905),
            .I(N__10895));
    InMux I__1747 (
            .O(N__10904),
            .I(N__10890));
    InMux I__1746 (
            .O(N__10903),
            .I(N__10890));
    InMux I__1745 (
            .O(N__10900),
            .I(N__10887));
    Span4Mux_h I__1744 (
            .O(N__10895),
            .I(N__10884));
    LocalMux I__1743 (
            .O(N__10890),
            .I(N__10881));
    LocalMux I__1742 (
            .O(N__10887),
            .I(N__10878));
    Odrv4 I__1741 (
            .O(N__10884),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__1740 (
            .O(N__10881),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__1739 (
            .O(N__10878),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    CascadeMux I__1738 (
            .O(N__10871),
            .I(N__10865));
    InMux I__1737 (
            .O(N__10870),
            .I(N__10857));
    InMux I__1736 (
            .O(N__10869),
            .I(N__10857));
    InMux I__1735 (
            .O(N__10868),
            .I(N__10857));
    InMux I__1734 (
            .O(N__10865),
            .I(N__10853));
    InMux I__1733 (
            .O(N__10864),
            .I(N__10850));
    LocalMux I__1732 (
            .O(N__10857),
            .I(N__10847));
    InMux I__1731 (
            .O(N__10856),
            .I(N__10844));
    LocalMux I__1730 (
            .O(N__10853),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_0 ));
    LocalMux I__1729 (
            .O(N__10850),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_0 ));
    Odrv4 I__1728 (
            .O(N__10847),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_0 ));
    LocalMux I__1727 (
            .O(N__10844),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_0 ));
    InMux I__1726 (
            .O(N__10835),
            .I(N__10832));
    LocalMux I__1725 (
            .O(N__10832),
            .I(\this_vga_signals.if_m16_0_o4 ));
    InMux I__1724 (
            .O(N__10829),
            .I(N__10824));
    InMux I__1723 (
            .O(N__10828),
            .I(N__10818));
    InMux I__1722 (
            .O(N__10827),
            .I(N__10815));
    LocalMux I__1721 (
            .O(N__10824),
            .I(N__10810));
    InMux I__1720 (
            .O(N__10823),
            .I(N__10807));
    InMux I__1719 (
            .O(N__10822),
            .I(N__10804));
    InMux I__1718 (
            .O(N__10821),
            .I(N__10801));
    LocalMux I__1717 (
            .O(N__10818),
            .I(N__10798));
    LocalMux I__1716 (
            .O(N__10815),
            .I(N__10795));
    InMux I__1715 (
            .O(N__10814),
            .I(N__10792));
    InMux I__1714 (
            .O(N__10813),
            .I(N__10787));
    Span4Mux_h I__1713 (
            .O(N__10810),
            .I(N__10784));
    LocalMux I__1712 (
            .O(N__10807),
            .I(N__10781));
    LocalMux I__1711 (
            .O(N__10804),
            .I(N__10772));
    LocalMux I__1710 (
            .O(N__10801),
            .I(N__10772));
    Span4Mux_v I__1709 (
            .O(N__10798),
            .I(N__10772));
    Span4Mux_v I__1708 (
            .O(N__10795),
            .I(N__10772));
    LocalMux I__1707 (
            .O(N__10792),
            .I(N__10769));
    InMux I__1706 (
            .O(N__10791),
            .I(N__10766));
    InMux I__1705 (
            .O(N__10790),
            .I(N__10763));
    LocalMux I__1704 (
            .O(N__10787),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv4 I__1703 (
            .O(N__10784),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv4 I__1702 (
            .O(N__10781),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv4 I__1701 (
            .O(N__10772),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv4 I__1700 (
            .O(N__10769),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__1699 (
            .O(N__10766),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__1698 (
            .O(N__10763),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    CascadeMux I__1697 (
            .O(N__10748),
            .I(N__10736));
    InMux I__1696 (
            .O(N__10747),
            .I(N__10726));
    InMux I__1695 (
            .O(N__10746),
            .I(N__10726));
    InMux I__1694 (
            .O(N__10745),
            .I(N__10723));
    InMux I__1693 (
            .O(N__10744),
            .I(N__10720));
    InMux I__1692 (
            .O(N__10743),
            .I(N__10715));
    InMux I__1691 (
            .O(N__10742),
            .I(N__10715));
    InMux I__1690 (
            .O(N__10741),
            .I(N__10712));
    InMux I__1689 (
            .O(N__10740),
            .I(N__10709));
    InMux I__1688 (
            .O(N__10739),
            .I(N__10704));
    InMux I__1687 (
            .O(N__10736),
            .I(N__10704));
    CascadeMux I__1686 (
            .O(N__10735),
            .I(N__10701));
    InMux I__1685 (
            .O(N__10734),
            .I(N__10697));
    InMux I__1684 (
            .O(N__10733),
            .I(N__10694));
    InMux I__1683 (
            .O(N__10732),
            .I(N__10689));
    InMux I__1682 (
            .O(N__10731),
            .I(N__10689));
    LocalMux I__1681 (
            .O(N__10726),
            .I(N__10684));
    LocalMux I__1680 (
            .O(N__10723),
            .I(N__10684));
    LocalMux I__1679 (
            .O(N__10720),
            .I(N__10673));
    LocalMux I__1678 (
            .O(N__10715),
            .I(N__10673));
    LocalMux I__1677 (
            .O(N__10712),
            .I(N__10673));
    LocalMux I__1676 (
            .O(N__10709),
            .I(N__10673));
    LocalMux I__1675 (
            .O(N__10704),
            .I(N__10673));
    InMux I__1674 (
            .O(N__10701),
            .I(N__10670));
    CascadeMux I__1673 (
            .O(N__10700),
            .I(N__10661));
    LocalMux I__1672 (
            .O(N__10697),
            .I(N__10648));
    LocalMux I__1671 (
            .O(N__10694),
            .I(N__10648));
    LocalMux I__1670 (
            .O(N__10689),
            .I(N__10648));
    Span4Mux_v I__1669 (
            .O(N__10684),
            .I(N__10648));
    Span4Mux_v I__1668 (
            .O(N__10673),
            .I(N__10648));
    LocalMux I__1667 (
            .O(N__10670),
            .I(N__10648));
    InMux I__1666 (
            .O(N__10669),
            .I(N__10645));
    InMux I__1665 (
            .O(N__10668),
            .I(N__10638));
    InMux I__1664 (
            .O(N__10667),
            .I(N__10638));
    InMux I__1663 (
            .O(N__10666),
            .I(N__10638));
    InMux I__1662 (
            .O(N__10665),
            .I(N__10633));
    InMux I__1661 (
            .O(N__10664),
            .I(N__10633));
    InMux I__1660 (
            .O(N__10661),
            .I(N__10630));
    Odrv4 I__1659 (
            .O(N__10648),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__1658 (
            .O(N__10645),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__1657 (
            .O(N__10638),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__1656 (
            .O(N__10633),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__1655 (
            .O(N__10630),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    InMux I__1654 (
            .O(N__10619),
            .I(N__10616));
    LocalMux I__1653 (
            .O(N__10616),
            .I(N__10612));
    InMux I__1652 (
            .O(N__10615),
            .I(N__10609));
    Odrv4 I__1651 (
            .O(N__10612),
            .I(\this_vga_signals.address_N_40 ));
    LocalMux I__1650 (
            .O(N__10609),
            .I(\this_vga_signals.address_N_40 ));
    InMux I__1649 (
            .O(N__10604),
            .I(N__10601));
    LocalMux I__1648 (
            .O(N__10601),
            .I(N__10598));
    Odrv4 I__1647 (
            .O(N__10598),
            .I(\this_vga_signals.if_m4_0_1_0_0 ));
    CascadeMux I__1646 (
            .O(N__10595),
            .I(N_11_0_cascade_));
    InMux I__1645 (
            .O(N__10592),
            .I(N__10586));
    InMux I__1644 (
            .O(N__10591),
            .I(N__10586));
    LocalMux I__1643 (
            .O(N__10586),
            .I(\this_vga_signals.N_5_i ));
    InMux I__1642 (
            .O(N__10583),
            .I(N__10580));
    LocalMux I__1641 (
            .O(N__10580),
            .I(\this_vga_signals.G_12_0_1 ));
    InMux I__1640 (
            .O(N__10577),
            .I(N__10574));
    LocalMux I__1639 (
            .O(N__10574),
            .I(\this_vga_signals.N_25 ));
    InMux I__1638 (
            .O(N__10571),
            .I(N__10562));
    InMux I__1637 (
            .O(N__10570),
            .I(N__10562));
    InMux I__1636 (
            .O(N__10569),
            .I(N__10557));
    InMux I__1635 (
            .O(N__10568),
            .I(N__10557));
    InMux I__1634 (
            .O(N__10567),
            .I(N__10554));
    LocalMux I__1633 (
            .O(N__10562),
            .I(\this_vga_signals.M_vstate_qZ0Z_0 ));
    LocalMux I__1632 (
            .O(N__10557),
            .I(\this_vga_signals.M_vstate_qZ0Z_0 ));
    LocalMux I__1631 (
            .O(N__10554),
            .I(\this_vga_signals.M_vstate_qZ0Z_0 ));
    InMux I__1630 (
            .O(N__10547),
            .I(N__10540));
    InMux I__1629 (
            .O(N__10546),
            .I(N__10540));
    CascadeMux I__1628 (
            .O(N__10545),
            .I(N__10535));
    LocalMux I__1627 (
            .O(N__10540),
            .I(N__10532));
    InMux I__1626 (
            .O(N__10539),
            .I(N__10528));
    InMux I__1625 (
            .O(N__10538),
            .I(N__10523));
    InMux I__1624 (
            .O(N__10535),
            .I(N__10523));
    Span4Mux_h I__1623 (
            .O(N__10532),
            .I(N__10514));
    InMux I__1622 (
            .O(N__10531),
            .I(N__10511));
    LocalMux I__1621 (
            .O(N__10528),
            .I(N__10508));
    LocalMux I__1620 (
            .O(N__10523),
            .I(N__10505));
    InMux I__1619 (
            .O(N__10522),
            .I(N__10502));
    InMux I__1618 (
            .O(N__10521),
            .I(N__10499));
    InMux I__1617 (
            .O(N__10520),
            .I(N__10494));
    InMux I__1616 (
            .O(N__10519),
            .I(N__10494));
    InMux I__1615 (
            .O(N__10518),
            .I(N__10491));
    InMux I__1614 (
            .O(N__10517),
            .I(N__10488));
    Odrv4 I__1613 (
            .O(N__10514),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__1612 (
            .O(N__10511),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__1611 (
            .O(N__10508),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv12 I__1610 (
            .O(N__10505),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__1609 (
            .O(N__10502),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__1608 (
            .O(N__10499),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__1607 (
            .O(N__10494),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__1606 (
            .O(N__10491),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__1605 (
            .O(N__10488),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    InMux I__1604 (
            .O(N__10469),
            .I(N__10466));
    LocalMux I__1603 (
            .O(N__10466),
            .I(\this_vga_signals.N_275 ));
    CascadeMux I__1602 (
            .O(N__10463),
            .I(\this_vga_signals.if_N_9_i_i_cascade_ ));
    InMux I__1601 (
            .O(N__10460),
            .I(N__10457));
    LocalMux I__1600 (
            .O(N__10457),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    CascadeMux I__1599 (
            .O(N__10454),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_ ));
    CascadeMux I__1598 (
            .O(N__10451),
            .I(N__10448));
    CascadeBuf I__1597 (
            .O(N__10448),
            .I(N__10445));
    CascadeMux I__1596 (
            .O(N__10445),
            .I(N__10442));
    CascadeBuf I__1595 (
            .O(N__10442),
            .I(N__10439));
    CascadeMux I__1594 (
            .O(N__10439),
            .I(N__10436));
    CascadeBuf I__1593 (
            .O(N__10436),
            .I(N__10433));
    CascadeMux I__1592 (
            .O(N__10433),
            .I(N__10430));
    CascadeBuf I__1591 (
            .O(N__10430),
            .I(N__10427));
    CascadeMux I__1590 (
            .O(N__10427),
            .I(N__10424));
    CascadeBuf I__1589 (
            .O(N__10424),
            .I(N__10421));
    CascadeMux I__1588 (
            .O(N__10421),
            .I(N__10418));
    CascadeBuf I__1587 (
            .O(N__10418),
            .I(N__10415));
    CascadeMux I__1586 (
            .O(N__10415),
            .I(N__10412));
    CascadeBuf I__1585 (
            .O(N__10412),
            .I(N__10409));
    CascadeMux I__1584 (
            .O(N__10409),
            .I(N__10406));
    CascadeBuf I__1583 (
            .O(N__10406),
            .I(N__10403));
    CascadeMux I__1582 (
            .O(N__10403),
            .I(N__10400));
    CascadeBuf I__1581 (
            .O(N__10400),
            .I(N__10397));
    CascadeMux I__1580 (
            .O(N__10397),
            .I(N__10394));
    CascadeBuf I__1579 (
            .O(N__10394),
            .I(N__10391));
    CascadeMux I__1578 (
            .O(N__10391),
            .I(N__10388));
    CascadeBuf I__1577 (
            .O(N__10388),
            .I(N__10385));
    CascadeMux I__1576 (
            .O(N__10385),
            .I(N__10382));
    CascadeBuf I__1575 (
            .O(N__10382),
            .I(N__10379));
    CascadeMux I__1574 (
            .O(N__10379),
            .I(N__10376));
    CascadeBuf I__1573 (
            .O(N__10376),
            .I(N__10373));
    CascadeMux I__1572 (
            .O(N__10373),
            .I(N__10370));
    CascadeBuf I__1571 (
            .O(N__10370),
            .I(N__10367));
    CascadeMux I__1570 (
            .O(N__10367),
            .I(N__10364));
    CascadeBuf I__1569 (
            .O(N__10364),
            .I(N__10361));
    CascadeMux I__1568 (
            .O(N__10361),
            .I(N__10358));
    InMux I__1567 (
            .O(N__10358),
            .I(N__10355));
    LocalMux I__1566 (
            .O(N__10355),
            .I(N__10352));
    Span12Mux_s5_v I__1565 (
            .O(N__10352),
            .I(N__10349));
    Span12Mux_h I__1564 (
            .O(N__10349),
            .I(N__10346));
    Odrv12 I__1563 (
            .O(N__10346),
            .I(M_this_vga_signals_address_8));
    CascadeMux I__1562 (
            .O(N__10343),
            .I(\this_vga_signals.address_m6_0_1_cascade_ ));
    InMux I__1561 (
            .O(N__10340),
            .I(N__10336));
    InMux I__1560 (
            .O(N__10339),
            .I(N__10330));
    LocalMux I__1559 (
            .O(N__10336),
            .I(N__10327));
    InMux I__1558 (
            .O(N__10335),
            .I(N__10320));
    InMux I__1557 (
            .O(N__10334),
            .I(N__10320));
    InMux I__1556 (
            .O(N__10333),
            .I(N__10320));
    LocalMux I__1555 (
            .O(N__10330),
            .I(\this_vga_signals.address_mZ0Z1 ));
    Odrv4 I__1554 (
            .O(N__10327),
            .I(\this_vga_signals.address_mZ0Z1 ));
    LocalMux I__1553 (
            .O(N__10320),
            .I(\this_vga_signals.address_mZ0Z1 ));
    CascadeMux I__1552 (
            .O(N__10313),
            .I(\this_vga_signals.G_12_0_3_cascade_ ));
    InMux I__1551 (
            .O(N__10310),
            .I(N__10307));
    LocalMux I__1550 (
            .O(N__10307),
            .I(N__10303));
    InMux I__1549 (
            .O(N__10306),
            .I(N__10300));
    Odrv4 I__1548 (
            .O(N__10303),
            .I(\this_vga_signals.if_m4_0_1 ));
    LocalMux I__1547 (
            .O(N__10300),
            .I(\this_vga_signals.if_m4_0_1 ));
    CascadeMux I__1546 (
            .O(N__10295),
            .I(this_vga_signals_un17_address_if_N_8_mux_cascade_));
    InMux I__1545 (
            .O(N__10292),
            .I(N__10289));
    LocalMux I__1544 (
            .O(N__10289),
            .I(\this_vga_signals.N_10_0 ));
    CascadeMux I__1543 (
            .O(N__10286),
            .I(N_6_i_cascade_));
    InMux I__1542 (
            .O(N__10283),
            .I(N__10280));
    LocalMux I__1541 (
            .O(N__10280),
            .I(N__10277));
    Odrv4 I__1540 (
            .O(N__10277),
            .I(\this_vga_signals.N_18_0 ));
    InMux I__1539 (
            .O(N__10274),
            .I(N__10271));
    LocalMux I__1538 (
            .O(N__10271),
            .I(N__10268));
    Odrv4 I__1537 (
            .O(N__10268),
            .I(\this_vga_signals.g0_6_1 ));
    InMux I__1536 (
            .O(N__10265),
            .I(N__10262));
    LocalMux I__1535 (
            .O(N__10262),
            .I(\this_vga_signals.G_12_0_x3_0 ));
    InMux I__1534 (
            .O(N__10259),
            .I(N__10256));
    LocalMux I__1533 (
            .O(N__10256),
            .I(N__10253));
    Span4Mux_h I__1532 (
            .O(N__10253),
            .I(N__10250));
    Odrv4 I__1531 (
            .O(N__10250),
            .I(\this_vga_signals.g0_6_0_0_1 ));
    CascadeMux I__1530 (
            .O(N__10247),
            .I(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_));
    CascadeMux I__1529 (
            .O(N__10244),
            .I(N__10236));
    InMux I__1528 (
            .O(N__10243),
            .I(N__10231));
    InMux I__1527 (
            .O(N__10242),
            .I(N__10226));
    InMux I__1526 (
            .O(N__10241),
            .I(N__10226));
    InMux I__1525 (
            .O(N__10240),
            .I(N__10219));
    InMux I__1524 (
            .O(N__10239),
            .I(N__10216));
    InMux I__1523 (
            .O(N__10236),
            .I(N__10213));
    InMux I__1522 (
            .O(N__10235),
            .I(N__10208));
    InMux I__1521 (
            .O(N__10234),
            .I(N__10208));
    LocalMux I__1520 (
            .O(N__10231),
            .I(N__10203));
    LocalMux I__1519 (
            .O(N__10226),
            .I(N__10203));
    InMux I__1518 (
            .O(N__10225),
            .I(N__10196));
    InMux I__1517 (
            .O(N__10224),
            .I(N__10196));
    InMux I__1516 (
            .O(N__10223),
            .I(N__10196));
    InMux I__1515 (
            .O(N__10222),
            .I(N__10193));
    LocalMux I__1514 (
            .O(N__10219),
            .I(\this_vga_signals.mult1_un61_sum_axb3 ));
    LocalMux I__1513 (
            .O(N__10216),
            .I(\this_vga_signals.mult1_un61_sum_axb3 ));
    LocalMux I__1512 (
            .O(N__10213),
            .I(\this_vga_signals.mult1_un61_sum_axb3 ));
    LocalMux I__1511 (
            .O(N__10208),
            .I(\this_vga_signals.mult1_un61_sum_axb3 ));
    Odrv4 I__1510 (
            .O(N__10203),
            .I(\this_vga_signals.mult1_un61_sum_axb3 ));
    LocalMux I__1509 (
            .O(N__10196),
            .I(\this_vga_signals.mult1_un61_sum_axb3 ));
    LocalMux I__1508 (
            .O(N__10193),
            .I(\this_vga_signals.mult1_un61_sum_axb3 ));
    CascadeMux I__1507 (
            .O(N__10178),
            .I(\this_vga_signals.if_m4_0_1_0_cascade_ ));
    InMux I__1506 (
            .O(N__10175),
            .I(N__10169));
    InMux I__1505 (
            .O(N__10174),
            .I(N__10169));
    LocalMux I__1504 (
            .O(N__10169),
            .I(\this_vga_signals.mult1_un54_sum_axbxc5 ));
    CascadeMux I__1503 (
            .O(N__10166),
            .I(N__10162));
    InMux I__1502 (
            .O(N__10165),
            .I(N__10151));
    InMux I__1501 (
            .O(N__10162),
            .I(N__10151));
    InMux I__1500 (
            .O(N__10161),
            .I(N__10151));
    InMux I__1499 (
            .O(N__10160),
            .I(N__10144));
    InMux I__1498 (
            .O(N__10159),
            .I(N__10144));
    InMux I__1497 (
            .O(N__10158),
            .I(N__10137));
    LocalMux I__1496 (
            .O(N__10151),
            .I(N__10134));
    CascadeMux I__1495 (
            .O(N__10150),
            .I(N__10131));
    InMux I__1494 (
            .O(N__10149),
            .I(N__10125));
    LocalMux I__1493 (
            .O(N__10144),
            .I(N__10122));
    InMux I__1492 (
            .O(N__10143),
            .I(N__10117));
    InMux I__1491 (
            .O(N__10142),
            .I(N__10117));
    InMux I__1490 (
            .O(N__10141),
            .I(N__10112));
    InMux I__1489 (
            .O(N__10140),
            .I(N__10112));
    LocalMux I__1488 (
            .O(N__10137),
            .I(N__10107));
    Span4Mux_v I__1487 (
            .O(N__10134),
            .I(N__10107));
    InMux I__1486 (
            .O(N__10131),
            .I(N__10102));
    InMux I__1485 (
            .O(N__10130),
            .I(N__10102));
    InMux I__1484 (
            .O(N__10129),
            .I(N__10097));
    InMux I__1483 (
            .O(N__10128),
            .I(N__10097));
    LocalMux I__1482 (
            .O(N__10125),
            .I(\this_vga_signals.un12_address_cry_7_c_RNI32HB ));
    Odrv4 I__1481 (
            .O(N__10122),
            .I(\this_vga_signals.un12_address_cry_7_c_RNI32HB ));
    LocalMux I__1480 (
            .O(N__10117),
            .I(\this_vga_signals.un12_address_cry_7_c_RNI32HB ));
    LocalMux I__1479 (
            .O(N__10112),
            .I(\this_vga_signals.un12_address_cry_7_c_RNI32HB ));
    Odrv4 I__1478 (
            .O(N__10107),
            .I(\this_vga_signals.un12_address_cry_7_c_RNI32HB ));
    LocalMux I__1477 (
            .O(N__10102),
            .I(\this_vga_signals.un12_address_cry_7_c_RNI32HB ));
    LocalMux I__1476 (
            .O(N__10097),
            .I(\this_vga_signals.un12_address_cry_7_c_RNI32HB ));
    CascadeMux I__1475 (
            .O(N__10082),
            .I(N__10079));
    InMux I__1474 (
            .O(N__10079),
            .I(N__10076));
    LocalMux I__1473 (
            .O(N__10076),
            .I(\this_vga_signals.if_m2_3_0 ));
    InMux I__1472 (
            .O(N__10073),
            .I(N__10070));
    LocalMux I__1471 (
            .O(N__10070),
            .I(\this_vga_signals.mult1_un61_sum_axb3_1 ));
    InMux I__1470 (
            .O(N__10067),
            .I(N__10064));
    LocalMux I__1469 (
            .O(N__10064),
            .I(\this_vga_signals.G_12_0_3_1 ));
    CascadeMux I__1468 (
            .O(N__10061),
            .I(\this_vga_signals.N_9_cascade_ ));
    CascadeMux I__1467 (
            .O(N__10058),
            .I(N__10055));
    InMux I__1466 (
            .O(N__10055),
            .I(N__10052));
    LocalMux I__1465 (
            .O(N__10052),
            .I(\this_vga_signals.g1_1 ));
    CascadeMux I__1464 (
            .O(N__10049),
            .I(\this_vga_signals.mult1_un61_sum_axb3_0_cascade_ ));
    CascadeMux I__1463 (
            .O(N__10046),
            .I(\this_vga_signals.g0_4_0_1_cascade_ ));
    InMux I__1462 (
            .O(N__10043),
            .I(N__10039));
    InMux I__1461 (
            .O(N__10042),
            .I(N__10036));
    LocalMux I__1460 (
            .O(N__10039),
            .I(N__10033));
    LocalMux I__1459 (
            .O(N__10036),
            .I(\this_vga_signals.g1_1_0 ));
    Odrv4 I__1458 (
            .O(N__10033),
            .I(\this_vga_signals.g1_1_0 ));
    InMux I__1457 (
            .O(N__10028),
            .I(N__10016));
    InMux I__1456 (
            .O(N__10027),
            .I(N__10016));
    InMux I__1455 (
            .O(N__10026),
            .I(N__10016));
    InMux I__1454 (
            .O(N__10025),
            .I(N__10013));
    InMux I__1453 (
            .O(N__10024),
            .I(N__10006));
    InMux I__1452 (
            .O(N__10023),
            .I(N__10006));
    LocalMux I__1451 (
            .O(N__10016),
            .I(N__10003));
    LocalMux I__1450 (
            .O(N__10013),
            .I(N__9992));
    InMux I__1449 (
            .O(N__10012),
            .I(N__9987));
    InMux I__1448 (
            .O(N__10011),
            .I(N__9987));
    LocalMux I__1447 (
            .O(N__10006),
            .I(N__9982));
    Span4Mux_v I__1446 (
            .O(N__10003),
            .I(N__9982));
    InMux I__1445 (
            .O(N__10002),
            .I(N__9977));
    InMux I__1444 (
            .O(N__10001),
            .I(N__9977));
    InMux I__1443 (
            .O(N__10000),
            .I(N__9968));
    InMux I__1442 (
            .O(N__9999),
            .I(N__9968));
    InMux I__1441 (
            .O(N__9998),
            .I(N__9968));
    InMux I__1440 (
            .O(N__9997),
            .I(N__9968));
    InMux I__1439 (
            .O(N__9996),
            .I(N__9963));
    InMux I__1438 (
            .O(N__9995),
            .I(N__9963));
    Odrv12 I__1437 (
            .O(N__9992),
            .I(\this_vga_signals.mult1_un54_sum_axb3_out ));
    LocalMux I__1436 (
            .O(N__9987),
            .I(\this_vga_signals.mult1_un54_sum_axb3_out ));
    Odrv4 I__1435 (
            .O(N__9982),
            .I(\this_vga_signals.mult1_un54_sum_axb3_out ));
    LocalMux I__1434 (
            .O(N__9977),
            .I(\this_vga_signals.mult1_un54_sum_axb3_out ));
    LocalMux I__1433 (
            .O(N__9968),
            .I(\this_vga_signals.mult1_un54_sum_axb3_out ));
    LocalMux I__1432 (
            .O(N__9963),
            .I(\this_vga_signals.mult1_un54_sum_axb3_out ));
    InMux I__1431 (
            .O(N__9950),
            .I(N__9947));
    LocalMux I__1430 (
            .O(N__9947),
            .I(N__9941));
    InMux I__1429 (
            .O(N__9946),
            .I(N__9938));
    InMux I__1428 (
            .O(N__9945),
            .I(N__9933));
    InMux I__1427 (
            .O(N__9944),
            .I(N__9933));
    Odrv4 I__1426 (
            .O(N__9941),
            .I(\this_vga_signals.mult1_un54_sum_axb4 ));
    LocalMux I__1425 (
            .O(N__9938),
            .I(\this_vga_signals.mult1_un54_sum_axb4 ));
    LocalMux I__1424 (
            .O(N__9933),
            .I(\this_vga_signals.mult1_un54_sum_axb4 ));
    CascadeMux I__1423 (
            .O(N__9926),
            .I(N__9922));
    InMux I__1422 (
            .O(N__9925),
            .I(N__9915));
    InMux I__1421 (
            .O(N__9922),
            .I(N__9912));
    InMux I__1420 (
            .O(N__9921),
            .I(N__9907));
    InMux I__1419 (
            .O(N__9920),
            .I(N__9907));
    InMux I__1418 (
            .O(N__9919),
            .I(N__9902));
    InMux I__1417 (
            .O(N__9918),
            .I(N__9902));
    LocalMux I__1416 (
            .O(N__9915),
            .I(\this_vga_signals.mult1_un47_sum_c5 ));
    LocalMux I__1415 (
            .O(N__9912),
            .I(\this_vga_signals.mult1_un47_sum_c5 ));
    LocalMux I__1414 (
            .O(N__9907),
            .I(\this_vga_signals.mult1_un47_sum_c5 ));
    LocalMux I__1413 (
            .O(N__9902),
            .I(\this_vga_signals.mult1_un47_sum_c5 ));
    InMux I__1412 (
            .O(N__9893),
            .I(N__9890));
    LocalMux I__1411 (
            .O(N__9890),
            .I(\this_vga_signals.mult1_un61_sum_axb4_x0 ));
    CascadeMux I__1410 (
            .O(N__9887),
            .I(\this_vga_signals.mult1_un54_sum_ac0_7_cascade_ ));
    InMux I__1409 (
            .O(N__9884),
            .I(N__9881));
    LocalMux I__1408 (
            .O(N__9881),
            .I(\this_vga_signals.mult1_un61_sum_axb4_x1 ));
    CascadeMux I__1407 (
            .O(N__9878),
            .I(\this_vga_signals.mult1_un61_sum_axb4_i_cascade_ ));
    CascadeMux I__1406 (
            .O(N__9875),
            .I(\this_vga_signals.mult1_un61_sum_ac0_5_cascade_ ));
    InMux I__1405 (
            .O(N__9872),
            .I(N__9869));
    LocalMux I__1404 (
            .O(N__9869),
            .I(\this_vga_signals.mult1_un61_sum_axb4_i ));
    InMux I__1403 (
            .O(N__9866),
            .I(N__9863));
    LocalMux I__1402 (
            .O(N__9863),
            .I(N__9859));
    InMux I__1401 (
            .O(N__9862),
            .I(N__9856));
    Span4Mux_h I__1400 (
            .O(N__9859),
            .I(N__9853));
    LocalMux I__1399 (
            .O(N__9856),
            .I(N__9850));
    Odrv4 I__1398 (
            .O(N__9853),
            .I(\this_vga_signals.M_vcounter_q_RNITV8S_2Z0Z_0 ));
    Odrv4 I__1397 (
            .O(N__9850),
            .I(\this_vga_signals.M_vcounter_q_RNITV8S_2Z0Z_0 ));
    CascadeMux I__1396 (
            .O(N__9845),
            .I(\this_vga_signals.M_vcounter_q_RNI8OSG6BZ0Z_2_cascade_ ));
    InMux I__1395 (
            .O(N__9842),
            .I(N__9836));
    InMux I__1394 (
            .O(N__9841),
            .I(N__9836));
    LocalMux I__1393 (
            .O(N__9836),
            .I(\this_vga_signals.mult1_un61_sum_axb1_0 ));
    InMux I__1392 (
            .O(N__9833),
            .I(N__9826));
    InMux I__1391 (
            .O(N__9832),
            .I(N__9826));
    InMux I__1390 (
            .O(N__9831),
            .I(N__9817));
    LocalMux I__1389 (
            .O(N__9826),
            .I(N__9814));
    InMux I__1388 (
            .O(N__9825),
            .I(N__9811));
    InMux I__1387 (
            .O(N__9824),
            .I(N__9806));
    InMux I__1386 (
            .O(N__9823),
            .I(N__9806));
    InMux I__1385 (
            .O(N__9822),
            .I(N__9799));
    InMux I__1384 (
            .O(N__9821),
            .I(N__9799));
    InMux I__1383 (
            .O(N__9820),
            .I(N__9799));
    LocalMux I__1382 (
            .O(N__9817),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    Odrv4 I__1381 (
            .O(N__9814),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    LocalMux I__1380 (
            .O(N__9811),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    LocalMux I__1379 (
            .O(N__9806),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    LocalMux I__1378 (
            .O(N__9799),
            .I(\this_vga_signals.mult1_un54_sum_c3 ));
    InMux I__1377 (
            .O(N__9788),
            .I(N__9785));
    LocalMux I__1376 (
            .O(N__9785),
            .I(\this_vga_signals.address_m35_1 ));
    InMux I__1375 (
            .O(N__9782),
            .I(N__9776));
    InMux I__1374 (
            .O(N__9781),
            .I(N__9773));
    InMux I__1373 (
            .O(N__9780),
            .I(N__9770));
    InMux I__1372 (
            .O(N__9779),
            .I(N__9767));
    LocalMux I__1371 (
            .O(N__9776),
            .I(N__9760));
    LocalMux I__1370 (
            .O(N__9773),
            .I(N__9757));
    LocalMux I__1369 (
            .O(N__9770),
            .I(N__9752));
    LocalMux I__1368 (
            .O(N__9767),
            .I(N__9752));
    InMux I__1367 (
            .O(N__9766),
            .I(N__9747));
    InMux I__1366 (
            .O(N__9765),
            .I(N__9747));
    InMux I__1365 (
            .O(N__9764),
            .I(N__9742));
    InMux I__1364 (
            .O(N__9763),
            .I(N__9742));
    Odrv4 I__1363 (
            .O(N__9760),
            .I(\this_vga_signals.N_75_mux ));
    Odrv4 I__1362 (
            .O(N__9757),
            .I(\this_vga_signals.N_75_mux ));
    Odrv4 I__1361 (
            .O(N__9752),
            .I(\this_vga_signals.N_75_mux ));
    LocalMux I__1360 (
            .O(N__9747),
            .I(\this_vga_signals.N_75_mux ));
    LocalMux I__1359 (
            .O(N__9742),
            .I(\this_vga_signals.N_75_mux ));
    CascadeMux I__1358 (
            .O(N__9731),
            .I(N__9728));
    InMux I__1357 (
            .O(N__9728),
            .I(N__9721));
    InMux I__1356 (
            .O(N__9727),
            .I(N__9716));
    InMux I__1355 (
            .O(N__9726),
            .I(N__9716));
    CascadeMux I__1354 (
            .O(N__9725),
            .I(N__9713));
    CascadeMux I__1353 (
            .O(N__9724),
            .I(N__9710));
    LocalMux I__1352 (
            .O(N__9721),
            .I(N__9706));
    LocalMux I__1351 (
            .O(N__9716),
            .I(N__9703));
    InMux I__1350 (
            .O(N__9713),
            .I(N__9700));
    InMux I__1349 (
            .O(N__9710),
            .I(N__9697));
    CascadeMux I__1348 (
            .O(N__9709),
            .I(N__9694));
    Span4Mux_v I__1347 (
            .O(N__9706),
            .I(N__9689));
    Span4Mux_v I__1346 (
            .O(N__9703),
            .I(N__9689));
    LocalMux I__1345 (
            .O(N__9700),
            .I(N__9686));
    LocalMux I__1344 (
            .O(N__9697),
            .I(N__9683));
    InMux I__1343 (
            .O(N__9694),
            .I(N__9680));
    Sp12to4 I__1342 (
            .O(N__9689),
            .I(N__9677));
    Span4Mux_h I__1341 (
            .O(N__9686),
            .I(N__9674));
    Sp12to4 I__1340 (
            .O(N__9683),
            .I(N__9669));
    LocalMux I__1339 (
            .O(N__9680),
            .I(N__9669));
    Odrv12 I__1338 (
            .O(N__9677),
            .I(\this_vga_signals.N_84 ));
    Odrv4 I__1337 (
            .O(N__9674),
            .I(\this_vga_signals.N_84 ));
    Odrv12 I__1336 (
            .O(N__9669),
            .I(\this_vga_signals.N_84 ));
    InMux I__1335 (
            .O(N__9662),
            .I(N__9659));
    LocalMux I__1334 (
            .O(N__9659),
            .I(N__9656));
    Span4Mux_h I__1333 (
            .O(N__9656),
            .I(N__9653));
    Odrv4 I__1332 (
            .O(N__9653),
            .I(\this_vga_signals.M_vcounter_q_RNO_0Z0Z_2 ));
    CascadeMux I__1331 (
            .O(N__9650),
            .I(N__9647));
    InMux I__1330 (
            .O(N__9647),
            .I(N__9644));
    LocalMux I__1329 (
            .O(N__9644),
            .I(\this_vga_signals.address_m31_1 ));
    InMux I__1328 (
            .O(N__9641),
            .I(N__9638));
    LocalMux I__1327 (
            .O(N__9638),
            .I(\this_vga_signals.address_i2_mux_4 ));
    CascadeMux I__1326 (
            .O(N__9635),
            .I(N__9630));
    InMux I__1325 (
            .O(N__9634),
            .I(N__9627));
    InMux I__1324 (
            .O(N__9633),
            .I(N__9622));
    InMux I__1323 (
            .O(N__9630),
            .I(N__9622));
    LocalMux I__1322 (
            .O(N__9627),
            .I(\this_vga_signals.M_vcounter_q_RNITV8S_1Z0Z_0 ));
    LocalMux I__1321 (
            .O(N__9622),
            .I(\this_vga_signals.M_vcounter_q_RNITV8S_1Z0Z_0 ));
    InMux I__1320 (
            .O(N__9617),
            .I(N__9614));
    LocalMux I__1319 (
            .O(N__9614),
            .I(\this_vga_signals.address_N_9_0 ));
    CascadeMux I__1318 (
            .O(N__9611),
            .I(\this_vga_signals.address_N_33_cascade_ ));
    InMux I__1317 (
            .O(N__9608),
            .I(N__9605));
    LocalMux I__1316 (
            .O(N__9605),
            .I(\this_vga_signals.address_N_34 ));
    InMux I__1315 (
            .O(N__9602),
            .I(N__9586));
    InMux I__1314 (
            .O(N__9601),
            .I(N__9586));
    InMux I__1313 (
            .O(N__9600),
            .I(N__9586));
    InMux I__1312 (
            .O(N__9599),
            .I(N__9586));
    InMux I__1311 (
            .O(N__9598),
            .I(N__9586));
    InMux I__1310 (
            .O(N__9597),
            .I(N__9583));
    LocalMux I__1309 (
            .O(N__9586),
            .I(\this_vga_signals.M_vstate_qZ0Z_1 ));
    LocalMux I__1308 (
            .O(N__9583),
            .I(\this_vga_signals.M_vstate_qZ0Z_1 ));
    CascadeMux I__1307 (
            .O(N__9578),
            .I(\this_vga_signals.m35_e_1_cascade_ ));
    InMux I__1306 (
            .O(N__9575),
            .I(N__9572));
    LocalMux I__1305 (
            .O(N__9572),
            .I(N__9568));
    InMux I__1304 (
            .O(N__9571),
            .I(N__9565));
    Odrv4 I__1303 (
            .O(N__9568),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_0 ));
    LocalMux I__1302 (
            .O(N__9565),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_0 ));
    InMux I__1301 (
            .O(N__9560),
            .I(N__9557));
    LocalMux I__1300 (
            .O(N__9557),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1 ));
    CascadeMux I__1299 (
            .O(N__9554),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1_cascade_ ));
    CascadeMux I__1298 (
            .O(N__9551),
            .I(N__9547));
    InMux I__1297 (
            .O(N__9550),
            .I(N__9544));
    InMux I__1296 (
            .O(N__9547),
            .I(N__9541));
    LocalMux I__1295 (
            .O(N__9544),
            .I(\this_vga_signals.mult1_un68_sum_c2 ));
    LocalMux I__1294 (
            .O(N__9541),
            .I(\this_vga_signals.mult1_un68_sum_c2 ));
    CascadeMux I__1293 (
            .O(N__9536),
            .I(\this_vga_signals.address_N_9_0_cascade_ ));
    InMux I__1292 (
            .O(N__9533),
            .I(N__9530));
    LocalMux I__1291 (
            .O(N__9530),
            .I(\this_vga_signals.address_N_10_0 ));
    InMux I__1290 (
            .O(N__9527),
            .I(N__9523));
    InMux I__1289 (
            .O(N__9526),
            .I(N__9520));
    LocalMux I__1288 (
            .O(N__9523),
            .I(\this_vga_signals.address_N_3 ));
    LocalMux I__1287 (
            .O(N__9520),
            .I(\this_vga_signals.address_N_3 ));
    IoInMux I__1286 (
            .O(N__9515),
            .I(N__9512));
    LocalMux I__1285 (
            .O(N__9512),
            .I(N__9509));
    IoSpan4Mux I__1284 (
            .O(N__9509),
            .I(N__9506));
    IoSpan4Mux I__1283 (
            .O(N__9506),
            .I(N__9503));
    Span4Mux_s3_v I__1282 (
            .O(N__9503),
            .I(N__9500));
    Span4Mux_v I__1281 (
            .O(N__9500),
            .I(N__9497));
    Span4Mux_v I__1280 (
            .O(N__9497),
            .I(N__9494));
    Odrv4 I__1279 (
            .O(N__9494),
            .I(vsync_c));
    CascadeMux I__1278 (
            .O(N__9491),
            .I(\this_vga_signals.N_52_cascade_ ));
    InMux I__1277 (
            .O(N__9488),
            .I(N__9485));
    LocalMux I__1276 (
            .O(N__9485),
            .I(\this_vga_signals.N_76_mux ));
    CascadeMux I__1275 (
            .O(N__9482),
            .I(\this_vga_signals.N_76_mux_cascade_ ));
    InMux I__1274 (
            .O(N__9479),
            .I(N__9473));
    InMux I__1273 (
            .O(N__9478),
            .I(N__9473));
    LocalMux I__1272 (
            .O(N__9473),
            .I(\this_vga_signals.N_72_mux ));
    CascadeMux I__1271 (
            .O(N__9470),
            .I(\this_vga_signals.N_55_cascade_ ));
    CascadeMux I__1270 (
            .O(N__9467),
            .I(\this_vga_signals.M_vstate_q_RNO_1Z0Z_0_cascade_ ));
    InMux I__1269 (
            .O(N__9464),
            .I(N__9461));
    LocalMux I__1268 (
            .O(N__9461),
            .I(\this_vga_signals.M_vstate_q_RNO_2Z0Z_0 ));
    InMux I__1267 (
            .O(N__9458),
            .I(N__9455));
    LocalMux I__1266 (
            .O(N__9455),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_3 ));
    CascadeMux I__1265 (
            .O(N__9452),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ));
    InMux I__1264 (
            .O(N__9449),
            .I(N__9446));
    LocalMux I__1263 (
            .O(N__9446),
            .I(\this_vga_signals.mult1_un54_sum_c4 ));
    CascadeMux I__1262 (
            .O(N__9443),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_4_cascade_ ));
    CascadeMux I__1261 (
            .O(N__9440),
            .I(\this_vga_signals.if_m4_0_1_cascade_ ));
    CascadeMux I__1260 (
            .O(N__9437),
            .I(\this_vga_signals.G_12_0_x3_0_cascade_ ));
    CascadeMux I__1259 (
            .O(N__9434),
            .I(N__9430));
    CascadeMux I__1258 (
            .O(N__9433),
            .I(N__9425));
    InMux I__1257 (
            .O(N__9430),
            .I(N__9417));
    InMux I__1256 (
            .O(N__9429),
            .I(N__9417));
    InMux I__1255 (
            .O(N__9428),
            .I(N__9408));
    InMux I__1254 (
            .O(N__9425),
            .I(N__9408));
    InMux I__1253 (
            .O(N__9424),
            .I(N__9408));
    InMux I__1252 (
            .O(N__9423),
            .I(N__9408));
    InMux I__1251 (
            .O(N__9422),
            .I(N__9405));
    LocalMux I__1250 (
            .O(N__9417),
            .I(\this_vga_signals.un12_address_cry_10_c_RNINP5K ));
    LocalMux I__1249 (
            .O(N__9408),
            .I(\this_vga_signals.un12_address_cry_10_c_RNINP5K ));
    LocalMux I__1248 (
            .O(N__9405),
            .I(\this_vga_signals.un12_address_cry_10_c_RNINP5K ));
    CascadeMux I__1247 (
            .O(N__9398),
            .I(\this_vga_signals.un12_address_cry_9_c_RNIVF1R_cascade_ ));
    CascadeMux I__1246 (
            .O(N__9395),
            .I(N__9387));
    CascadeMux I__1245 (
            .O(N__9394),
            .I(N__9384));
    InMux I__1244 (
            .O(N__9393),
            .I(N__9378));
    InMux I__1243 (
            .O(N__9392),
            .I(N__9378));
    InMux I__1242 (
            .O(N__9391),
            .I(N__9369));
    InMux I__1241 (
            .O(N__9390),
            .I(N__9369));
    InMux I__1240 (
            .O(N__9387),
            .I(N__9369));
    InMux I__1239 (
            .O(N__9384),
            .I(N__9369));
    InMux I__1238 (
            .O(N__9383),
            .I(N__9366));
    LocalMux I__1237 (
            .O(N__9378),
            .I(\this_vga_signals.un12_address_cry_9_c_RNIEJOE ));
    LocalMux I__1236 (
            .O(N__9369),
            .I(\this_vga_signals.un12_address_cry_9_c_RNIEJOE ));
    LocalMux I__1235 (
            .O(N__9366),
            .I(\this_vga_signals.un12_address_cry_9_c_RNIEJOE ));
    CascadeMux I__1234 (
            .O(N__9359),
            .I(\this_vga_signals.mult1_un47_sum_c5_cascade_ ));
    CascadeMux I__1233 (
            .O(N__9356),
            .I(\this_vga_signals.mult1_un61_sum_axb3_x1_cascade_ ));
    CascadeMux I__1232 (
            .O(N__9353),
            .I(\this_vga_signals.mult1_un61_sum_axb3_cascade_ ));
    InMux I__1231 (
            .O(N__9350),
            .I(N__9347));
    LocalMux I__1230 (
            .O(N__9347),
            .I(\this_vga_signals.if_m5_sn ));
    CascadeMux I__1229 (
            .O(N__9344),
            .I(\this_vga_signals.if_m5_rn_0_cascade_ ));
    CascadeMux I__1228 (
            .O(N__9341),
            .I(\this_vga_signals.mult1_un68_sum_c5_cascade_ ));
    CascadeMux I__1227 (
            .O(N__9338),
            .I(N__9335));
    CascadeBuf I__1226 (
            .O(N__9335),
            .I(N__9332));
    CascadeMux I__1225 (
            .O(N__9332),
            .I(N__9329));
    CascadeBuf I__1224 (
            .O(N__9329),
            .I(N__9326));
    CascadeMux I__1223 (
            .O(N__9326),
            .I(N__9323));
    CascadeBuf I__1222 (
            .O(N__9323),
            .I(N__9320));
    CascadeMux I__1221 (
            .O(N__9320),
            .I(N__9317));
    CascadeBuf I__1220 (
            .O(N__9317),
            .I(N__9314));
    CascadeMux I__1219 (
            .O(N__9314),
            .I(N__9311));
    CascadeBuf I__1218 (
            .O(N__9311),
            .I(N__9308));
    CascadeMux I__1217 (
            .O(N__9308),
            .I(N__9305));
    CascadeBuf I__1216 (
            .O(N__9305),
            .I(N__9302));
    CascadeMux I__1215 (
            .O(N__9302),
            .I(N__9299));
    CascadeBuf I__1214 (
            .O(N__9299),
            .I(N__9296));
    CascadeMux I__1213 (
            .O(N__9296),
            .I(N__9293));
    CascadeBuf I__1212 (
            .O(N__9293),
            .I(N__9290));
    CascadeMux I__1211 (
            .O(N__9290),
            .I(N__9287));
    CascadeBuf I__1210 (
            .O(N__9287),
            .I(N__9284));
    CascadeMux I__1209 (
            .O(N__9284),
            .I(N__9281));
    CascadeBuf I__1208 (
            .O(N__9281),
            .I(N__9278));
    CascadeMux I__1207 (
            .O(N__9278),
            .I(N__9275));
    CascadeBuf I__1206 (
            .O(N__9275),
            .I(N__9272));
    CascadeMux I__1205 (
            .O(N__9272),
            .I(N__9269));
    CascadeBuf I__1204 (
            .O(N__9269),
            .I(N__9266));
    CascadeMux I__1203 (
            .O(N__9266),
            .I(N__9263));
    CascadeBuf I__1202 (
            .O(N__9263),
            .I(N__9260));
    CascadeMux I__1201 (
            .O(N__9260),
            .I(N__9257));
    CascadeBuf I__1200 (
            .O(N__9257),
            .I(N__9254));
    CascadeMux I__1199 (
            .O(N__9254),
            .I(N__9251));
    CascadeBuf I__1198 (
            .O(N__9251),
            .I(N__9248));
    CascadeMux I__1197 (
            .O(N__9248),
            .I(N__9245));
    InMux I__1196 (
            .O(N__9245),
            .I(N__9242));
    LocalMux I__1195 (
            .O(N__9242),
            .I(N__9239));
    Span12Mux_h I__1194 (
            .O(N__9239),
            .I(N__9236));
    Span12Mux_v I__1193 (
            .O(N__9236),
            .I(N__9233));
    Odrv12 I__1192 (
            .O(N__9233),
            .I(M_this_vga_signals_address_4));
    CascadeMux I__1191 (
            .O(N__9230),
            .I(\this_vga_signals.mult1_un54_sum_ac0_8_cascade_ ));
    InMux I__1190 (
            .O(N__9227),
            .I(N__9224));
    LocalMux I__1189 (
            .O(N__9224),
            .I(\this_vga_signals.g1_1_1 ));
    InMux I__1188 (
            .O(N__9221),
            .I(N__9217));
    InMux I__1187 (
            .O(N__9220),
            .I(N__9211));
    LocalMux I__1186 (
            .O(N__9217),
            .I(N__9206));
    InMux I__1185 (
            .O(N__9216),
            .I(N__9201));
    InMux I__1184 (
            .O(N__9215),
            .I(N__9201));
    InMux I__1183 (
            .O(N__9214),
            .I(N__9197));
    LocalMux I__1182 (
            .O(N__9211),
            .I(N__9194));
    InMux I__1181 (
            .O(N__9210),
            .I(N__9189));
    InMux I__1180 (
            .O(N__9209),
            .I(N__9189));
    Span4Mux_h I__1179 (
            .O(N__9206),
            .I(N__9184));
    LocalMux I__1178 (
            .O(N__9201),
            .I(N__9184));
    InMux I__1177 (
            .O(N__9200),
            .I(N__9181));
    LocalMux I__1176 (
            .O(N__9197),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    Odrv4 I__1175 (
            .O(N__9194),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    LocalMux I__1174 (
            .O(N__9189),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    Odrv4 I__1173 (
            .O(N__9184),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    LocalMux I__1172 (
            .O(N__9181),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    InMux I__1171 (
            .O(N__9170),
            .I(N__9166));
    InMux I__1170 (
            .O(N__9169),
            .I(N__9163));
    LocalMux I__1169 (
            .O(N__9166),
            .I(N__9158));
    LocalMux I__1168 (
            .O(N__9163),
            .I(N__9158));
    Odrv12 I__1167 (
            .O(N__9158),
            .I(\this_vga_signals.M_hcounter_q_i_11 ));
    InMux I__1166 (
            .O(N__9155),
            .I(N__9149));
    InMux I__1165 (
            .O(N__9154),
            .I(N__9149));
    LocalMux I__1164 (
            .O(N__9149),
            .I(\this_vga_signals.un12_address_cry_9_THRU_CO ));
    InMux I__1163 (
            .O(N__9146),
            .I(N__9136));
    InMux I__1162 (
            .O(N__9145),
            .I(N__9136));
    InMux I__1161 (
            .O(N__9144),
            .I(N__9127));
    InMux I__1160 (
            .O(N__9143),
            .I(N__9127));
    InMux I__1159 (
            .O(N__9142),
            .I(N__9127));
    InMux I__1158 (
            .O(N__9141),
            .I(N__9127));
    LocalMux I__1157 (
            .O(N__9136),
            .I(\this_vga_signals.un12_address_cry_9_c_RNIVF1R ));
    LocalMux I__1156 (
            .O(N__9127),
            .I(\this_vga_signals.un12_address_cry_9_c_RNIVF1R ));
    CascadeMux I__1155 (
            .O(N__9122),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_cascade_ ));
    CascadeMux I__1154 (
            .O(N__9119),
            .I(N__9114));
    InMux I__1153 (
            .O(N__9118),
            .I(N__9108));
    InMux I__1152 (
            .O(N__9117),
            .I(N__9108));
    InMux I__1151 (
            .O(N__9114),
            .I(N__9103));
    InMux I__1150 (
            .O(N__9113),
            .I(N__9103));
    LocalMux I__1149 (
            .O(N__9108),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    LocalMux I__1148 (
            .O(N__9103),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    InMux I__1147 (
            .O(N__9098),
            .I(N__9092));
    InMux I__1146 (
            .O(N__9097),
            .I(N__9092));
    LocalMux I__1145 (
            .O(N__9092),
            .I(\this_vga_signals.mult1_un61_sum_c2 ));
    CascadeMux I__1144 (
            .O(N__9089),
            .I(N__9086));
    InMux I__1143 (
            .O(N__9086),
            .I(N__9083));
    LocalMux I__1142 (
            .O(N__9083),
            .I(\this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2 ));
    InMux I__1141 (
            .O(N__9080),
            .I(N__9077));
    LocalMux I__1140 (
            .O(N__9077),
            .I(\this_vga_signals.address_i3_mux_i ));
    CascadeMux I__1139 (
            .O(N__9074),
            .I(\this_vga_signals.address_m27_ns_1_cascade_ ));
    CascadeMux I__1138 (
            .O(N__9071),
            .I(\this_vga_signals.address_i2_mux_3_cascade_ ));
    InMux I__1137 (
            .O(N__9068),
            .I(N__9065));
    LocalMux I__1136 (
            .O(N__9065),
            .I(\this_vga_signals.address_i2_mux_2 ));
    InMux I__1135 (
            .O(N__9062),
            .I(N__9059));
    LocalMux I__1134 (
            .O(N__9059),
            .I(N__9056));
    Span4Mux_h I__1133 (
            .O(N__9056),
            .I(N__9053));
    Odrv4 I__1132 (
            .O(N__9053),
            .I(\this_vga_signals.M_vcounter_q_RNO_0Z0Z_1 ));
    IoInMux I__1131 (
            .O(N__9050),
            .I(N__9047));
    LocalMux I__1130 (
            .O(N__9047),
            .I(N__9044));
    Span4Mux_s3_h I__1129 (
            .O(N__9044),
            .I(N__9041));
    Span4Mux_v I__1128 (
            .O(N__9041),
            .I(N__9037));
    IoInMux I__1127 (
            .O(N__9040),
            .I(N__9034));
    Span4Mux_v I__1126 (
            .O(N__9037),
            .I(N__9031));
    LocalMux I__1125 (
            .O(N__9034),
            .I(N__9028));
    Span4Mux_v I__1124 (
            .O(N__9031),
            .I(N__9023));
    Span4Mux_s3_h I__1123 (
            .O(N__9028),
            .I(N__9023));
    Span4Mux_v I__1122 (
            .O(N__9023),
            .I(N__9020));
    Span4Mux_h I__1121 (
            .O(N__9020),
            .I(N__9017));
    Odrv4 I__1120 (
            .O(N__9017),
            .I(rgb_c_0));
    InMux I__1119 (
            .O(N__9014),
            .I(N__9009));
    CascadeMux I__1118 (
            .O(N__9013),
            .I(N__9004));
    InMux I__1117 (
            .O(N__9012),
            .I(N__8997));
    LocalMux I__1116 (
            .O(N__9009),
            .I(N__8993));
    InMux I__1115 (
            .O(N__9008),
            .I(N__8988));
    InMux I__1114 (
            .O(N__9007),
            .I(N__8988));
    InMux I__1113 (
            .O(N__9004),
            .I(N__8985));
    CascadeMux I__1112 (
            .O(N__9003),
            .I(N__8982));
    InMux I__1111 (
            .O(N__9002),
            .I(N__8979));
    CascadeMux I__1110 (
            .O(N__9001),
            .I(N__8976));
    InMux I__1109 (
            .O(N__9000),
            .I(N__8973));
    LocalMux I__1108 (
            .O(N__8997),
            .I(N__8970));
    InMux I__1107 (
            .O(N__8996),
            .I(N__8967));
    Span4Mux_v I__1106 (
            .O(N__8993),
            .I(N__8962));
    LocalMux I__1105 (
            .O(N__8988),
            .I(N__8962));
    LocalMux I__1104 (
            .O(N__8985),
            .I(N__8959));
    InMux I__1103 (
            .O(N__8982),
            .I(N__8956));
    LocalMux I__1102 (
            .O(N__8979),
            .I(N__8953));
    InMux I__1101 (
            .O(N__8976),
            .I(N__8950));
    LocalMux I__1100 (
            .O(N__8973),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__1099 (
            .O(N__8970),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__1098 (
            .O(N__8967),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__1097 (
            .O(N__8962),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__1096 (
            .O(N__8959),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__1095 (
            .O(N__8956),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv12 I__1094 (
            .O(N__8953),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__1093 (
            .O(N__8950),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    InMux I__1092 (
            .O(N__8933),
            .I(N__8930));
    LocalMux I__1091 (
            .O(N__8930),
            .I(\this_vga_signals.address_m1_1_1 ));
    InMux I__1090 (
            .O(N__8927),
            .I(N__8923));
    InMux I__1089 (
            .O(N__8926),
            .I(N__8920));
    LocalMux I__1088 (
            .O(N__8923),
            .I(\this_vga_signals.mult1_un54_sum_c2 ));
    LocalMux I__1087 (
            .O(N__8920),
            .I(\this_vga_signals.mult1_un54_sum_c2 ));
    CascadeMux I__1086 (
            .O(N__8915),
            .I(\this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2_cascade_ ));
    CascadeMux I__1085 (
            .O(N__8912),
            .I(N__8909));
    InMux I__1084 (
            .O(N__8909),
            .I(N__8906));
    LocalMux I__1083 (
            .O(N__8906),
            .I(\this_vga_signals.mult1_un61_sum_c3_1 ));
    CascadeMux I__1082 (
            .O(N__8903),
            .I(\this_vga_signals.mult1_un61_sum_c3_cascade_ ));
    InMux I__1081 (
            .O(N__8900),
            .I(N__8890));
    InMux I__1080 (
            .O(N__8899),
            .I(N__8885));
    InMux I__1079 (
            .O(N__8898),
            .I(N__8885));
    InMux I__1078 (
            .O(N__8897),
            .I(N__8874));
    InMux I__1077 (
            .O(N__8896),
            .I(N__8874));
    InMux I__1076 (
            .O(N__8895),
            .I(N__8874));
    InMux I__1075 (
            .O(N__8894),
            .I(N__8874));
    InMux I__1074 (
            .O(N__8893),
            .I(N__8874));
    LocalMux I__1073 (
            .O(N__8890),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1072 (
            .O(N__8885),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1071 (
            .O(N__8874),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    InMux I__1070 (
            .O(N__8867),
            .I(N__8861));
    InMux I__1069 (
            .O(N__8866),
            .I(N__8861));
    LocalMux I__1068 (
            .O(N__8861),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_0 ));
    InMux I__1067 (
            .O(N__8858),
            .I(N__8855));
    LocalMux I__1066 (
            .O(N__8855),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_3_2 ));
    InMux I__1065 (
            .O(N__8852),
            .I(N__8848));
    InMux I__1064 (
            .O(N__8851),
            .I(N__8843));
    LocalMux I__1063 (
            .O(N__8848),
            .I(N__8840));
    InMux I__1062 (
            .O(N__8847),
            .I(N__8837));
    CascadeMux I__1061 (
            .O(N__8846),
            .I(N__8833));
    LocalMux I__1060 (
            .O(N__8843),
            .I(N__8825));
    Span4Mux_v I__1059 (
            .O(N__8840),
            .I(N__8825));
    LocalMux I__1058 (
            .O(N__8837),
            .I(N__8825));
    InMux I__1057 (
            .O(N__8836),
            .I(N__8822));
    InMux I__1056 (
            .O(N__8833),
            .I(N__8819));
    InMux I__1055 (
            .O(N__8832),
            .I(N__8816));
    Span4Mux_h I__1054 (
            .O(N__8825),
            .I(N__8813));
    LocalMux I__1053 (
            .O(N__8822),
            .I(N__8808));
    LocalMux I__1052 (
            .O(N__8819),
            .I(N__8808));
    LocalMux I__1051 (
            .O(N__8816),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__1050 (
            .O(N__8813),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv12 I__1049 (
            .O(N__8808),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    InMux I__1048 (
            .O(N__8801),
            .I(N__8797));
    CascadeMux I__1047 (
            .O(N__8800),
            .I(N__8794));
    LocalMux I__1046 (
            .O(N__8797),
            .I(N__8791));
    InMux I__1045 (
            .O(N__8794),
            .I(N__8788));
    Span4Mux_h I__1044 (
            .O(N__8791),
            .I(N__8785));
    LocalMux I__1043 (
            .O(N__8788),
            .I(N__8782));
    Odrv4 I__1042 (
            .O(N__8785),
            .I(\this_vga_signals.N_27 ));
    Odrv4 I__1041 (
            .O(N__8782),
            .I(\this_vga_signals.N_27 ));
    CascadeMux I__1040 (
            .O(N__8777),
            .I(N__8770));
    InMux I__1039 (
            .O(N__8776),
            .I(N__8765));
    InMux I__1038 (
            .O(N__8775),
            .I(N__8765));
    InMux I__1037 (
            .O(N__8774),
            .I(N__8762));
    InMux I__1036 (
            .O(N__8773),
            .I(N__8759));
    InMux I__1035 (
            .O(N__8770),
            .I(N__8756));
    LocalMux I__1034 (
            .O(N__8765),
            .I(N__8752));
    LocalMux I__1033 (
            .O(N__8762),
            .I(N__8749));
    LocalMux I__1032 (
            .O(N__8759),
            .I(N__8746));
    LocalMux I__1031 (
            .O(N__8756),
            .I(N__8743));
    InMux I__1030 (
            .O(N__8755),
            .I(N__8740));
    Span4Mux_h I__1029 (
            .O(N__8752),
            .I(N__8737));
    Span4Mux_v I__1028 (
            .O(N__8749),
            .I(N__8730));
    Span4Mux_v I__1027 (
            .O(N__8746),
            .I(N__8730));
    Span4Mux_v I__1026 (
            .O(N__8743),
            .I(N__8730));
    LocalMux I__1025 (
            .O(N__8740),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1024 (
            .O(N__8737),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1023 (
            .O(N__8730),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    InMux I__1022 (
            .O(N__8723),
            .I(N__8720));
    LocalMux I__1021 (
            .O(N__8720),
            .I(N__8717));
    Odrv4 I__1020 (
            .O(N__8717),
            .I(\this_vga_signals.hvisible_i_a2_2_0 ));
    IoInMux I__1019 (
            .O(N__8714),
            .I(N__8711));
    LocalMux I__1018 (
            .O(N__8711),
            .I(N__8708));
    Span4Mux_s2_h I__1017 (
            .O(N__8708),
            .I(N__8704));
    IoInMux I__1016 (
            .O(N__8707),
            .I(N__8701));
    Span4Mux_h I__1015 (
            .O(N__8704),
            .I(N__8698));
    LocalMux I__1014 (
            .O(N__8701),
            .I(N__8695));
    Span4Mux_h I__1013 (
            .O(N__8698),
            .I(N__8692));
    Span12Mux_s10_h I__1012 (
            .O(N__8695),
            .I(N__8689));
    Span4Mux_v I__1011 (
            .O(N__8692),
            .I(N__8686));
    Odrv12 I__1010 (
            .O(N__8689),
            .I(rgb_c_4));
    Odrv4 I__1009 (
            .O(N__8686),
            .I(rgb_c_4));
    InMux I__1008 (
            .O(N__8681),
            .I(N__8678));
    LocalMux I__1007 (
            .O(N__8678),
            .I(\this_vga_signals.m30_3 ));
    CascadeMux I__1006 (
            .O(N__8675),
            .I(\this_vga_signals.m30_4_cascade_ ));
    InMux I__1005 (
            .O(N__8672),
            .I(N__8667));
    InMux I__1004 (
            .O(N__8671),
            .I(N__8661));
    InMux I__1003 (
            .O(N__8670),
            .I(N__8658));
    LocalMux I__1002 (
            .O(N__8667),
            .I(N__8655));
    CascadeMux I__1001 (
            .O(N__8666),
            .I(N__8652));
    CascadeMux I__1000 (
            .O(N__8665),
            .I(N__8649));
    CascadeMux I__999 (
            .O(N__8664),
            .I(N__8643));
    LocalMux I__998 (
            .O(N__8661),
            .I(N__8639));
    LocalMux I__997 (
            .O(N__8658),
            .I(N__8636));
    Span4Mux_h I__996 (
            .O(N__8655),
            .I(N__8633));
    InMux I__995 (
            .O(N__8652),
            .I(N__8630));
    InMux I__994 (
            .O(N__8649),
            .I(N__8625));
    InMux I__993 (
            .O(N__8648),
            .I(N__8625));
    InMux I__992 (
            .O(N__8647),
            .I(N__8622));
    InMux I__991 (
            .O(N__8646),
            .I(N__8617));
    InMux I__990 (
            .O(N__8643),
            .I(N__8617));
    InMux I__989 (
            .O(N__8642),
            .I(N__8614));
    Odrv4 I__988 (
            .O(N__8639),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__987 (
            .O(N__8636),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__986 (
            .O(N__8633),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__985 (
            .O(N__8630),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__984 (
            .O(N__8625),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__983 (
            .O(N__8622),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__982 (
            .O(N__8617),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__981 (
            .O(N__8614),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    InMux I__980 (
            .O(N__8597),
            .I(N__8593));
    CascadeMux I__979 (
            .O(N__8596),
            .I(N__8584));
    LocalMux I__978 (
            .O(N__8593),
            .I(N__8580));
    InMux I__977 (
            .O(N__8592),
            .I(N__8577));
    InMux I__976 (
            .O(N__8591),
            .I(N__8574));
    InMux I__975 (
            .O(N__8590),
            .I(N__8571));
    InMux I__974 (
            .O(N__8589),
            .I(N__8568));
    InMux I__973 (
            .O(N__8588),
            .I(N__8565));
    InMux I__972 (
            .O(N__8587),
            .I(N__8558));
    InMux I__971 (
            .O(N__8584),
            .I(N__8558));
    InMux I__970 (
            .O(N__8583),
            .I(N__8558));
    Span4Mux_v I__969 (
            .O(N__8580),
            .I(N__8553));
    LocalMux I__968 (
            .O(N__8577),
            .I(N__8553));
    LocalMux I__967 (
            .O(N__8574),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__966 (
            .O(N__8571),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__965 (
            .O(N__8568),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__964 (
            .O(N__8565),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__963 (
            .O(N__8558),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__962 (
            .O(N__8553),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    InMux I__961 (
            .O(N__8540),
            .I(N__8535));
    InMux I__960 (
            .O(N__8539),
            .I(N__8532));
    InMux I__959 (
            .O(N__8538),
            .I(N__8526));
    LocalMux I__958 (
            .O(N__8535),
            .I(N__8518));
    LocalMux I__957 (
            .O(N__8532),
            .I(N__8515));
    InMux I__956 (
            .O(N__8531),
            .I(N__8508));
    InMux I__955 (
            .O(N__8530),
            .I(N__8505));
    InMux I__954 (
            .O(N__8529),
            .I(N__8502));
    LocalMux I__953 (
            .O(N__8526),
            .I(N__8499));
    InMux I__952 (
            .O(N__8525),
            .I(N__8494));
    InMux I__951 (
            .O(N__8524),
            .I(N__8494));
    InMux I__950 (
            .O(N__8523),
            .I(N__8489));
    InMux I__949 (
            .O(N__8522),
            .I(N__8489));
    InMux I__948 (
            .O(N__8521),
            .I(N__8486));
    Span4Mux_h I__947 (
            .O(N__8518),
            .I(N__8483));
    Span4Mux_h I__946 (
            .O(N__8515),
            .I(N__8480));
    InMux I__945 (
            .O(N__8514),
            .I(N__8477));
    InMux I__944 (
            .O(N__8513),
            .I(N__8470));
    InMux I__943 (
            .O(N__8512),
            .I(N__8470));
    InMux I__942 (
            .O(N__8511),
            .I(N__8470));
    LocalMux I__941 (
            .O(N__8508),
            .I(N__8465));
    LocalMux I__940 (
            .O(N__8505),
            .I(N__8465));
    LocalMux I__939 (
            .O(N__8502),
            .I(N__8462));
    Span4Mux_h I__938 (
            .O(N__8499),
            .I(N__8455));
    LocalMux I__937 (
            .O(N__8494),
            .I(N__8455));
    LocalMux I__936 (
            .O(N__8489),
            .I(N__8455));
    LocalMux I__935 (
            .O(N__8486),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__934 (
            .O(N__8483),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__933 (
            .O(N__8480),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__932 (
            .O(N__8477),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__931 (
            .O(N__8470),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__930 (
            .O(N__8465),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv12 I__929 (
            .O(N__8462),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__928 (
            .O(N__8455),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    CascadeMux I__927 (
            .O(N__8438),
            .I(\this_vga_signals.N_3_0_cascade_ ));
    InMux I__926 (
            .O(N__8435),
            .I(N__8430));
    CascadeMux I__925 (
            .O(N__8434),
            .I(N__8421));
    CascadeMux I__924 (
            .O(N__8433),
            .I(N__8418));
    LocalMux I__923 (
            .O(N__8430),
            .I(N__8415));
    InMux I__922 (
            .O(N__8429),
            .I(N__8412));
    InMux I__921 (
            .O(N__8428),
            .I(N__8409));
    InMux I__920 (
            .O(N__8427),
            .I(N__8404));
    InMux I__919 (
            .O(N__8426),
            .I(N__8404));
    InMux I__918 (
            .O(N__8425),
            .I(N__8401));
    InMux I__917 (
            .O(N__8424),
            .I(N__8398));
    InMux I__916 (
            .O(N__8421),
            .I(N__8393));
    InMux I__915 (
            .O(N__8418),
            .I(N__8393));
    Odrv4 I__914 (
            .O(N__8415),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__913 (
            .O(N__8412),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__912 (
            .O(N__8409),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__911 (
            .O(N__8404),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__910 (
            .O(N__8401),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__909 (
            .O(N__8398),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__908 (
            .O(N__8393),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    InMux I__907 (
            .O(N__8378),
            .I(\this_vga_signals.un12_address_cry_10 ));
    InMux I__906 (
            .O(N__8375),
            .I(N__8372));
    LocalMux I__905 (
            .O(N__8372),
            .I(N__8367));
    CascadeMux I__904 (
            .O(N__8371),
            .I(N__8364));
    InMux I__903 (
            .O(N__8370),
            .I(N__8361));
    Span4Mux_v I__902 (
            .O(N__8367),
            .I(N__8358));
    InMux I__901 (
            .O(N__8364),
            .I(N__8355));
    LocalMux I__900 (
            .O(N__8361),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__899 (
            .O(N__8358),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__898 (
            .O(N__8355),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    InMux I__897 (
            .O(N__8348),
            .I(N__8345));
    LocalMux I__896 (
            .O(N__8345),
            .I(N__8341));
    InMux I__895 (
            .O(N__8344),
            .I(N__8338));
    Span4Mux_h I__894 (
            .O(N__8341),
            .I(N__8335));
    LocalMux I__893 (
            .O(N__8338),
            .I(\this_vga_signals.N_49 ));
    Odrv4 I__892 (
            .O(N__8335),
            .I(\this_vga_signals.N_49 ));
    CascadeMux I__891 (
            .O(N__8330),
            .I(N__8325));
    InMux I__890 (
            .O(N__8329),
            .I(N__8320));
    InMux I__889 (
            .O(N__8328),
            .I(N__8317));
    InMux I__888 (
            .O(N__8325),
            .I(N__8314));
    InMux I__887 (
            .O(N__8324),
            .I(N__8309));
    InMux I__886 (
            .O(N__8323),
            .I(N__8309));
    LocalMux I__885 (
            .O(N__8320),
            .I(\this_vga_signals.M_hcounter_qZ0Z_11 ));
    LocalMux I__884 (
            .O(N__8317),
            .I(\this_vga_signals.M_hcounter_qZ0Z_11 ));
    LocalMux I__883 (
            .O(N__8314),
            .I(\this_vga_signals.M_hcounter_qZ0Z_11 ));
    LocalMux I__882 (
            .O(N__8309),
            .I(\this_vga_signals.M_hcounter_qZ0Z_11 ));
    IoInMux I__881 (
            .O(N__8300),
            .I(N__8297));
    LocalMux I__880 (
            .O(N__8297),
            .I(N__8294));
    Span4Mux_s3_v I__879 (
            .O(N__8294),
            .I(N__8291));
    Span4Mux_h I__878 (
            .O(N__8291),
            .I(N__8287));
    InMux I__877 (
            .O(N__8290),
            .I(N__8284));
    Sp12to4 I__876 (
            .O(N__8287),
            .I(N__8281));
    LocalMux I__875 (
            .O(N__8284),
            .I(N__8278));
    Span12Mux_v I__874 (
            .O(N__8281),
            .I(N__8274));
    Span12Mux_s10_h I__873 (
            .O(N__8278),
            .I(N__8271));
    InMux I__872 (
            .O(N__8277),
            .I(N__8268));
    Odrv12 I__871 (
            .O(N__8274),
            .I(N_16));
    Odrv12 I__870 (
            .O(N__8271),
            .I(N_16));
    LocalMux I__869 (
            .O(N__8268),
            .I(N_16));
    CascadeMux I__868 (
            .O(N__8261),
            .I(\this_vga_signals.mult1_un61_sum_ac0_7_0_3_1_1_cascade_ ));
    CascadeMux I__867 (
            .O(N__8258),
            .I(N__8253));
    InMux I__866 (
            .O(N__8257),
            .I(N__8250));
    InMux I__865 (
            .O(N__8256),
            .I(N__8247));
    InMux I__864 (
            .O(N__8253),
            .I(N__8244));
    LocalMux I__863 (
            .O(N__8250),
            .I(N__8241));
    LocalMux I__862 (
            .O(N__8247),
            .I(N__8236));
    LocalMux I__861 (
            .O(N__8244),
            .I(N__8236));
    Span4Mux_h I__860 (
            .O(N__8241),
            .I(N__8233));
    Span4Mux_v I__859 (
            .O(N__8236),
            .I(N__8230));
    Odrv4 I__858 (
            .O(N__8233),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__857 (
            .O(N__8230),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__856 (
            .O(N__8225),
            .I(\this_vga_signals.un12_address_cry_1 ));
    CascadeMux I__855 (
            .O(N__8222),
            .I(N__8219));
    InMux I__854 (
            .O(N__8219),
            .I(N__8214));
    InMux I__853 (
            .O(N__8218),
            .I(N__8211));
    InMux I__852 (
            .O(N__8217),
            .I(N__8208));
    LocalMux I__851 (
            .O(N__8214),
            .I(N__8205));
    LocalMux I__850 (
            .O(N__8211),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__849 (
            .O(N__8208),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__848 (
            .O(N__8205),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__847 (
            .O(N__8198),
            .I(\this_vga_signals.un12_address_cry_2 ));
    CascadeMux I__846 (
            .O(N__8195),
            .I(N__8190));
    InMux I__845 (
            .O(N__8194),
            .I(N__8187));
    InMux I__844 (
            .O(N__8193),
            .I(N__8184));
    InMux I__843 (
            .O(N__8190),
            .I(N__8181));
    LocalMux I__842 (
            .O(N__8187),
            .I(N__8178));
    LocalMux I__841 (
            .O(N__8184),
            .I(N__8173));
    LocalMux I__840 (
            .O(N__8181),
            .I(N__8173));
    Span4Mux_h I__839 (
            .O(N__8178),
            .I(N__8170));
    Span4Mux_h I__838 (
            .O(N__8173),
            .I(N__8167));
    Odrv4 I__837 (
            .O(N__8170),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__836 (
            .O(N__8167),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__835 (
            .O(N__8162),
            .I(\this_vga_signals.un12_address_cry_3 ));
    CascadeMux I__834 (
            .O(N__8159),
            .I(N__8155));
    CascadeMux I__833 (
            .O(N__8158),
            .I(N__8151));
    InMux I__832 (
            .O(N__8155),
            .I(N__8148));
    InMux I__831 (
            .O(N__8154),
            .I(N__8145));
    InMux I__830 (
            .O(N__8151),
            .I(N__8142));
    LocalMux I__829 (
            .O(N__8148),
            .I(N__8139));
    LocalMux I__828 (
            .O(N__8145),
            .I(N__8134));
    LocalMux I__827 (
            .O(N__8142),
            .I(N__8134));
    Span4Mux_h I__826 (
            .O(N__8139),
            .I(N__8131));
    Span4Mux_h I__825 (
            .O(N__8134),
            .I(N__8128));
    Odrv4 I__824 (
            .O(N__8131),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__823 (
            .O(N__8128),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    InMux I__822 (
            .O(N__8123),
            .I(\this_vga_signals.un12_address_cry_4 ));
    InMux I__821 (
            .O(N__8120),
            .I(\this_vga_signals.un12_address_cry_5 ));
    InMux I__820 (
            .O(N__8117),
            .I(N__8111));
    CascadeMux I__819 (
            .O(N__8116),
            .I(N__8108));
    InMux I__818 (
            .O(N__8115),
            .I(N__8103));
    InMux I__817 (
            .O(N__8114),
            .I(N__8103));
    LocalMux I__816 (
            .O(N__8111),
            .I(N__8100));
    InMux I__815 (
            .O(N__8108),
            .I(N__8097));
    LocalMux I__814 (
            .O(N__8103),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__813 (
            .O(N__8100),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__812 (
            .O(N__8097),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__811 (
            .O(N__8090),
            .I(\this_vga_signals.un12_address_cry_6 ));
    InMux I__810 (
            .O(N__8087),
            .I(bfn_11_18_0_));
    InMux I__809 (
            .O(N__8084),
            .I(\this_vga_signals.un12_address_cry_8 ));
    InMux I__808 (
            .O(N__8081),
            .I(\this_vga_signals.un12_address_cry_9 ));
    CascadeMux I__807 (
            .O(N__8078),
            .I(\this_vga_signals.address_m24_ns_1Z0Z_0_cascade_ ));
    InMux I__806 (
            .O(N__8075),
            .I(N__8072));
    LocalMux I__805 (
            .O(N__8072),
            .I(N__8068));
    InMux I__804 (
            .O(N__8071),
            .I(N__8060));
    Span4Mux_v I__803 (
            .O(N__8068),
            .I(N__8057));
    InMux I__802 (
            .O(N__8067),
            .I(N__8054));
    InMux I__801 (
            .O(N__8066),
            .I(N__8049));
    InMux I__800 (
            .O(N__8065),
            .I(N__8049));
    InMux I__799 (
            .O(N__8064),
            .I(N__8044));
    InMux I__798 (
            .O(N__8063),
            .I(N__8044));
    LocalMux I__797 (
            .O(N__8060),
            .I(N__8041));
    Odrv4 I__796 (
            .O(N__8057),
            .I(\this_vga_signals.mult1_un40_sum_c3 ));
    LocalMux I__795 (
            .O(N__8054),
            .I(\this_vga_signals.mult1_un40_sum_c3 ));
    LocalMux I__794 (
            .O(N__8049),
            .I(\this_vga_signals.mult1_un40_sum_c3 ));
    LocalMux I__793 (
            .O(N__8044),
            .I(\this_vga_signals.mult1_un40_sum_c3 ));
    Odrv4 I__792 (
            .O(N__8041),
            .I(\this_vga_signals.mult1_un40_sum_c3 ));
    CascadeMux I__791 (
            .O(N__8030),
            .I(\this_vga_signals.mult1_un54_sum_c2_cascade_ ));
    CascadeMux I__790 (
            .O(N__8027),
            .I(N__8024));
    InMux I__789 (
            .O(N__8024),
            .I(N__8017));
    InMux I__788 (
            .O(N__8023),
            .I(N__8017));
    InMux I__787 (
            .O(N__8022),
            .I(N__8014));
    LocalMux I__786 (
            .O(N__8017),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    LocalMux I__785 (
            .O(N__8014),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    CascadeMux I__784 (
            .O(N__8009),
            .I(\this_vga_signals.mult1_un54_sum_c3_cascade_ ));
    InMux I__783 (
            .O(N__8006),
            .I(N__8003));
    LocalMux I__782 (
            .O(N__8003),
            .I(\this_vga_signals.M_vcounter_q_RNO_0Z0Z_0 ));
    CascadeMux I__781 (
            .O(N__8000),
            .I(N__7995));
    InMux I__780 (
            .O(N__7999),
            .I(N__7991));
    InMux I__779 (
            .O(N__7998),
            .I(N__7988));
    InMux I__778 (
            .O(N__7995),
            .I(N__7985));
    InMux I__777 (
            .O(N__7994),
            .I(N__7982));
    LocalMux I__776 (
            .O(N__7991),
            .I(N__7975));
    LocalMux I__775 (
            .O(N__7988),
            .I(N__7975));
    LocalMux I__774 (
            .O(N__7985),
            .I(N__7975));
    LocalMux I__773 (
            .O(N__7982),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    Odrv4 I__772 (
            .O(N__7975),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    InMux I__771 (
            .O(N__7970),
            .I(N__7966));
    CascadeMux I__770 (
            .O(N__7969),
            .I(N__7962));
    LocalMux I__769 (
            .O(N__7966),
            .I(N__7959));
    CascadeMux I__768 (
            .O(N__7965),
            .I(N__7956));
    InMux I__767 (
            .O(N__7962),
            .I(N__7953));
    Span4Mux_h I__766 (
            .O(N__7959),
            .I(N__7950));
    InMux I__765 (
            .O(N__7956),
            .I(N__7947));
    LocalMux I__764 (
            .O(N__7953),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__763 (
            .O(N__7950),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__762 (
            .O(N__7947),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    InMux I__761 (
            .O(N__7940),
            .I(\this_vga_signals.un12_address_cry_0 ));
    InMux I__760 (
            .O(N__7937),
            .I(N__7931));
    InMux I__759 (
            .O(N__7936),
            .I(N__7924));
    InMux I__758 (
            .O(N__7935),
            .I(N__7924));
    InMux I__757 (
            .O(N__7934),
            .I(N__7924));
    LocalMux I__756 (
            .O(N__7931),
            .I(N__7919));
    LocalMux I__755 (
            .O(N__7924),
            .I(N__7916));
    InMux I__754 (
            .O(N__7923),
            .I(N__7911));
    InMux I__753 (
            .O(N__7922),
            .I(N__7911));
    Odrv4 I__752 (
            .O(N__7919),
            .I(\this_vga_signals.N_70 ));
    Odrv4 I__751 (
            .O(N__7916),
            .I(\this_vga_signals.N_70 ));
    LocalMux I__750 (
            .O(N__7911),
            .I(\this_vga_signals.N_70 ));
    InMux I__749 (
            .O(N__7904),
            .I(N__7900));
    InMux I__748 (
            .O(N__7903),
            .I(N__7897));
    LocalMux I__747 (
            .O(N__7900),
            .I(\this_vga_signals.SUM_0 ));
    LocalMux I__746 (
            .O(N__7897),
            .I(\this_vga_signals.SUM_0 ));
    InMux I__745 (
            .O(N__7892),
            .I(N__7889));
    LocalMux I__744 (
            .O(N__7889),
            .I(\this_vga_signals.mult1_un40_sum_axbxc1 ));
    InMux I__743 (
            .O(N__7886),
            .I(N__7883));
    LocalMux I__742 (
            .O(N__7883),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_c ));
    CascadeMux I__741 (
            .O(N__7880),
            .I(\this_vga_signals.mult1_un40_sum_axbxc1_cascade_ ));
    InMux I__740 (
            .O(N__7877),
            .I(N__7873));
    InMux I__739 (
            .O(N__7876),
            .I(N__7870));
    LocalMux I__738 (
            .O(N__7873),
            .I(\this_vga_signals.mult1_un47_sum_ac0_1 ));
    LocalMux I__737 (
            .O(N__7870),
            .I(\this_vga_signals.mult1_un47_sum_ac0_1 ));
    CascadeMux I__736 (
            .O(N__7865),
            .I(\this_vga_signals.mult1_un47_sum_c3_cascade_ ));
    CascadeMux I__735 (
            .O(N__7862),
            .I(N__7859));
    InMux I__734 (
            .O(N__7859),
            .I(N__7853));
    InMux I__733 (
            .O(N__7858),
            .I(N__7853));
    LocalMux I__732 (
            .O(N__7853),
            .I(N__7850));
    Odrv4 I__731 (
            .O(N__7850),
            .I(\this_vga_signals.N_13_0 ));
    InMux I__730 (
            .O(N__7847),
            .I(N__7841));
    InMux I__729 (
            .O(N__7846),
            .I(N__7841));
    LocalMux I__728 (
            .O(N__7841),
            .I(\this_vga_signals.if_i1_mux ));
    InMux I__727 (
            .O(N__7838),
            .I(N__7835));
    LocalMux I__726 (
            .O(N__7835),
            .I(N__7832));
    Odrv4 I__725 (
            .O(N__7832),
            .I(\this_vga_signals.M_vcounter_q_RNO_0Z0Z_3 ));
    CascadeMux I__724 (
            .O(N__7829),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_ ));
    CascadeMux I__723 (
            .O(N__7826),
            .I(\this_vga_signals.i9_mux_cascade_ ));
    InMux I__722 (
            .O(N__7823),
            .I(N__7820));
    LocalMux I__721 (
            .O(N__7820),
            .I(\this_vga_signals.i9_mux ));
    InMux I__720 (
            .O(N__7817),
            .I(N__7810));
    InMux I__719 (
            .O(N__7816),
            .I(N__7810));
    InMux I__718 (
            .O(N__7815),
            .I(N__7807));
    LocalMux I__717 (
            .O(N__7810),
            .I(\this_vga_signals.address_1_c5_i ));
    LocalMux I__716 (
            .O(N__7807),
            .I(\this_vga_signals.address_1_c5_i ));
    IoInMux I__715 (
            .O(N__7802),
            .I(N__7799));
    LocalMux I__714 (
            .O(N__7799),
            .I(N__7795));
    InMux I__713 (
            .O(N__7798),
            .I(N__7792));
    IoSpan4Mux I__712 (
            .O(N__7795),
            .I(N__7789));
    LocalMux I__711 (
            .O(N__7792),
            .I(N__7786));
    Span4Mux_s1_h I__710 (
            .O(N__7789),
            .I(N__7783));
    Span4Mux_v I__709 (
            .O(N__7786),
            .I(N__7779));
    Span4Mux_h I__708 (
            .O(N__7783),
            .I(N__7776));
    InMux I__707 (
            .O(N__7782),
            .I(N__7773));
    Span4Mux_h I__706 (
            .O(N__7779),
            .I(N__7770));
    Span4Mux_h I__705 (
            .O(N__7776),
            .I(N__7765));
    LocalMux I__704 (
            .O(N__7773),
            .I(N__7765));
    Span4Mux_v I__703 (
            .O(N__7770),
            .I(N__7760));
    Span4Mux_v I__702 (
            .O(N__7765),
            .I(N__7760));
    Odrv4 I__701 (
            .O(N__7760),
            .I(port_nmib_c));
    InMux I__700 (
            .O(N__7757),
            .I(N__7752));
    InMux I__699 (
            .O(N__7756),
            .I(N__7747));
    InMux I__698 (
            .O(N__7755),
            .I(N__7747));
    LocalMux I__697 (
            .O(N__7752),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    LocalMux I__696 (
            .O(N__7747),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    InMux I__695 (
            .O(N__7742),
            .I(N__7736));
    InMux I__694 (
            .O(N__7741),
            .I(N__7736));
    LocalMux I__693 (
            .O(N__7736),
            .I(N__7733));
    Odrv4 I__692 (
            .O(N__7733),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCNZ0 ));
    InMux I__691 (
            .O(N__7730),
            .I(N__7726));
    InMux I__690 (
            .O(N__7729),
            .I(N__7723));
    LocalMux I__689 (
            .O(N__7726),
            .I(N__7720));
    LocalMux I__688 (
            .O(N__7723),
            .I(N__7717));
    Span4Mux_h I__687 (
            .O(N__7720),
            .I(N__7714));
    Span4Mux_h I__686 (
            .O(N__7717),
            .I(N__7711));
    Odrv4 I__685 (
            .O(N__7714),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBNZ0 ));
    Odrv4 I__684 (
            .O(N__7711),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBNZ0 ));
    InMux I__683 (
            .O(N__7706),
            .I(N__7700));
    InMux I__682 (
            .O(N__7705),
            .I(N__7695));
    InMux I__681 (
            .O(N__7704),
            .I(N__7695));
    InMux I__680 (
            .O(N__7703),
            .I(N__7692));
    LocalMux I__679 (
            .O(N__7700),
            .I(N__7689));
    LocalMux I__678 (
            .O(N__7695),
            .I(N__7684));
    LocalMux I__677 (
            .O(N__7692),
            .I(N__7684));
    Span4Mux_v I__676 (
            .O(N__7689),
            .I(N__7679));
    Span4Mux_v I__675 (
            .O(N__7684),
            .I(N__7679));
    Sp12to4 I__674 (
            .O(N__7679),
            .I(N__7676));
    Span12Mux_h I__673 (
            .O(N__7676),
            .I(N__7673));
    Span12Mux_v I__672 (
            .O(N__7673),
            .I(N__7670));
    Odrv12 I__671 (
            .O(N__7670),
            .I(rst_n_c));
    InMux I__670 (
            .O(N__7667),
            .I(N__7664));
    LocalMux I__669 (
            .O(N__7664),
            .I(N__7661));
    Odrv4 I__668 (
            .O(N__7661),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__667 (
            .O(N__7658),
            .I(N__7655));
    LocalMux I__666 (
            .O(N__7655),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    CascadeMux I__665 (
            .O(N__7652),
            .I(\this_vga_signals.address_1_c4_cascade_ ));
    InMux I__664 (
            .O(N__7649),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_9 ));
    CascadeMux I__663 (
            .O(N__7646),
            .I(N__7642));
    InMux I__662 (
            .O(N__7645),
            .I(N__7636));
    InMux I__661 (
            .O(N__7642),
            .I(N__7633));
    InMux I__660 (
            .O(N__7641),
            .I(N__7630));
    InMux I__659 (
            .O(N__7640),
            .I(N__7627));
    InMux I__658 (
            .O(N__7639),
            .I(N__7624));
    LocalMux I__657 (
            .O(N__7636),
            .I(N__7619));
    LocalMux I__656 (
            .O(N__7633),
            .I(N__7619));
    LocalMux I__655 (
            .O(N__7630),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    LocalMux I__654 (
            .O(N__7627),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    LocalMux I__653 (
            .O(N__7624),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    Odrv12 I__652 (
            .O(N__7619),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    InMux I__651 (
            .O(N__7610),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_10 ));
    CascadeMux I__650 (
            .O(N__7607),
            .I(\this_vga_signals.g1_0_0_a2_0_cascade_ ));
    CascadeMux I__649 (
            .O(N__7604),
            .I(\this_vga_signals.g0_11_1_cascade_ ));
    CascadeMux I__648 (
            .O(N__7601),
            .I(N__7598));
    InMux I__647 (
            .O(N__7598),
            .I(N__7592));
    InMux I__646 (
            .O(N__7597),
            .I(N__7592));
    LocalMux I__645 (
            .O(N__7592),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    InMux I__644 (
            .O(N__7589),
            .I(N__7586));
    LocalMux I__643 (
            .O(N__7586),
            .I(N__7582));
    InMux I__642 (
            .O(N__7585),
            .I(N__7579));
    Span4Mux_v I__641 (
            .O(N__7582),
            .I(N__7574));
    LocalMux I__640 (
            .O(N__7579),
            .I(N__7574));
    Odrv4 I__639 (
            .O(N__7574),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KANZ0 ));
    InMux I__638 (
            .O(N__7571),
            .I(N__7562));
    InMux I__637 (
            .O(N__7570),
            .I(N__7562));
    InMux I__636 (
            .O(N__7569),
            .I(N__7562));
    LocalMux I__635 (
            .O(N__7562),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    CascadeMux I__634 (
            .O(N__7559),
            .I(N__7556));
    InMux I__633 (
            .O(N__7556),
            .I(N__7553));
    LocalMux I__632 (
            .O(N__7553),
            .I(\this_vga_signals.N_2 ));
    InMux I__631 (
            .O(N__7550),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__630 (
            .O(N__7547),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_0 ));
    InMux I__629 (
            .O(N__7544),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_1 ));
    InMux I__628 (
            .O(N__7541),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_2 ));
    InMux I__627 (
            .O(N__7538),
            .I(N__7535));
    LocalMux I__626 (
            .O(N__7535),
            .I(N__7531));
    InMux I__625 (
            .O(N__7534),
            .I(N__7528));
    Odrv4 I__624 (
            .O(N__7531),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7NZ0 ));
    LocalMux I__623 (
            .O(N__7528),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7NZ0 ));
    InMux I__622 (
            .O(N__7523),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_3 ));
    InMux I__621 (
            .O(N__7520),
            .I(N__7517));
    LocalMux I__620 (
            .O(N__7517),
            .I(N__7513));
    InMux I__619 (
            .O(N__7516),
            .I(N__7510));
    Odrv4 I__618 (
            .O(N__7513),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8NZ0 ));
    LocalMux I__617 (
            .O(N__7510),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8NZ0 ));
    InMux I__616 (
            .O(N__7505),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_4 ));
    InMux I__615 (
            .O(N__7502),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_5 ));
    InMux I__614 (
            .O(N__7499),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_6 ));
    InMux I__613 (
            .O(N__7496),
            .I(bfn_9_24_0_));
    InMux I__612 (
            .O(N__7493),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_8 ));
    InMux I__611 (
            .O(N__7490),
            .I(N__7487));
    LocalMux I__610 (
            .O(N__7487),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1 ));
    CascadeMux I__609 (
            .O(N__7484),
            .I(\this_vga_signals.mult1_un40_sum_c3_cascade_ ));
    CascadeMux I__608 (
            .O(N__7481),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_ ));
    CascadeMux I__607 (
            .O(N__7478),
            .I(\this_vga_signals.mult1_un47_sum_ac0_2_cascade_ ));
    CascadeMux I__606 (
            .O(N__7475),
            .I(\this_vga_signals.N_2_cascade_ ));
    InMux I__605 (
            .O(N__7472),
            .I(N__7468));
    InMux I__604 (
            .O(N__7471),
            .I(N__7465));
    LocalMux I__603 (
            .O(N__7468),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__602 (
            .O(N__7465),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    CascadeMux I__601 (
            .O(N__7460),
            .I(\this_vga_signals.N_70_cascade_ ));
    InMux I__600 (
            .O(N__7457),
            .I(N__7454));
    LocalMux I__599 (
            .O(N__7454),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_1_0 ));
    InMux I__598 (
            .O(N__7451),
            .I(N__7445));
    InMux I__597 (
            .O(N__7450),
            .I(N__7445));
    LocalMux I__596 (
            .O(N__7445),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    InMux I__595 (
            .O(N__7442),
            .I(N__7439));
    LocalMux I__594 (
            .O(N__7439),
            .I(\this_vga_signals.m44_0_0 ));
    CascadeMux I__593 (
            .O(N__7436),
            .I(\this_vga_signals.M_vcounter_q_RNIQE2J1Z0Z_9_cascade_ ));
    InMux I__592 (
            .O(N__7433),
            .I(N__7430));
    LocalMux I__591 (
            .O(N__7430),
            .I(\this_vga_signals.M_vcounter_q_fast_RNI3BJLZ0Z_4 ));
    InMux I__590 (
            .O(N__7427),
            .I(N__7424));
    LocalMux I__589 (
            .O(N__7424),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__588 (
            .O(N__7421),
            .I(N__7417));
    InMux I__587 (
            .O(N__7420),
            .I(N__7414));
    LocalMux I__586 (
            .O(N__7417),
            .I(N__7411));
    LocalMux I__585 (
            .O(N__7414),
            .I(N__7408));
    Span4Mux_h I__584 (
            .O(N__7411),
            .I(N__7405));
    Span4Mux_h I__583 (
            .O(N__7408),
            .I(N__7402));
    Odrv4 I__582 (
            .O(N__7405),
            .I(\this_vga_signals.N_32 ));
    Odrv4 I__581 (
            .O(N__7402),
            .I(\this_vga_signals.N_32 ));
    InMux I__580 (
            .O(N__7397),
            .I(N__7392));
    InMux I__579 (
            .O(N__7396),
            .I(N__7389));
    InMux I__578 (
            .O(N__7395),
            .I(N__7385));
    LocalMux I__577 (
            .O(N__7392),
            .I(N__7382));
    LocalMux I__576 (
            .O(N__7389),
            .I(N__7379));
    InMux I__575 (
            .O(N__7388),
            .I(N__7376));
    LocalMux I__574 (
            .O(N__7385),
            .I(N__7373));
    Span4Mux_v I__573 (
            .O(N__7382),
            .I(N__7370));
    Odrv4 I__572 (
            .O(N__7379),
            .I(\this_vga_signals.M_hstate_qZ0Z_0 ));
    LocalMux I__571 (
            .O(N__7376),
            .I(\this_vga_signals.M_hstate_qZ0Z_0 ));
    Odrv4 I__570 (
            .O(N__7373),
            .I(\this_vga_signals.M_hstate_qZ0Z_0 ));
    Odrv4 I__569 (
            .O(N__7370),
            .I(\this_vga_signals.M_hstate_qZ0Z_0 ));
    CascadeMux I__568 (
            .O(N__7361),
            .I(N__7358));
    InMux I__567 (
            .O(N__7358),
            .I(N__7355));
    LocalMux I__566 (
            .O(N__7355),
            .I(\this_vga_signals.N_26 ));
    CascadeMux I__565 (
            .O(N__7352),
            .I(\this_vga_signals.N_26_cascade_ ));
    InMux I__564 (
            .O(N__7349),
            .I(N__7346));
    LocalMux I__563 (
            .O(N__7346),
            .I(N__7342));
    InMux I__562 (
            .O(N__7345),
            .I(N__7339));
    Span4Mux_v I__561 (
            .O(N__7342),
            .I(N__7336));
    LocalMux I__560 (
            .O(N__7339),
            .I(N__7333));
    Sp12to4 I__559 (
            .O(N__7336),
            .I(N__7329));
    Span4Mux_h I__558 (
            .O(N__7333),
            .I(N__7326));
    InMux I__557 (
            .O(N__7332),
            .I(N__7323));
    Odrv12 I__556 (
            .O(N__7329),
            .I(\this_vga_signals.N_51 ));
    Odrv4 I__555 (
            .O(N__7326),
            .I(\this_vga_signals.N_51 ));
    LocalMux I__554 (
            .O(N__7323),
            .I(\this_vga_signals.N_51 ));
    InMux I__553 (
            .O(N__7316),
            .I(N__7310));
    InMux I__552 (
            .O(N__7315),
            .I(N__7310));
    LocalMux I__551 (
            .O(N__7310),
            .I(N__7307));
    Span4Mux_h I__550 (
            .O(N__7307),
            .I(N__7304));
    Odrv4 I__549 (
            .O(N__7304),
            .I(\this_vga_signals.N_273 ));
    CascadeMux I__548 (
            .O(N__7301),
            .I(\this_vga_signals.N_18_cascade_ ));
    IoInMux I__547 (
            .O(N__7298),
            .I(N__7295));
    LocalMux I__546 (
            .O(N__7295),
            .I(N__7292));
    IoSpan4Mux I__545 (
            .O(N__7292),
            .I(N__7289));
    Span4Mux_s2_v I__544 (
            .O(N__7289),
            .I(N__7286));
    Span4Mux_v I__543 (
            .O(N__7286),
            .I(N__7283));
    Span4Mux_v I__542 (
            .O(N__7283),
            .I(N__7280));
    Odrv4 I__541 (
            .O(N__7280),
            .I(this_vga_signals_N_274_i));
    CascadeMux I__540 (
            .O(N__7277),
            .I(\this_vga_signals.hvisible_i_a2_0_3_0_cascade_ ));
    InMux I__539 (
            .O(N__7274),
            .I(N__7266));
    InMux I__538 (
            .O(N__7273),
            .I(N__7266));
    InMux I__537 (
            .O(N__7272),
            .I(N__7263));
    InMux I__536 (
            .O(N__7271),
            .I(N__7258));
    LocalMux I__535 (
            .O(N__7266),
            .I(N__7253));
    LocalMux I__534 (
            .O(N__7263),
            .I(N__7253));
    InMux I__533 (
            .O(N__7262),
            .I(N__7250));
    InMux I__532 (
            .O(N__7261),
            .I(N__7247));
    LocalMux I__531 (
            .O(N__7258),
            .I(N__7242));
    Span4Mux_h I__530 (
            .O(N__7253),
            .I(N__7242));
    LocalMux I__529 (
            .O(N__7250),
            .I(\this_vga_signals.M_hstate_qZ0Z_1 ));
    LocalMux I__528 (
            .O(N__7247),
            .I(\this_vga_signals.M_hstate_qZ0Z_1 ));
    Odrv4 I__527 (
            .O(N__7242),
            .I(\this_vga_signals.M_hstate_qZ0Z_1 ));
    CascadeMux I__526 (
            .O(N__7235),
            .I(\this_vga_signals.N_49_cascade_ ));
    CascadeMux I__525 (
            .O(N__7232),
            .I(\this_vga_signals.N_29_cascade_ ));
    CascadeMux I__524 (
            .O(N__7229),
            .I(\this_vga_signals.N_40_cascade_ ));
    InMux I__523 (
            .O(N__7226),
            .I(N__7223));
    LocalMux I__522 (
            .O(N__7223),
            .I(N__7220));
    Odrv4 I__521 (
            .O(N__7220),
            .I(\this_vga_signals.N_20 ));
    IoInMux I__520 (
            .O(N__7217),
            .I(N__7214));
    LocalMux I__519 (
            .O(N__7214),
            .I(port_rw_c_i));
    IoInMux I__518 (
            .O(N__7211),
            .I(N__7208));
    LocalMux I__517 (
            .O(N__7208),
            .I(N__7205));
    Odrv12 I__516 (
            .O(N__7205),
            .I(port_nmib_c_i));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\this_vga_signals.un12_address_cry_7 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_6_cry_7 ),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_19_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_23_0_));
    defparam IN_MUX_bfv_19_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_24_0_ (
            .carryinitin(un1_M_current_address_q_cry_7),
            .carryinitout(bfn_19_24_0_));
    ICE_GB \this_reset_cond.M_stage_q_RNI6VB7_3  (
            .USERSIGNALTOGLOBALBUFFER(N__17739),
            .GLOBALBUFFEROUTPUT(N_339_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam port_data_rw_obuf_RNO_LC_1_21_2.C_ON=1'b0;
    defparam port_data_rw_obuf_RNO_LC_1_21_2.SEQ_MODE=4'b0000;
    defparam port_data_rw_obuf_RNO_LC_1_21_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 port_data_rw_obuf_RNO_LC_1_21_2 (
            .in0(N__19705),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(port_rw_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIL6FA3_0_9_LC_5_30_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIL6FA3_0_9_LC_5_30_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIL6FA3_0_9_LC_5_30_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIL6FA3_0_9_LC_5_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7798),
            .lcout(port_nmib_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_6_LC_7_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_6_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_7_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13486),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17351),
            .ce(),
            .sr(N__15473));
    defparam \this_vga_signals.M_hstate_q_RNO_2_0_LC_7_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_2_0_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_2_0_LC_7_18_3 .LUT_INIT=16'b1110111001110111;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_2_0_LC_7_18_3  (
            .in0(N__7273),
            .in1(N__8832),
            .in2(_gnd_net_),
            .in3(N__8755),
            .lcout(),
            .ltout(\this_vga_signals.N_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_1_0_LC_7_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_1_0_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_1_0_LC_7_18_4 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_1_0_LC_7_18_4  (
            .in0(N__8801),
            .in1(N__7395),
            .in2(N__7232),
            .in3(N__9221),
            .lcout(),
            .ltout(\this_vga_signals.N_40_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_0_0_LC_7_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_0_0_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_0_0_LC_7_18_5 .LUT_INIT=16'b1111101111110001;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_0_0_LC_7_18_5  (
            .in0(N__7274),
            .in1(N__7420),
            .in2(N__7229),
            .in3(N__7345),
            .lcout(\this_vga_signals.N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_9_LC_7_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_9_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_9_LC_7_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_9_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10025),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17351),
            .ce(),
            .sr(N__15473));
    defparam \this_vga_signals.M_hcounter_q_2_LC_7_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_2_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_7_19_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__14012),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17357),
            .ce(),
            .sr(N__15471));
    defparam \this_vga_signals.M_hcounter_q_4_LC_7_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_4_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_7_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12977),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17357),
            .ce(),
            .sr(N__15471));
    defparam \this_vga_signals.M_hcounter_q_5_LC_7_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_5_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13762),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17357),
            .ce(),
            .sr(N__15471));
    defparam \this_vga_signals.M_hstate_q_0_LC_7_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_0_LC_7_20_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hstate_q_0_LC_7_20_0 .LUT_INIT=16'b0000011100000010;
    LogicCell40 \this_vga_signals.M_hstate_q_0_LC_7_20_0  (
            .in0(N__7315),
            .in1(N__7226),
            .in2(N__17737),
            .in3(N__7388),
            .lcout(\this_vga_signals.M_hstate_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17362),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_0_1_LC_7_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_0_1_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_0_1_LC_7_20_3 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_0_1_LC_7_20_3  (
            .in0(N__7421),
            .in1(N__7261),
            .in2(_gnd_net_),
            .in3(N__7349),
            .lcout(),
            .ltout(\this_vga_signals.N_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_1_LC_7_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_1_LC_7_20_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hstate_q_1_LC_7_20_4 .LUT_INIT=16'b0000000001001110;
    LogicCell40 \this_vga_signals.M_hstate_q_1_LC_7_20_4  (
            .in0(N__7316),
            .in1(N__7262),
            .in2(N__7301),
            .in3(N__17738),
            .lcout(\this_vga_signals.M_hstate_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17362),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNI1P4R_0_LC_7_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNI1P4R_0_LC_7_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNI1P4R_0_LC_7_22_7 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \this_vga_signals.M_hstate_q_RNI1P4R_0_LC_7_22_7  (
            .in0(N__7396),
            .in1(N__7271),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_N_274_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_13_LC_9_15_0 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_13_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_13_LC_9_15_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vram.mem_radreg_13_LC_9_15_0  (
            .in0(N__7782),
            .in1(N__8290),
            .in2(_gnd_net_),
            .in3(N__8075),
            .lcout(\this_vram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17323),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_3_LC_9_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_3_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_9_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14042),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17336),
            .ce(),
            .sr(N__15472));
    defparam \this_vga_signals.M_hcounter_q_0_LC_9_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_9_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7999),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17336),
            .ce(),
            .sr(N__15472));
    defparam \this_vga_signals.M_hcounter_q_RNI84D41_1_LC_9_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI84D41_1_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI84D41_1_LC_9_18_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI84D41_1_LC_9_18_0  (
            .in0(N__8194),
            .in1(N__8257),
            .in2(N__8159),
            .in3(N__7970),
            .lcout(),
            .ltout(\this_vga_signals.hvisible_i_a2_0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI9JJM1_0_LC_9_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI9JJM1_0_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI9JJM1_0_LC_9_18_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI9JJM1_0_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__8217),
            .in2(N__7277),
            .in3(N__7994),
            .lcout(\this_vga_signals.N_49 ),
            .ltout(\this_vga_signals.N_49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI5RNE4_11_LC_9_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI5RNE4_11_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI5RNE4_11_LC_9_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI5RNE4_11_LC_9_18_2  (
            .in0(N__7272),
            .in1(N__7332),
            .in2(N__7235),
            .in3(N__8324),
            .lcout(\this_vga_signals.M_hstate_d_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_9_18_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_9_18_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_9_18_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_9_18_4  (
            .in0(N__7703),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17340),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIHS8C_11_LC_9_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIHS8C_11_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIHS8C_11_LC_9_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIHS8C_11_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8323),
            .lcout(\this_vga_signals.M_hcounter_q_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_9_19_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_9_19_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_9_19_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__7706),
            .in2(_gnd_net_),
            .in3(N__7427),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17346),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIAU8U1_6_LC_9_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIAU8U1_6_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIAU8U1_6_LC_9_19_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIAU8U1_6_LC_9_19_2  (
            .in0(N__8776),
            .in1(N__9210),
            .in2(N__7361),
            .in3(N__8851),
            .lcout(\this_vga_signals.N_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNID7PV_0_LC_9_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNID7PV_0_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNID7PV_0_LC_9_19_4 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \this_vga_signals.M_hstate_q_RNID7PV_0_LC_9_19_4  (
            .in0(N__7397),
            .in1(N__8375),
            .in2(_gnd_net_),
            .in3(N__8117),
            .lcout(\this_vga_signals.N_26 ),
            .ltout(\this_vga_signals.N_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIAU8U1_0_6_LC_9_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIAU8U1_0_6_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIAU8U1_0_6_LC_9_19_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIAU8U1_0_6_LC_9_19_5  (
            .in0(N__9209),
            .in1(N__8847),
            .in2(N__7352),
            .in3(N__8775),
            .lcout(\this_vga_signals.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_9_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_9_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__8344),
            .in2(_gnd_net_),
            .in3(N__8328),
            .lcout(\this_vga_signals.N_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_5_LC_9_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_5_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_5_LC_9_20_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_5_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__15508),
            .in2(_gnd_net_),
            .in3(N__7520),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17352),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_1_1_0_LC_9_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_1_1_0_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_1_1_0_LC_9_20_3 .LUT_INIT=16'b0101000011110101;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_1_1_0_LC_9_20_3  (
            .in0(N__7570),
            .in1(_gnd_net_),
            .in2(N__7601),
            .in3(N__7755),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_RNI3JK8_8_LC_9_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_RNI3JK8_8_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_RNI3JK8_8_LC_9_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_RNI3JK8_8_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__7597),
            .in2(_gnd_net_),
            .in3(N__7569),
            .lcout(\this_vga_signals.N_2 ),
            .ltout(\this_vga_signals.N_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_RNI3BJL_4_LC_9_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_RNI3BJL_4_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_RNI3BJL_4_LC_9_20_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_RNI3BJL_4_LC_9_20_5  (
            .in0(N__7451),
            .in1(N__7756),
            .in2(N__7475),
            .in3(N__7472),
            .lcout(\this_vga_signals.M_vcounter_q_fast_RNI3BJLZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_RNITCK8_4_LC_9_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_RNITCK8_4_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_RNITCK8_4_LC_9_20_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_RNITCK8_4_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__7471),
            .in2(_gnd_net_),
            .in3(N__7450),
            .lcout(\this_vga_signals.N_70 ),
            .ltout(\this_vga_signals.N_70_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_RNI61891_7_LC_9_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_RNI61891_7_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_RNI61891_7_LC_9_20_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_RNI61891_7_LC_9_20_7  (
            .in0(N__7571),
            .in1(N__8592),
            .in2(N__7460),
            .in3(N__8529),
            .lcout(\this_vga_signals.address_1_c5_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_1_LC_9_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_1_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_1_LC_9_21_0 .LUT_INIT=16'b0010001001000000;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_1_LC_9_21_0  (
            .in0(N__8524),
            .in1(N__7457),
            .in2(N__8596),
            .in3(N__7923),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_RNIVBOE1_9_LC_9_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_RNIVBOE1_9_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_RNIVBOE1_9_LC_9_21_1 .LUT_INIT=16'b1100110001111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_RNIVBOE1_9_LC_9_21_1  (
            .in0(N__8523),
            .in1(N__8583),
            .in2(N__8664),
            .in3(N__7757),
            .lcout(\this_vga_signals.m44_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_4_LC_9_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_4_LC_9_21_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_4_LC_9_21_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_4_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__15507),
            .in2(_gnd_net_),
            .in3(N__7538),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17358),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_LC_9_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_LC_9_21_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_LC_9_21_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_LC_9_21_3  (
            .in0(N__7585),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17710),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17358),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQE2J1_9_LC_9_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQE2J1_9_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQE2J1_9_LC_9_21_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQE2J1_9_LC_9_21_4  (
            .in0(N__8642),
            .in1(N__8522),
            .in2(N__8433),
            .in3(N__7922),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_RNIQE2J1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_RNI27M05_4_LC_9_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_RNI27M05_4_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_RNI27M05_4_LC_9_21_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_RNI27M05_4_LC_9_21_5  (
            .in0(N__7442),
            .in1(N__7815),
            .in2(N__7436),
            .in3(N__7433),
            .lcout(\this_vga_signals.SUM_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_LC_9_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_LC_9_21_6 .LUT_INIT=16'b1111111101000010;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_LC_9_21_6  (
            .in0(N__8587),
            .in1(N__8646),
            .in2(N__8434),
            .in3(N__7490),
            .lcout(\this_vga_signals.mult1_un40_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_1_LC_9_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_1_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_1_LC_9_21_7 .LUT_INIT=16'b0110000000000110;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_1_LC_9_21_7  (
            .in0(N__10518),
            .in1(N__9002),
            .in2(N__7484),
            .in3(N__8525),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_9_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_9_22_0 .LUT_INIT=16'b0111011110011001;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_9_22_0  (
            .in0(N__8648),
            .in1(N__8424),
            .in2(_gnd_net_),
            .in3(N__8588),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_c_0_LC_9_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_c_0_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_c_0_LC_9_22_1 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_c_0_LC_9_22_1  (
            .in0(N__7935),
            .in1(_gnd_net_),
            .in2(N__7481),
            .in3(N__8512),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_LC_9_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_LC_9_22_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_LC_9_22_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_LC_9_22_3  (
            .in0(N__15506),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7516),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17363),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_2_LC_9_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_2_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_2_LC_9_22_4 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_2_LC_9_22_4  (
            .in0(N__8513),
            .in1(N__8065),
            .in2(_gnd_net_),
            .in3(N__7936),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_ac0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc3_1_0_LC_9_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc3_1_0_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc3_1_0_LC_9_22_5 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc3_1_0_LC_9_22_5  (
            .in0(N__8066),
            .in1(N__7892),
            .in2(N__7478),
            .in3(N__7877),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_m3_LC_9_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_m3_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_m3_LC_9_22_6 .LUT_INIT=16'b0111111000000110;
    LogicCell40 \this_vga_signals.un5_address_if_m3_LC_9_22_6  (
            .in0(N__8511),
            .in1(N__7934),
            .in2(N__8665),
            .in3(N__7903),
            .lcout(\this_vga_signals.if_i1_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_LC_9_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_LC_9_22_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_LC_9_22_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_LC_9_22_7  (
            .in0(N__15505),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7534),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17363),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNO_0_0_LC_9_23_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_RNO_0_0_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNO_0_0_LC_9_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNO_0_0_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__10813),
            .in2(N__7646),
            .in3(N__7645),
            .lcout(\this_vga_signals.M_vcounter_q_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNO_0_1_LC_9_23_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_RNO_0_1_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNO_0_1_LC_9_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNO_0_1_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__10922),
            .in2(_gnd_net_),
            .in3(N__7547),
            .lcout(\this_vga_signals.M_vcounter_q_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNO_0_2_LC_9_23_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_RNO_0_2_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNO_0_2_LC_9_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNO_0_2_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__11030),
            .in2(_gnd_net_),
            .in3(N__7544),
            .lcout(\this_vga_signals.M_vcounter_q_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNO_0_3_LC_9_23_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_RNO_0_3_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNO_0_3_LC_9_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNO_0_3_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__10734),
            .in2(_gnd_net_),
            .in3(N__7541),
            .lcout(\this_vga_signals.M_vcounter_q_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7N_LC_9_23_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7N_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7N_LC_9_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7N_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__10531),
            .in2(_gnd_net_),
            .in3(N__7523),
            .lcout(\this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7NZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8N_LC_9_23_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8N_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8N_LC_9_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8N_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__9000),
            .in2(_gnd_net_),
            .in3(N__7505),
            .lcout(\this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8NZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_LC_9_23_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_6_LC_9_23_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_LC_9_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_LC_9_23_6  (
            .in0(N__15504),
            .in1(N__8521),
            .in2(_gnd_net_),
            .in3(N__7502),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_6 ),
            .clk(N__17368),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KAN_LC_9_23_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KAN_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KAN_LC_9_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KAN_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(N__8671),
            .in2(_gnd_net_),
            .in3(N__7499),
            .lcout(\this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KANZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBN_LC_9_24_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBN_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBN_LC_9_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBN_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__8597),
            .in2(_gnd_net_),
            .in3(N__7496),
            .lcout(\this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBNZ0 ),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCN_LC_9_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCN_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCN_LC_9_24_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCN_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__8435),
            .in2(_gnd_net_),
            .in3(N__7493),
            .lcout(\this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_10_17_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_10_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__7998),
            .in2(N__7969),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_2_c_LC_10_17_1 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_2_c_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_2_c_LC_10_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_2_c_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__8256),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_3_c_LC_10_17_2 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_3_c_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_3_c_LC_10_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_3_c_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__8218),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_4_c_LC_10_17_3 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_4_c_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_4_c_LC_10_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_4_c_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__8193),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_5_c_LC_10_17_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_5_c_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_5_c_LC_10_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_5_c_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__8154),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_6_c_LC_10_17_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_6_c_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_6_c_LC_10_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_6_c_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__8774),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_7_LC_10_17_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_10_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_10_17_6  (
            .in0(N__7641),
            .in1(N__8115),
            .in2(_gnd_net_),
            .in3(N__7550),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__17324),
            .ce(),
            .sr(N__15470));
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_8_LC_10_17_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_8_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIDR6I_8_LC_10_17_7 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIDR6I_8_LC_10_17_7  (
            .in0(N__8114),
            .in1(N__8370),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.N_27 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_9_c_LC_10_18_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_9_c_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_9_c_LC_10_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_9_c_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__8836),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_10_LC_10_18_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_10_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_10_LC_10_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_10_LC_10_18_1  (
            .in0(N__7640),
            .in1(N__9214),
            .in2(_gnd_net_),
            .in3(N__7649),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_10 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_9 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_10 ),
            .clk(N__17329),
            .ce(),
            .sr(N__15468));
    defparam \this_vga_signals.M_hcounter_q_11_LC_10_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_11_LC_10_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_11_LC_10_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_11_LC_10_18_2  (
            .in0(N__7639),
            .in1(N__8329),
            .in2(_gnd_net_),
            .in3(N__7610),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17329),
            .ce(),
            .sr(N__15468));
    defparam \this_vga_signals.un17_address_g1_0_0_a2_0_LC_10_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g1_0_0_a2_0_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g1_0_0_a2_0_LC_10_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un17_address_g1_0_0_a2_0_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__13761),
            .in2(_gnd_net_),
            .in3(N__12667),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g1_0_0_a2_LC_10_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g1_0_0_a2_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g1_0_0_a2_LC_10_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g1_0_0_a2_LC_10_19_2  (
            .in0(N__13465),
            .in1(N__18345),
            .in2(N__7607),
            .in3(N__13071),
            .lcout(\this_vga_signals.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_11_1_LC_10_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_11_1_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_11_1_LC_10_19_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un17_address_g0_11_1_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12677),
            .in3(N__18346),
            .lcout(),
            .ltout(\this_vga_signals.g0_11_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_11_LC_10_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_11_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_11_LC_10_19_7 .LUT_INIT=16'b0010000110110111;
    LogicCell40 \this_vga_signals.un17_address_g0_11_LC_10_19_7  (
            .in0(N__13072),
            .in1(N__13760),
            .in2(N__7604),
            .in3(N__13466),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_8_LC_10_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_8_LC_10_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_8_LC_10_20_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_8_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__17685),
            .in2(_gnd_net_),
            .in3(N__7730),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17341),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_7_LC_10_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_7_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_7_LC_10_20_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_7_LC_10_20_2  (
            .in0(N__17686),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7589),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17341),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIPD2J1_5_LC_10_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIPD2J1_5_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIPD2J1_5_LC_10_20_3 .LUT_INIT=16'b0000111101111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIPD2J1_5_LC_10_20_3  (
            .in0(N__9012),
            .in1(N__10539),
            .in2(N__7559),
            .in3(N__8538),
            .lcout(\this_vga_signals.i9_mux ),
            .ltout(\this_vga_signals.i9_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIOO3P7_9_LC_10_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIOO3P7_9_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIOO3P7_9_LC_10_20_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIOO3P7_9_LC_10_20_4  (
            .in0(N__8277),
            .in1(N__8426),
            .in2(N__7826),
            .in3(N__7816),
            .lcout(\this_vga_signals.rgb72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIL6FA3_9_LC_10_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIL6FA3_9_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIL6FA3_9_LC_10_20_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIL6FA3_9_LC_10_20_6  (
            .in0(N__7823),
            .in1(N__8427),
            .in2(_gnd_net_),
            .in3(N__7817),
            .lcout(port_nmib_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_9_LC_10_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_9_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_9_LC_10_21_0 .LUT_INIT=16'b0100011100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_9_LC_10_21_0  (
            .in0(N__9766),
            .in1(N__9727),
            .in2(N__17712),
            .in3(N__7742),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17347),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_10_21_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_10_21_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_10_21_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__7705),
            .in2(_gnd_net_),
            .in3(N__7658),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17347),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_9_LC_10_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_LC_10_21_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_9_LC_10_21_2 .LUT_INIT=16'b0100011100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_LC_10_21_2  (
            .in0(N__9765),
            .in1(N__9726),
            .in2(N__17711),
            .in3(N__7741),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17347),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_8_LC_10_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_LC_10_21_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_LC_10_21_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__17687),
            .in2(_gnd_net_),
            .in3(N__7729),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17347),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_10_21_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_10_21_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_10_21_4 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_10_21_4  (
            .in0(N__7704),
            .in1(N__7667),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17347),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIAGIO1_5_LC_10_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIAGIO1_5_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIAGIO1_5_LC_10_21_6 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIAGIO1_5_LC_10_21_6  (
            .in0(N__10517),
            .in1(N__8647),
            .in2(N__9001),
            .in3(N__8530),
            .lcout(),
            .ltout(\this_vga_signals.address_1_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNILURK2_9_LC_10_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNILURK2_9_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNILURK2_9_LC_10_21_7 .LUT_INIT=16'b1100111111110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNILURK2_9_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__8425),
            .in2(N__7652),
            .in3(N__8589),
            .lcout(\this_vga_signals.N_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_axbxc3_1_LC_10_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_axbxc3_1_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_axbxc3_1_LC_10_22_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_axbxc3_1_LC_10_22_1  (
            .in0(N__7858),
            .in1(N__8063),
            .in2(_gnd_net_),
            .in3(N__7846),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_axbxc1_LC_10_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_axbxc1_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_axbxc1_LC_10_22_2 .LUT_INIT=16'b0111100010000111;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_axbxc1_LC_10_22_2  (
            .in0(N__8531),
            .in1(N__7937),
            .in2(N__8666),
            .in3(N__7904),
            .lcout(\this_vga_signals.mult1_un40_sum_axbxc1 ),
            .ltout(\this_vga_signals.mult1_un40_sum_axbxc1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_10_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_10_22_3 .LUT_INIT=16'b1111111011101010;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_10_22_3  (
            .in0(N__7886),
            .in1(N__8064),
            .in2(N__7880),
            .in3(N__7876),
            .lcout(\this_vga_signals.mult1_un47_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un47_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_10_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_10_22_4 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_10_22_4  (
            .in0(N__9571),
            .in1(_gnd_net_),
            .in2(N__7865),
            .in3(N__11565),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI5CJTF_9_LC_10_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI5CJTF_9_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI5CJTF_9_LC_10_22_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI5CJTF_9_LC_10_22_5  (
            .in0(N__8067),
            .in1(N__8022),
            .in2(N__7862),
            .in3(N__7847),
            .lcout(\this_vga_signals.address_m1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c3_1_LC_10_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c3_1_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c3_1_LC_10_22_6 .LUT_INIT=16'b0001011100101011;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c3_1_LC_10_22_6  (
            .in0(N__8996),
            .in1(N__10522),
            .in2(N__10700),
            .in3(N__11615),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_3_LC_10_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_3_LC_10_23_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_10_23_0 .LUT_INIT=16'b0011010100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_10_23_0  (
            .in0(N__15512),
            .in1(N__9781),
            .in2(N__9725),
            .in3(N__7838),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17359),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc3_1_0_LC_10_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc3_1_0_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc3_1_0_LC_10_23_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc3_1_0_LC_10_23_1  (
            .in0(N__11614),
            .in1(N__8927),
            .in2(N__8027),
            .in3(N__11564),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_m24_ns_1_0_LC_10_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.address_m24_ns_1_0_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_m24_ns_1_0_LC_10_23_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.address_m24_ns_1_0_LC_10_23_2  (
            .in0(N__8899),
            .in1(N__14348),
            .in2(N__7829),
            .in3(N__9825),
            .lcout(),
            .ltout(\this_vga_signals.address_m24_ns_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIS78CB9_2_LC_10_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIS78CB9_2_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIS78CB9_2_LC_10_23_3 .LUT_INIT=16'b0011111011011101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIS78CB9_2_LC_10_23_3  (
            .in0(N__10665),
            .in1(N__9862),
            .in2(N__8078),
            .in3(N__11029),
            .lcout(\this_vga_signals.address_i2_mux_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_axbxc1_LC_10_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_axbxc1_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_axbxc1_LC_10_23_4 .LUT_INIT=16'b0011011011001001;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_axbxc1_LC_10_23_4  (
            .in0(N__10519),
            .in1(N__8514),
            .in2(N__9003),
            .in3(N__8071),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_c2_LC_10_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_c2_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_c2_LC_10_23_5 .LUT_INIT=16'b0011010110010100;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_c2_LC_10_23_5  (
            .in0(N__10521),
            .in1(N__11611),
            .in2(N__9013),
            .in3(N__11562),
            .lcout(\this_vga_signals.mult1_un54_sum_c2 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_c3_LC_10_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_c3_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_c3_LC_10_23_6 .LUT_INIT=16'b1111100110010000;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_c3_LC_10_23_6  (
            .in0(N__11563),
            .in1(N__11613),
            .in2(N__8030),
            .in3(N__8023),
            .lcout(\this_vga_signals.mult1_un54_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c2_LC_10_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c2_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c2_LC_10_23_7 .LUT_INIT=16'b1000111011101000;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c2_LC_10_23_7  (
            .in0(N__10664),
            .in1(N__10520),
            .in2(N__8009),
            .in3(N__8898),
            .lcout(\this_vga_signals.mult1_un61_sum_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_10_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_0_LC_10_24_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_10_24_1 .LUT_INIT=16'b0000010011000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_10_24_1  (
            .in0(N__15511),
            .in1(N__8006),
            .in2(N__9731),
            .in3(N__9780),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17364),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_2_0_LC_10_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_2_0_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_2_0_LC_10_24_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNITV8S_2_0_LC_10_24_3  (
            .in0(_gnd_net_),
            .in1(N__10669),
            .in2(_gnd_net_),
            .in3(N__10791),
            .lcout(\this_vga_signals.M_vcounter_q_RNITV8S_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_0_c_LC_11_17_0 .C_ON=1'b1;
    defparam \this_vga_signals.un12_address_un12_address_cry_0_c_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_0_c_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_0_c_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8000),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\this_vga_signals.un12_address_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_11_17_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_1_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_11_17_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7965),
            .in3(N__7940),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un12_address_cry_0 ),
            .carryout(\this_vga_signals.un12_address_cry_1 ),
            .clk(N__17318),
            .ce(),
            .sr(N__15469));
    defparam \this_vga_signals.un12_address_un12_address_cry_1_c_RNINFAB_LC_11_17_2 .C_ON=1'b1;
    defparam \this_vga_signals.un12_address_un12_address_cry_1_c_RNINFAB_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_1_c_RNINFAB_LC_11_17_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_1_c_RNINFAB_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8258),
            .in3(N__8225),
            .lcout(\this_vga_signals.un12_address_cry_1_c_RNINFAB ),
            .ltout(),
            .carryin(\this_vga_signals.un12_address_cry_1 ),
            .carryout(\this_vga_signals.un12_address_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_2_c_RNIPIBB_LC_11_17_3 .C_ON=1'b1;
    defparam \this_vga_signals.un12_address_un12_address_cry_2_c_RNIPIBB_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_2_c_RNIPIBB_LC_11_17_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_2_c_RNIPIBB_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8222),
            .in3(N__8198),
            .lcout(\this_vga_signals.un12_address_cry_2_c_RNIPIBB ),
            .ltout(),
            .carryin(\this_vga_signals.un12_address_cry_2 ),
            .carryout(\this_vga_signals.un12_address_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIRLCB_LC_11_17_4 .C_ON=1'b1;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIRLCB_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIRLCB_LC_11_17_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_3_c_RNIRLCB_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8195),
            .in3(N__8162),
            .lcout(\this_vga_signals.un12_address_cry_3_c_RNIRLCB ),
            .ltout(),
            .carryin(\this_vga_signals.un12_address_cry_3 ),
            .carryout(\this_vga_signals.un12_address_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNITODB_LC_11_17_5 .C_ON=1'b1;
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNITODB_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNITODB_LC_11_17_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_4_c_RNITODB_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8158),
            .in3(N__8123),
            .lcout(\this_vga_signals.un12_address_cry_4_c_RNITODB ),
            .ltout(),
            .carryin(\this_vga_signals.un12_address_cry_4 ),
            .carryout(\this_vga_signals.un12_address_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_5_c_RNIVREB_LC_11_17_6 .C_ON=1'b1;
    defparam \this_vga_signals.un12_address_un12_address_cry_5_c_RNIVREB_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_5_c_RNIVREB_LC_11_17_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_5_c_RNIVREB_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8777),
            .in3(N__8120),
            .lcout(\this_vga_signals.un12_address_cry_5_c_RNIVREB ),
            .ltout(),
            .carryin(\this_vga_signals.un12_address_cry_5 ),
            .carryout(\this_vga_signals.un12_address_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_6_c_RNI1VFB_LC_11_17_7 .C_ON=1'b1;
    defparam \this_vga_signals.un12_address_un12_address_cry_6_c_RNI1VFB_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_6_c_RNI1VFB_LC_11_17_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_6_c_RNI1VFB_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8116),
            .in3(N__8090),
            .lcout(\this_vga_signals.if_m1_0_0 ),
            .ltout(),
            .carryin(\this_vga_signals.un12_address_cry_6 ),
            .carryout(\this_vga_signals.un12_address_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_7_c_RNI32HB_LC_11_18_0 .C_ON=1'b1;
    defparam \this_vga_signals.un12_address_un12_address_cry_7_c_RNI32HB_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_7_c_RNI32HB_LC_11_18_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_7_c_RNI32HB_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8371),
            .in3(N__8087),
            .lcout(\this_vga_signals.un12_address_cry_7_c_RNI32HB ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\this_vga_signals.un12_address_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_8_c_RNI55IB_LC_11_18_1 .C_ON=1'b1;
    defparam \this_vga_signals.un12_address_un12_address_cry_8_c_RNI55IB_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_8_c_RNI55IB_LC_11_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_8_c_RNI55IB_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__18650),
            .in2(N__8846),
            .in3(N__8084),
            .lcout(\this_vga_signals.mult1_un54_sum_axb3_out ),
            .ltout(),
            .carryin(\this_vga_signals.un12_address_cry_8 ),
            .carryout(\this_vga_signals.un12_address_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_cry_9_THRU_LUT4_0_LC_11_18_2 .C_ON=1'b1;
    defparam \this_vga_signals.un12_address_cry_9_THRU_LUT4_0_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_cry_9_THRU_LUT4_0_LC_11_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.un12_address_cry_9_THRU_LUT4_0_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__9200),
            .in2(N__18673),
            .in3(N__8081),
            .lcout(\this_vga_signals.un12_address_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\this_vga_signals.un12_address_cry_9 ),
            .carryout(\this_vga_signals.un12_address_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_10_c_RNINP5K_LC_11_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_10_c_RNINP5K_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_10_c_RNINP5K_LC_11_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_10_c_RNINP5K_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__9170),
            .in2(_gnd_net_),
            .in3(N__8378),
            .lcout(\this_vga_signals.un12_address_cry_10_c_RNINP5K ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10149),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17325),
            .ce(),
            .sr(N__15467));
    defparam \this_vga_signals.M_hcounter_q_RNI3IKE4_11_LC_11_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI3IKE4_11_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI3IKE4_11_LC_11_19_0 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI3IKE4_11_LC_11_19_0  (
            .in0(N__9146),
            .in1(N__8348),
            .in2(N__8330),
            .in3(N__8723),
            .lcout(N_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_1_0_LC_11_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_1_0_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_1_0_LC_11_19_1 .LUT_INIT=16'b1110000111000011;
    LogicCell40 \this_vga_signals.un17_address_g0_1_0_LC_11_19_1  (
            .in0(N__12030),
            .in1(N__11832),
            .in2(N__13452),
            .in3(N__10239),
            .lcout(\this_vga_signals.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_2L1_LC_11_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_2L1_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_2L1_LC_11_19_2 .LUT_INIT=16'b0011001101100110;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_2L1_LC_11_19_2  (
            .in0(N__11833),
            .in1(N__12031),
            .in2(_gnd_net_),
            .in3(N__11760),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axbxc5_LC_11_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axbxc5_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axbxc5_LC_11_19_3 .LUT_INIT=16'b0000000000111111;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axbxc5_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__11989),
            .in2(N__10244),
            .in3(N__11831),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_1_1_LC_11_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_1_1_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_1_1_LC_11_19_4 .LUT_INIT=16'b0110011011011101;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_1_1_LC_11_19_4  (
            .in0(N__10002),
            .in1(N__9392),
            .in2(_gnd_net_),
            .in3(N__9429),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_7_0_3_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_LC_11_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_LC_11_19_5 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_LC_11_19_5  (
            .in0(N__10140),
            .in1(N__8858),
            .in2(N__8261),
            .in3(N__9145),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_7_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_7_c_RNI8RAPK_LC_11_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_7_c_RNI8RAPK_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_7_c_RNI8RAPK_LC_11_19_6 .LUT_INIT=16'b0100101000011010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_7_c_RNI8RAPK_LC_11_19_6  (
            .in0(N__11834),
            .in1(N__9227),
            .in2(N__12025),
            .in3(N__10141),
            .lcout(\this_vga_signals.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_2_LC_11_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_2_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_2_LC_11_19_7 .LUT_INIT=16'b0101000000001010;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_2_LC_11_19_7  (
            .in0(N__9393),
            .in1(_gnd_net_),
            .in2(N__9434),
            .in3(N__10001),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_7_0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIAIMG1_6_LC_11_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIAIMG1_6_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIAIMG1_6_LC_11_20_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIAIMG1_6_LC_11_20_3  (
            .in0(N__9220),
            .in1(N__8852),
            .in2(N__8800),
            .in3(N__8773),
            .lcout(\this_vga_signals.hvisible_i_a2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_26_LC_11_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_26_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_26_LC_11_20_5 .LUT_INIT=16'b0011001101000100;
    LogicCell40 \this_vga_signals.un17_address_g0_26_LC_11_20_5  (
            .in0(N__10243),
            .in1(N__12032),
            .in2(_gnd_net_),
            .in3(N__11847),
            .lcout(\this_vga_signals.g0_6_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI7A9S_7_LC_11_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI7A9S_7_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI7A9S_7_LC_11_21_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI7A9S_7_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__8670),
            .in2(_gnd_net_),
            .in3(N__8540),
            .lcout(\this_vga_signals.m30_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI0FV6Q_11_LC_11_21_1 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI0FV6Q_11_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI0FV6Q_11_LC_11_21_1 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \this_vram.mem_radreg_RNI0FV6Q_11_LC_11_21_1  (
            .in0(N__16984),
            .in1(N__17799),
            .in2(N__14500),
            .in3(N__17011),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI39IO1_1_LC_11_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI39IO1_1_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI39IO1_1_LC_11_21_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI39IO1_1_LC_11_21_4  (
            .in0(N__10823),
            .in1(N__9014),
            .in2(N__10913),
            .in3(N__8428),
            .lcout(),
            .ltout(\this_vga_signals.m30_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIEQ4H3_8_LC_11_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIEQ4H3_8_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIEQ4H3_8_LC_11_21_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIEQ4H3_8_LC_11_21_5  (
            .in0(N__8681),
            .in1(N__11026),
            .in2(N__8675),
            .in3(N__8591),
            .lcout(\this_vga_signals.N_75_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIS0EA1_8_LC_11_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIS0EA1_8_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIS0EA1_8_LC_11_22_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIS0EA1_8_LC_11_22_0  (
            .in0(N__8672),
            .in1(N__8590),
            .in2(_gnd_net_),
            .in3(N__8539),
            .lcout(),
            .ltout(\this_vga_signals.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIHQRK2_9_LC_11_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIHQRK2_9_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIHQRK2_9_LC_11_22_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIHQRK2_9_LC_11_22_1  (
            .in0(N__10829),
            .in1(N__9008),
            .in2(N__8438),
            .in3(N__8429),
            .lcout(\this_vga_signals.N_72_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_11_LC_11_22_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_11_LC_11_22_2 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_11_LC_11_22_2 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \this_vram.mem_radreg_11_LC_11_22_2  (
            .in0(N__19946),
            .in1(N__8900),
            .in2(_gnd_net_),
            .in3(N__9831),
            .lcout(\this_vram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17348),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI0FV6Q_0_11_LC_11_22_3 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI0FV6Q_0_11_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI0FV6Q_0_11_LC_11_22_3 .LUT_INIT=16'b0100000001110000;
    LogicCell40 \this_vram.mem_radreg_RNI0FV6Q_0_11_LC_11_22_3  (
            .in0(N__16985),
            .in1(N__17798),
            .in2(N__14501),
            .in3(N__17015),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_22_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_22_4  (
            .in0(N__9007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11612),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_11_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_11_23_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_11_23_0  (
            .in0(N__9098),
            .in1(N__8897),
            .in2(N__9119),
            .in3(N__9824),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQVOIR1_2_LC_11_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQVOIR1_2_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQVOIR1_2_LC_11_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQVOIR1_2_LC_11_23_1  (
            .in0(N__8933),
            .in1(N__11622),
            .in2(N__11016),
            .in3(N__8926),
            .lcout(\this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2 ),
            .ltout(\this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI495CI5_2_LC_11_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI495CI5_2_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI495CI5_2_LC_11_23_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI495CI5_2_LC_11_23_2  (
            .in0(N__9822),
            .in1(N__9117),
            .in2(N__8915),
            .in3(N__8895),
            .lcout(\this_vga_signals.address_i3_mux_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c3_LC_11_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c3_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c3_LC_11_23_3 .LUT_INIT=16'b1000111001001101;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c3_LC_11_23_3  (
            .in0(N__8894),
            .in1(N__9113),
            .in2(N__8912),
            .in3(N__9820),
            .lcout(\this_vga_signals.mult1_un61_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_m1_LC_11_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.address_m1_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_m1_LC_11_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.address_m1_LC_11_23_4  (
            .in0(N__8867),
            .in1(N__8896),
            .in2(N__8903),
            .in3(N__9823),
            .lcout(\this_vga_signals.address_mZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_11_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_11_23_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_11_23_5  (
            .in0(N__8893),
            .in1(N__9821),
            .in2(_gnd_net_),
            .in3(N__8866),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_c2_LC_11_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_c2_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_c2_LC_11_23_6 .LUT_INIT=16'b0100110111010100;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_c2_LC_11_23_6  (
            .in0(N__10733),
            .in1(N__10986),
            .in2(N__9122),
            .in3(N__14353),
            .lcout(\this_vga_signals.mult1_un68_sum_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI9MJK5B_2_LC_11_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI9MJK5B_2_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI9MJK5B_2_LC_11_23_7 .LUT_INIT=16'b0000011010011111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI9MJK5B_2_LC_11_23_7  (
            .in0(N__9118),
            .in1(N__9097),
            .in2(N__9089),
            .in3(N__9080),
            .lcout(\this_vga_signals.address_N_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIDN3UA9_3_LC_11_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIDN3UA9_3_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIDN3UA9_3_LC_11_24_0 .LUT_INIT=16'b0011010111000101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIDN3UA9_3_LC_11_24_0  (
            .in0(N__10667),
            .in1(N__14352),
            .in2(N__9635),
            .in3(N__14289),
            .lcout(),
            .ltout(\this_vga_signals.address_m27_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI2U4THK_2_LC_11_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI2U4THK_2_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI2U4THK_2_LC_11_24_1 .LUT_INIT=16'b0100000101110001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI2U4THK_2_LC_11_24_1  (
            .in0(N__11002),
            .in1(N__9633),
            .in2(N__9074),
            .in3(N__9527),
            .lcout(),
            .ltout(\this_vga_signals.address_i2_mux_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNICBPF381_2_LC_11_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNICBPF381_2_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNICBPF381_2_LC_11_24_2 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNICBPF381_2_LC_11_24_2  (
            .in0(N__11048),
            .in1(N__10856),
            .in2(N__9071),
            .in3(N__9068),
            .lcout(\this_vga_signals.address_m35_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_1_0_LC_11_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_1_0_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_1_0_LC_11_24_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNITV8S_1_0_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__10790),
            .in2(_gnd_net_),
            .in3(N__10666),
            .lcout(\this_vga_signals.M_vcounter_q_RNITV8S_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_0_LC_11_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_0_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_0_LC_11_24_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNITV8S_0_LC_11_24_4  (
            .in0(N__10668),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10821),
            .lcout(\this_vga_signals.address_m31_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_1_LC_11_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_1_LC_11_24_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_11_24_5 .LUT_INIT=16'b0101001100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_11_24_5  (
            .in0(N__9779),
            .in1(N__15510),
            .in2(N__9724),
            .in3(N__9062),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17360),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axb4_LC_12_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axb4_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axb4_LC_12_17_0 .LUT_INIT=16'b1101101110110110;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axb4_LC_12_17_0  (
            .in0(N__9998),
            .in1(N__9424),
            .in2(N__9395),
            .in3(N__9142),
            .lcout(\this_vga_signals.mult1_un54_sum_axb4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g1_LC_12_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g1_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g1_LC_12_17_1 .LUT_INIT=16'b0000101001010000;
    LogicCell40 \this_vga_signals.un17_address_g1_LC_12_17_1  (
            .in0(N__9143),
            .in1(_gnd_net_),
            .in2(N__9433),
            .in3(N__9390),
            .lcout(\this_vga_signals.g1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_30_LC_12_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_30_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_30_LC_12_17_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \this_vga_signals.un17_address_g0_30_LC_12_17_2  (
            .in0(N__13399),
            .in1(N__11954),
            .in2(_gnd_net_),
            .in3(N__10240),
            .lcout(\this_vga_signals.if_m4_0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_ac0_8_LC_12_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_ac0_8_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_ac0_8_LC_12_17_4 .LUT_INIT=16'b0010000000001000;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_ac0_8_LC_12_17_4  (
            .in0(N__9997),
            .in1(N__9423),
            .in2(N__9394),
            .in3(N__9141),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_8 ),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_x0_LC_12_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_x0_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_x0_LC_12_17_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_x0_LC_12_17_5  (
            .in0(N__10128),
            .in1(N__9999),
            .in2(N__9230),
            .in3(N__9919),
            .lcout(\this_vga_signals.mult1_un61_sum_axb4_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g1_1_LC_12_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g1_1_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g1_1_LC_12_17_6 .LUT_INIT=16'b0010001001000100;
    LogicCell40 \this_vga_signals.un17_address_g1_1_LC_12_17_6  (
            .in0(N__9391),
            .in1(N__9428),
            .in2(_gnd_net_),
            .in3(N__9144),
            .lcout(\this_vga_signals.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_x1_LC_12_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_x1_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_x1_LC_12_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_x1_LC_12_17_7  (
            .in0(N__10129),
            .in1(N__10000),
            .in2(_gnd_net_),
            .in3(N__9918),
            .lcout(\this_vga_signals.mult1_un61_sum_axb4_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axbxc5_LC_12_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axbxc5_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axbxc5_LC_12_18_0 .LUT_INIT=16'b1001110000111001;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axbxc5_LC_12_18_0  (
            .in0(N__9996),
            .in1(N__9945),
            .in2(N__10150),
            .in3(N__9925),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_9_c_RNIEJOE_LC_12_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_9_c_RNIEJOE_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_9_c_RNIEJOE_LC_12_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_9_c_RNIEJOE_LC_12_18_1  (
            .in0(N__9216),
            .in1(N__18646),
            .in2(_gnd_net_),
            .in3(N__9155),
            .lcout(\this_vga_signals.un12_address_cry_9_c_RNIEJOE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g1_2_LC_12_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g1_2_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g1_2_LC_12_18_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \this_vga_signals.un17_address_g1_2_LC_12_18_2  (
            .in0(N__11401),
            .in1(N__10042),
            .in2(_gnd_net_),
            .in3(N__10024),
            .lcout(\this_vga_signals.g1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_9_c_RNIVF1R_LC_12_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_9_c_RNIVF1R_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_9_c_RNIVF1R_LC_12_18_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_9_c_RNIVF1R_LC_12_18_3  (
            .in0(N__9215),
            .in1(N__9169),
            .in2(_gnd_net_),
            .in3(N__9154),
            .lcout(\this_vga_signals.un12_address_cry_9_c_RNIVF1R ),
            .ltout(\this_vga_signals.un12_address_cry_9_c_RNIVF1R_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un47_sum_ac0_7_LC_12_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un47_sum_ac0_7_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un47_sum_ac0_7_LC_12_18_4 .LUT_INIT=16'b1011001000101100;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un47_sum_ac0_7_LC_12_18_4  (
            .in0(N__9995),
            .in1(N__9422),
            .in2(N__9398),
            .in3(N__9383),
            .lcout(\this_vga_signals.mult1_un47_sum_c5 ),
            .ltout(\this_vga_signals.mult1_un47_sum_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb3_x1_LC_12_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb3_x1_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb3_x1_LC_12_18_5 .LUT_INIT=16'b0011001110000001;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb3_x1_LC_12_18_5  (
            .in0(N__10023),
            .in1(N__10130),
            .in2(N__9359),
            .in3(N__12231),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axb3_x1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb3_ns_LC_12_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb3_ns_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb3_ns_LC_12_18_6 .LUT_INIT=16'b1111000001100110;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb3_ns_LC_12_18_6  (
            .in0(N__12232),
            .in1(N__10158),
            .in2(N__9356),
            .in3(N__9944),
            .lcout(\this_vga_signals.mult1_un61_sum_axb3 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axb3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m5_sn_LC_12_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m5_sn_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m5_sn_LC_12_18_7 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \this_vga_signals.un17_address_if_m5_sn_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__13349),
            .in2(N__9353),
            .in3(N__11953),
            .lcout(\this_vga_signals.if_m5_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m5_rn_LC_12_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m5_rn_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m5_rn_LC_12_19_0 .LUT_INIT=16'b0000111111111010;
    LogicCell40 \this_vga_signals.un17_address_if_m5_rn_LC_12_19_0  (
            .in0(N__13400),
            .in1(_gnd_net_),
            .in2(N__12034),
            .in3(N__10235),
            .lcout(),
            .ltout(\this_vga_signals.if_m5_rn_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m5_mb_LC_12_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m5_mb_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m5_mb_LC_12_19_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \this_vga_signals.un17_address_if_m5_mb_LC_12_19_1  (
            .in0(N__11724),
            .in1(N__9350),
            .in2(N__9344),
            .in3(N__11835),
            .lcout(\this_vga_signals.mult1_un68_sum_c5 ),
            .ltout(\this_vga_signals.mult1_un68_sum_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un75_sum_axb3_LC_12_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un75_sum_axb3_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un75_sum_axb3_LC_12_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un75_sum_axb3_LC_12_19_2  (
            .in0(N__13401),
            .in1(N__12589),
            .in2(N__9341),
            .in3(N__18310),
            .lcout(\this_vga_signals.mult1_un75_sum_axb3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_c4_LC_12_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_c4_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_c4_LC_12_19_3 .LUT_INIT=16'b0010001010111011;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_c4_LC_12_19_3  (
            .in0(N__10142),
            .in1(N__10011),
            .in2(_gnd_net_),
            .in3(N__9920),
            .lcout(\this_vga_signals.mult1_un54_sum_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIAFTT93_9_LC_12_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIAFTT93_9_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIAFTT93_9_LC_12_19_4 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIAFTT93_9_LC_12_19_4  (
            .in0(N__12637),
            .in1(N__18311),
            .in2(N__19985),
            .in3(N__13062),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_12_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_12_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_12_19_5  (
            .in0(N__10143),
            .in1(N__10012),
            .in2(_gnd_net_),
            .in3(N__9921),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_4_LC_12_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_4_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_4_LC_12_19_6 .LUT_INIT=16'b1110110011011100;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_4_LC_12_19_6  (
            .in0(N__9950),
            .in1(N__9458),
            .in2(N__9452),
            .in3(N__9449),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_7_0_4 ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_7_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m1_0_LC_12_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m1_0_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m1_0_LC_12_19_7 .LUT_INIT=16'b0000010111110000;
    LogicCell40 \this_vga_signals.un17_address_if_m1_0_LC_12_19_7  (
            .in0(N__10234),
            .in1(_gnd_net_),
            .in2(N__9443),
            .in3(N__12017),
            .lcout(\this_vga_signals.if_m1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_i_o2_0_x2_LC_12_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_i_o2_0_x2_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_i_o2_0_x2_LC_12_20_0 .LUT_INIT=16'b1010100101010110;
    LogicCell40 \this_vga_signals.un17_address_g0_i_o2_0_x2_LC_12_20_0  (
            .in0(N__13042),
            .in1(N__11851),
            .in2(N__11761),
            .in3(N__12675),
            .lcout(\this_vga_signals.N_26_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m4_0_1_LC_12_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m4_0_1_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m4_0_1_LC_12_20_1 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \this_vga_signals.un17_address_if_m4_0_1_LC_12_20_1  (
            .in0(N__13402),
            .in1(N__11993),
            .in2(_gnd_net_),
            .in3(N__10241),
            .lcout(\this_vga_signals.if_m4_0_1 ),
            .ltout(\this_vga_signals.if_m4_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_25_LC_12_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_25_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_25_LC_12_20_2 .LUT_INIT=16'b1111111011100000;
    LogicCell40 \this_vga_signals.un17_address_g0_25_LC_12_20_2  (
            .in0(N__11755),
            .in1(N__11852),
            .in2(N__9440),
            .in3(N__11995),
            .lcout(\this_vga_signals.if_N_8_mux_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_6_c_RNIGPBEN_LC_12_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_6_c_RNIGPBEN_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_6_c_RNIGPBEN_LC_12_20_3 .LUT_INIT=16'b0001111000111100;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_6_c_RNIGPBEN_LC_12_20_3  (
            .in0(N__11994),
            .in1(N__11839),
            .in2(N__13451),
            .in3(N__10242),
            .lcout(\this_vga_signals.G_12_0_x3_0 ),
            .ltout(\this_vga_signals.G_12_0_x3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNI913733_LC_12_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNI913733_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNI913733_LC_12_20_4 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_3_c_RNI913733_LC_12_20_4  (
            .in0(N__13043),
            .in1(N__12907),
            .in2(N__9437),
            .in3(N__13300),
            .lcout(\this_vga_signals.G_12_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_38_LC_12_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_38_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_38_LC_12_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un17_address_g0_38_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(N__12651),
            .in2(N__18348),
            .in3(N__13041),
            .lcout(\this_vga_signals.g0_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_2_LC_12_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_2_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_2_LC_12_20_7 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_0_2_LC_12_20_7  (
            .in0(N__11996),
            .in1(N__11840),
            .in2(N__12945),
            .in3(N__11756),
            .lcout(\this_vga_signals.g0_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNITHP2_0_LC_12_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNITHP2_0_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNITHP2_0_LC_12_21_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNITHP2_0_LC_12_21_0  (
            .in0(N__10571),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9602),
            .lcout(vsync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_0_1_LC_12_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_0_1_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_0_1_LC_12_21_1 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_0_1_LC_12_21_1  (
            .in0(N__9600),
            .in1(N__9764),
            .in2(_gnd_net_),
            .in3(N__9488),
            .lcout(),
            .ltout(\this_vga_signals.N_52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_1_LC_12_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_1_LC_12_21_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vstate_q_1_LC_12_21_2 .LUT_INIT=16'b0000000001001110;
    LogicCell40 \this_vga_signals.M_vstate_q_1_LC_12_21_2  (
            .in0(N__10469),
            .in1(N__9601),
            .in2(N__9491),
            .in3(N__17709),
            .lcout(\this_vga_signals.M_vstate_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17337),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIEQ4H3_1_LC_12_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIEQ4H3_1_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIEQ4H3_1_LC_12_21_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIEQ4H3_1_LC_12_21_3  (
            .in0(N__9479),
            .in1(N__10904),
            .in2(_gnd_net_),
            .in3(N__11027),
            .lcout(\this_vga_signals.N_76_mux ),
            .ltout(\this_vga_signals.N_76_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_2_0_LC_12_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_2_0_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_2_0_LC_12_21_4 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_2_0_LC_12_21_4  (
            .in0(N__9763),
            .in1(N__9598),
            .in2(N__9482),
            .in3(N__10743),
            .lcout(\this_vga_signals.M_vstate_q_RNO_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_3_0_LC_12_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_3_0_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_3_0_LC_12_21_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_3_0_LC_12_21_5  (
            .in0(N__9478),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10903),
            .lcout(),
            .ltout(\this_vga_signals.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_1_0_LC_12_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_1_0_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_1_0_LC_12_21_6 .LUT_INIT=16'b0111111111101111;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_1_0_LC_12_21_6  (
            .in0(N__11028),
            .in1(N__9599),
            .in2(N__9470),
            .in3(N__10742),
            .lcout(),
            .ltout(\this_vga_signals.M_vstate_q_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_0_0_LC_12_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_0_0_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_0_0_LC_12_21_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_0_0_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(N__10570),
            .in2(N__9467),
            .in3(N__9464),
            .lcout(\this_vga_signals.N_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI149S_4_LC_12_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI149S_4_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI149S_4_LC_12_22_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI149S_4_LC_12_22_0  (
            .in0(N__10538),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10739),
            .lcout(),
            .ltout(\this_vga_signals.m35_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNI4LE61_0_LC_12_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNI4LE61_0_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNI4LE61_0_LC_12_22_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNI4LE61_0_LC_12_22_1  (
            .in0(N__9597),
            .in1(N__10567),
            .in2(N__9578),
            .in3(N__15503),
            .lcout(\this_vga_signals.N_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_12_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_12_22_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_12_22_4  (
            .in0(N__14285),
            .in1(N__9560),
            .in2(N__9551),
            .in3(N__14357),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIV7VFA9_0_2_LC_12_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIV7VFA9_0_2_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIV7VFA9_0_2_LC_12_22_5 .LUT_INIT=16'b1001010001100001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIV7VFA9_0_2_LC_12_22_5  (
            .in0(N__11023),
            .in1(N__14351),
            .in2(N__10748),
            .in3(N__14284),
            .lcout(\this_vga_signals.address_N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axb1_0_LC_12_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axb1_0_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axb1_0_LC_12_22_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axb1_0_LC_12_22_6  (
            .in0(N__9575),
            .in1(N__11623),
            .in2(N__10545),
            .in3(N__11572),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_12_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_12_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_12_23_0  (
            .in0(N__9833),
            .in1(N__10732),
            .in2(_gnd_net_),
            .in3(N__9842),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_c3_LC_12_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_c3_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_c3_LC_12_23_1 .LUT_INIT=16'b1111100110010000;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_c3_LC_12_23_1  (
            .in0(N__14288),
            .in1(N__14358),
            .in2(N__9554),
            .in3(N__9550),
            .lcout(\this_vga_signals.mult1_un68_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIV7VFA9_1_2_LC_12_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIV7VFA9_1_2_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIV7VFA9_1_2_LC_12_23_2 .LUT_INIT=16'b0100001000011000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIV7VFA9_1_2_LC_12_23_2  (
            .in0(N__10992),
            .in1(N__14349),
            .in2(N__10735),
            .in3(N__14286),
            .lcout(\this_vga_signals.address_N_9_0 ),
            .ltout(\this_vga_signals.address_N_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIBU2ELI_0_0_LC_12_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIBU2ELI_0_0_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIBU2ELI_0_0_LC_12_23_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIBU2ELI_0_0_LC_12_23_3  (
            .in0(N__10828),
            .in1(_gnd_net_),
            .in2(N__9536),
            .in3(N__9533),
            .lcout(\this_vga_signals.address_N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI8OSG6B_2_LC_12_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI8OSG6B_2_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI8OSG6B_2_LC_12_23_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI8OSG6B_2_LC_12_23_4  (
            .in0(N__10993),
            .in1(N__10731),
            .in2(_gnd_net_),
            .in3(N__9526),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_RNI8OSG6BZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI5UR0HK_2_LC_12_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI5UR0HK_2_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI5UR0HK_2_LC_12_23_5 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI5UR0HK_2_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(N__9866),
            .in2(N__9845),
            .in3(N__10339),
            .lcout(\this_vga_signals.address_i2_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_12_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_12_23_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_12_23_6  (
            .in0(N__10864),
            .in1(N__14350),
            .in2(_gnd_net_),
            .in3(N__14287),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axb1_LC_12_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axb1_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axb1_LC_12_23_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axb1_LC_12_23_7  (
            .in0(N__9841),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9832),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI4G7F3B2_0_LC_12_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI4G7F3B2_0_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI4G7F3B2_0_LC_12_24_1 .LUT_INIT=16'b1010000011001111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI4G7F3B2_0_LC_12_24_1  (
            .in0(N__9641),
            .in1(N__9608),
            .in2(N__10871),
            .in3(N__9788),
            .lcout(\this_vga_signals.address_N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_2_LC_12_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_2_LC_12_24_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_12_24_2 .LUT_INIT=16'b0011010100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_12_24_2  (
            .in0(N__15509),
            .in1(N__9782),
            .in2(N__9709),
            .in3(N__9662),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17353),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI9MCQB9_2_LC_12_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI9MCQB9_2_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI9MCQB9_2_LC_12_24_4 .LUT_INIT=16'b1100110000101111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI9MCQB9_2_LC_12_24_4  (
            .in0(N__10619),
            .in1(N__10998),
            .in2(N__9650),
            .in3(N__10334),
            .lcout(\this_vga_signals.address_i2_mux_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIS78CB9_0_2_LC_12_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIS78CB9_0_2_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIS78CB9_0_2_LC_12_24_5 .LUT_INIT=16'b0000100100111000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIS78CB9_0_2_LC_12_24_5  (
            .in0(N__10335),
            .in1(N__9634),
            .in2(N__11024),
            .in3(N__10747),
            .lcout(\this_vga_signals.address_i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIV7VFA9_2_LC_12_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIV7VFA9_2_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIV7VFA9_2_LC_12_24_6 .LUT_INIT=16'b1011101101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIV7VFA9_2_LC_12_24_6  (
            .in0(N__10746),
            .in1(N__10997),
            .in2(_gnd_net_),
            .in3(N__10333),
            .lcout(),
            .ltout(\this_vga_signals.address_N_33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIBU2ELI_0_LC_12_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIBU2ELI_0_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIBU2ELI_0_LC_12_24_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIBU2ELI_0_LC_12_24_7  (
            .in0(N__9617),
            .in1(_gnd_net_),
            .in2(N__9611),
            .in3(N__10822),
            .lcout(\this_vga_signals.address_N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_4_LC_13_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_4_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_4_LC_13_17_0 .LUT_INIT=16'b0001001111101100;
    LogicCell40 \this_vga_signals.un17_address_g0_4_LC_13_17_0  (
            .in0(N__10028),
            .in1(N__11394),
            .in2(N__10058),
            .in3(N__10165),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axb3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_4_0_1_LC_13_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_4_0_1_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_4_0_1_LC_13_17_1 .LUT_INIT=16'b0001000100001000;
    LogicCell40 \this_vga_signals.un17_address_g0_4_0_1_LC_13_17_1  (
            .in0(N__12023),
            .in1(N__10310),
            .in2(N__10049),
            .in3(N__11864),
            .lcout(),
            .ltout(\this_vga_signals.g0_4_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_4_0_LC_13_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_4_0_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_4_0_LC_13_17_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un17_address_g0_4_0_LC_13_17_2  (
            .in0(N__13449),
            .in1(N__12628),
            .in2(N__10046),
            .in3(N__13083),
            .lcout(\this_vga_signals.g0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_2_LC_13_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_2_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_2_LC_13_17_3 .LUT_INIT=16'b0001111001011010;
    LogicCell40 \this_vga_signals.un17_address_g0_2_LC_13_17_3  (
            .in0(N__11393),
            .in1(N__10027),
            .in2(N__10166),
            .in3(N__10043),
            .lcout(\this_vga_signals.mult1_un61_sum_axb3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_ac0_7_LC_13_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_ac0_7_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_ac0_7_LC_13_17_4 .LUT_INIT=16'b0100110000000100;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_ac0_7_LC_13_17_4  (
            .in0(N__10026),
            .in1(N__9946),
            .in2(N__9926),
            .in3(N__10161),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_7 ),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_ns_LC_13_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_ns_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_ns_LC_13_17_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_ns_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__9893),
            .in2(N__9887),
            .in3(N__9884),
            .lcout(\this_vga_signals.mult1_un61_sum_axb4_i ),
            .ltout(\this_vga_signals.mult1_un61_sum_axb4_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m2_3_0_LC_13_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m2_3_0_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m2_3_0_LC_13_17_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un17_address_if_m2_3_0_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9878),
            .in3(N__10222),
            .lcout(\this_vga_signals.if_m2_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_5_LC_13_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_5_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_5_LC_13_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_5_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__12000),
            .in2(_gnd_net_),
            .in3(N__10223),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_5 ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_13_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_13_18_1 .LUT_INIT=16'b1111010000001011;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_13_18_1  (
            .in0(N__10159),
            .in1(N__10174),
            .in2(N__9875),
            .in3(N__9872),
            .lcout(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0),
            .ltout(this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_0_a2_1_LC_13_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_0_a2_1_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_0_a2_1_LC_13_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_0_0_a2_1_LC_13_18_2  (
            .in0(N__10259),
            .in1(N__12832),
            .in2(N__10247),
            .in3(N__12806),
            .lcout(\this_vga_signals.g0_0_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_21_LC_13_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_21_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_21_LC_13_18_3 .LUT_INIT=16'b0000111101010000;
    LogicCell40 \this_vga_signals.un17_address_g0_21_LC_13_18_3  (
            .in0(N__10224),
            .in1(_gnd_net_),
            .in2(N__12029),
            .in3(N__11845),
            .lcout(\this_vga_signals.g0_6_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_41_LC_13_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_41_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_41_LC_13_18_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \this_vga_signals.un17_address_g0_41_LC_13_18_4  (
            .in0(N__12012),
            .in1(N__13471),
            .in2(_gnd_net_),
            .in3(N__10225),
            .lcout(),
            .ltout(\this_vga_signals.if_m4_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_15_LC_13_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_15_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_15_LC_13_18_5 .LUT_INIT=16'b1111110011101000;
    LogicCell40 \this_vga_signals.un17_address_g0_15_LC_13_18_5  (
            .in0(N__11723),
            .in1(N__12013),
            .in2(N__10178),
            .in3(N__11846),
            .lcout(\this_vga_signals.if_N_8_mux_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m2_3_LC_13_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m2_3_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m2_3_LC_13_18_6 .LUT_INIT=16'b0000111111010010;
    LogicCell40 \this_vga_signals.un17_address_if_m2_3_LC_13_18_6  (
            .in0(N__10175),
            .in1(N__10160),
            .in2(N__10082),
            .in3(N__11722),
            .lcout(\this_vga_signals.if_N_3_3_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_6_1_LC_13_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_6_1_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_6_1_LC_13_18_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \this_vga_signals.un17_address_g0_6_1_LC_13_18_7  (
            .in0(N__13470),
            .in1(N__10073),
            .in2(_gnd_net_),
            .in3(N__11844),
            .lcout(\this_vga_signals.g0_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_16_LC_13_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_16_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_16_LC_13_19_0 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \this_vga_signals.un17_address_g0_16_LC_13_19_0  (
            .in0(N__11728),
            .in1(N__11837),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.N_21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNIU8UQ04_0_LC_13_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNIU8UQ04_0_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNIU8UQ04_0_LC_13_19_1 .LUT_INIT=16'b1001000101100100;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_4_c_RNIU8UQ04_0_LC_13_19_1  (
            .in0(N__12600),
            .in1(N__12315),
            .in2(N__13802),
            .in3(N__12805),
            .lcout(),
            .ltout(\this_vga_signals.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIKCM73C_LC_13_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIKCM73C_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIKCM73C_LC_13_19_2 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_3_c_RNIKCM73C_LC_13_19_2  (
            .in0(N__10292),
            .in1(N__10067),
            .in2(N__10061),
            .in3(N__13288),
            .lcout(),
            .ltout(\this_vga_signals.G_12_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIRBMU931_LC_13_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIRBMU931_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIRBMU931_LC_13_19_3 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_3_c_RNIRBMU931_LC_13_19_3  (
            .in0(N__13554),
            .in1(N__10283),
            .in2(N__10313),
            .in3(N__10583),
            .lcout(\this_vga_signals.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m4_0_LC_13_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m4_0_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m4_0_LC_13_19_4 .LUT_INIT=16'b1111111010101000;
    LogicCell40 \this_vga_signals.un17_address_if_m4_0_LC_13_19_4  (
            .in0(N__12021),
            .in1(N__11836),
            .in2(N__11747),
            .in3(N__10306),
            .lcout(this_vga_signals_un17_address_if_N_8_mux),
            .ltout(this_vga_signals_un17_address_if_N_8_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNIU8UQ04_LC_13_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNIU8UQ04_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNIU8UQ04_LC_13_19_5 .LUT_INIT=16'b1010010001001010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_4_c_RNIU8UQ04_LC_13_19_5  (
            .in0(N__12599),
            .in1(N__13748),
            .in2(N__10295),
            .in3(N__12804),
            .lcout(\this_vga_signals.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_i_x4_4_a3_1_LC_13_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_i_x4_4_a3_1_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_i_x4_4_a3_1_LC_13_19_6 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_i_x4_4_a3_1_LC_13_19_6  (
            .in0(N__12022),
            .in1(N__13553),
            .in2(N__11748),
            .in3(N__11838),
            .lcout(\this_vga_signals.g0_i_x4_4_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g1_2_0_a2_0_LC_13_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g1_2_0_a2_0_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g1_2_0_a2_0_LC_13_19_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un17_address_g1_2_0_a2_0_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12650),
            .in3(N__13035),
            .lcout(\this_vga_signals.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam G_12_0_x2_0_LC_13_20_0.C_ON=1'b0;
    defparam G_12_0_x2_0_LC_13_20_0.SEQ_MODE=4'b0000;
    defparam G_12_0_x2_0_LC_13_20_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 G_12_0_x2_0_LC_13_20_0 (
            .in0(N__12308),
            .in1(N__12794),
            .in2(_gnd_net_),
            .in3(N__13281),
            .lcout(),
            .ltout(N_6_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNID4564B_LC_13_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNID4564B_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_4_c_RNID4564B_LC_13_20_1 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_4_c_RNID4564B_LC_13_20_1  (
            .in0(N__10592),
            .in1(N__13773),
            .in2(N__10286),
            .in3(N__13552),
            .lcout(\this_vga_signals.N_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_6_LC_13_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_6_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_6_LC_13_20_2 .LUT_INIT=16'b0011011011001001;
    LogicCell40 \this_vga_signals.un17_address_g0_6_LC_13_20_2  (
            .in0(N__10274),
            .in1(N__12795),
            .in2(N__12035),
            .in3(N__13045),
            .lcout(\this_vga_signals.g0_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_6_c_RNIHI8G23_LC_13_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_6_c_RNIHI8G23_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_6_c_RNIHI8G23_LC_13_20_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_6_c_RNIHI8G23_LC_13_20_4  (
            .in0(N__10265),
            .in1(N__12652),
            .in2(_gnd_net_),
            .in3(N__13044),
            .lcout(\this_vga_signals.N_5_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam G_12_0_o7_1_LC_13_20_5.C_ON=1'b0;
    defparam G_12_0_o7_1_LC_13_20_5.SEQ_MODE=4'b0000;
    defparam G_12_0_o7_1_LC_13_20_5.LUT_INIT=16'b0000100101100000;
    LogicCell40 G_12_0_o7_1_LC_13_20_5 (
            .in0(N__12796),
            .in1(N__12309),
            .in2(N__12674),
            .in3(N__13282),
            .lcout(),
            .ltout(N_11_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIPAA128_LC_13_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIPAA128_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNIPAA128_LC_13_20_6 .LUT_INIT=16'b0010000011101100;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_3_c_RNIPAA128_LC_13_20_6  (
            .in0(N__12950),
            .in1(N__13772),
            .in2(N__10595),
            .in3(N__10591),
            .lcout(\this_vga_signals.G_12_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_0_LC_13_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_0_LC_13_21_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vstate_q_0_LC_13_21_0 .LUT_INIT=16'b0000100000001101;
    LogicCell40 \this_vga_signals.M_vstate_q_0_LC_13_21_0  (
            .in0(N__10547),
            .in1(N__10569),
            .in2(N__17727),
            .in3(N__10577),
            .lcout(\this_vga_signals.M_vstate_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17330),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNO_1_1_LC_13_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNO_1_1_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNO_1_1_LC_13_21_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNO_1_1_LC_13_21_7  (
            .in0(N__10568),
            .in1(N__10744),
            .in2(_gnd_net_),
            .in3(N__10546),
            .lcout(\this_vga_signals.N_275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_m16_0_x4_LC_13_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_m16_0_x4_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_m16_0_x4_LC_13_22_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_address_if_m16_0_x4_LC_13_22_3  (
            .in0(N__10741),
            .in1(N__14368),
            .in2(_gnd_net_),
            .in3(N__14300),
            .lcout(),
            .ltout(\this_vga_signals.if_N_9_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_13_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_13_22_4 .LUT_INIT=16'b1010001101011100;
    LogicCell40 \this_vga_signals.un5_address_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_13_22_4  (
            .in0(N__11025),
            .in1(N__10835),
            .in2(N__10463),
            .in3(N__10460),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIO5SOPF2_9_LC_13_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIO5SOPF2_9_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIO5SOPF2_9_LC_13_22_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIO5SOPF2_9_LC_13_22_5  (
            .in0(N__19986),
            .in1(N__11524),
            .in2(N__10454),
            .in3(N__11539),
            .lcout(M_this_vga_signals_address_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_3_0_LC_13_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_3_0_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_3_0_LC_13_23_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNITV8S_3_0_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__10827),
            .in2(_gnd_net_),
            .in3(N__10740),
            .lcout(),
            .ltout(\this_vga_signals.address_m6_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI9MCQB9_0_2_LC_13_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI9MCQB9_0_2_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI9MCQB9_0_2_LC_13_23_1 .LUT_INIT=16'b0000011111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI9MCQB9_0_2_LC_13_23_1  (
            .in0(N__10615),
            .in1(N__11004),
            .in2(N__10343),
            .in3(N__10340),
            .lcout(),
            .ltout(\this_vga_signals.address_i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI2QRE761_0_LC_13_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI2QRE761_0_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI2QRE761_0_LC_13_23_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI2QRE761_0_LC_13_23_2  (
            .in0(N__11046),
            .in1(N__10868),
            .in2(N__11189),
            .in3(N__11186),
            .lcout(),
            .ltout(\this_vga_signals.address_m21_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI7GUI2B2_2_LC_13_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI7GUI2B2_2_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI7GUI2B2_2_LC_13_23_3 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI7GUI2B2_2_LC_13_23_3  (
            .in0(N__10870),
            .in1(N__11180),
            .in2(N__11174),
            .in3(N__11171),
            .lcout(),
            .ltout(\this_vga_signals.address_N_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIH8E9EM_1_LC_13_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIH8E9EM_1_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIH8E9EM_1_LC_13_23_4 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIH8E9EM_1_LC_13_23_4  (
            .in0(N__10917),
            .in1(N__20008),
            .in2(N__11165),
            .in3(N__11162),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_address_if_m16_0_o4_LC_13_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_address_if_m16_0_o4_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_address_if_m16_0_o4_LC_13_23_6 .LUT_INIT=16'b1110100011010100;
    LogicCell40 \this_vga_signals.un5_address_if_m16_0_o4_LC_13_23_6  (
            .in0(N__11047),
            .in1(N__11003),
            .in2(N__10921),
            .in3(N__10869),
            .lcout(\this_vga_signals.if_m16_0_o4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_0_0_LC_13_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_0_0_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNITV8S_0_0_LC_13_24_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNITV8S_0_0_LC_13_24_7  (
            .in0(N__10814),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10745),
            .lcout(\this_vga_signals.address_N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_20_LC_14_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_20_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_20_LC_14_17_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un17_address_g0_20_LC_14_17_0  (
            .in0(N__13082),
            .in1(_gnd_net_),
            .in2(N__12661),
            .in3(N__18355),
            .lcout(\this_vga_signals.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_14_LC_14_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_14_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_14_LC_14_17_2 .LUT_INIT=16'b1111111011001000;
    LogicCell40 \this_vga_signals.un17_address_g0_14_LC_14_17_2  (
            .in0(N__11743),
            .in1(N__12024),
            .in2(N__11870),
            .in3(N__10604),
            .lcout(\this_vga_signals.if_N_8_mux_2_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_3L3_LC_14_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_3L3_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_3L3_LC_14_17_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_3L3_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__12620),
            .in2(N__18361),
            .in3(N__13081),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_3L3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_4L5_LC_14_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_4L5_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_4L5_LC_14_17_4 .LUT_INIT=16'b0111100111110011;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_4L5_LC_14_17_4  (
            .in0(N__13709),
            .in1(N__13448),
            .in2(N__11234),
            .in3(N__12481),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5 ),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_14_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_14_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__11231),
            .in2(N__11219),
            .in3(N__13575),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc5_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_10_i_o2_LC_14_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_10_i_o2_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_10_i_o2_LC_14_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.un17_address_g0_10_i_o2_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__11865),
            .in2(_gnd_net_),
            .in3(N__11742),
            .lcout(\this_vga_signals.N_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_16_0_LC_14_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_16_0_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_16_0_LC_14_18_0 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un17_address_g0_16_0_LC_14_18_0  (
            .in0(N__13478),
            .in1(N__11881),
            .in2(N__13816),
            .in3(N__11678),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_3_LC_14_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_3_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_3_LC_14_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_3_LC_14_18_1  (
            .in0(N__11216),
            .in1(N__13283),
            .in2(N__13488),
            .in3(N__13084),
            .lcout(\this_vga_signals.g0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_9_LC_14_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_9_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_9_LC_14_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un17_address_g0_9_LC_14_18_3  (
            .in0(N__12799),
            .in1(N__12314),
            .in2(_gnd_net_),
            .in3(N__12626),
            .lcout(\this_vga_signals.N_20_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_0_LC_14_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_0_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_0_LC_14_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_0_0_LC_14_18_4  (
            .in0(N__12625),
            .in1(N__12798),
            .in2(N__11210),
            .in3(N__11198),
            .lcout(\this_vga_signals.g0_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_22_LC_14_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_22_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_22_LC_14_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_22_LC_14_18_5  (
            .in0(N__12797),
            .in1(N__12313),
            .in2(N__13823),
            .in3(N__12624),
            .lcout(\this_vga_signals.N_3_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axb3_LC_14_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axb3_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axb3_LC_14_18_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axb3_LC_14_18_6  (
            .in0(N__12627),
            .in1(N__12800),
            .in2(N__13817),
            .in3(N__12316),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_axb3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_ac0_7_0_LC_14_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_ac0_7_0_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_ac0_7_0_LC_14_18_7 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_ac0_7_0_LC_14_18_7  (
            .in0(N__12980),
            .in1(N__12401),
            .in2(N__11192),
            .in3(N__12713),
            .lcout(\this_vga_signals.mult1_un82_sum_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_i_x4_4_a3_LC_14_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_i_x4_4_a3_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_i_x4_4_a3_LC_14_19_0 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_i_x4_4_a3_LC_14_19_0  (
            .in0(N__11375),
            .in1(N__11369),
            .in2(N__11654),
            .in3(N__12041),
            .lcout(\this_vga_signals.g0_i_x4_4_a3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m5_2_LC_14_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m5_2_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m5_2_LC_14_19_1 .LUT_INIT=16'b0111011001100010;
    LogicCell40 \this_vga_signals.un17_address_if_m5_2_LC_14_19_1  (
            .in0(N__11363),
            .in1(N__13463),
            .in2(N__13784),
            .in3(N__11354),
            .lcout(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5),
            .ltout(this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un75_sum_axbxc5_LC_14_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un75_sum_axbxc5_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un75_sum_axbxc5_LC_14_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un75_sum_axbxc5_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__12602),
            .in2(N__11348),
            .in3(N__12298),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m2_2_LC_14_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m2_2_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m2_2_LC_14_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_if_m2_2_LC_14_19_3  (
            .in0(N__12299),
            .in1(N__13271),
            .in2(N__12814),
            .in3(N__12465),
            .lcout(\this_vga_signals.if_N_3_2_i ),
            .ltout(\this_vga_signals.if_N_3_2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_ac0_7_0_1_0_LC_14_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_ac0_7_0_1_0_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_ac0_7_0_1_0_LC_14_19_4 .LUT_INIT=16'b0011000001100110;
    LogicCell40 \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_ac0_7_0_1_0_LC_14_19_4  (
            .in0(N__12466),
            .in1(N__13733),
            .in2(N__11345),
            .in3(N__13574),
            .lcout(\this_vga_signals.mult1_un82_sum_ac0_7_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_2_0_a3_LC_14_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_2_0_a3_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_2_0_a3_LC_14_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_2_0_a3_LC_14_19_5  (
            .in0(N__13464),
            .in1(N__18347),
            .in2(N__13785),
            .in3(N__11676),
            .lcout(\this_vga_signals.g1_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_if_m2_2_0_LC_14_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_if_m2_2_0_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_if_m2_2_0_LC_14_19_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un17_address_if_m2_2_0_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__13729),
            .in2(_gnd_net_),
            .in3(N__12601),
            .lcout(this_vga_signals_un17_address_if_m2_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIP8K884_9_LC_14_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIP8K884_9_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIP8K884_9_LC_14_19_7 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIP8K884_9_LC_14_19_7  (
            .in0(N__12603),
            .in1(N__12317),
            .in2(N__20012),
            .in3(N__12812),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g1_0_0_LC_14_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g1_0_0_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g1_0_0_LC_14_20_0 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \this_vga_signals.un17_address_g1_0_0_LC_14_20_0  (
            .in0(N__13771),
            .in1(N__12660),
            .in2(N__12978),
            .in3(N__13189),
            .lcout(\this_vga_signals.g1_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_0_a2_2_LC_14_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_0_a2_2_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_0_a2_2_LC_14_20_1 .LUT_INIT=16'b0101011010101001;
    LogicCell40 \this_vga_signals.un17_address_g0_0_0_a2_2_LC_14_20_1  (
            .in0(N__13453),
            .in1(N__11869),
            .in2(N__11762),
            .in3(N__12302),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_0_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_12_0_a3_LC_14_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_12_0_a3_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_12_0_a3_LC_14_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_12_0_a3_LC_14_20_2  (
            .in0(N__12790),
            .in1(N__11677),
            .in2(N__11660),
            .in3(N__13278),
            .lcout(),
            .ltout(\this_vga_signals.if_N_3_2_i_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_0_a2_3_LC_14_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_0_a2_3_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_0_a2_3_LC_14_20_3 .LUT_INIT=16'b1000000001000000;
    LogicCell40 \this_vga_signals.un17_address_g0_0_0_a2_3_LC_14_20_3  (
            .in0(N__13769),
            .in1(N__12949),
            .in2(N__11657),
            .in3(N__11645),
            .lcout(\this_vga_signals.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_14_0_a2_i_x2_LC_14_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_14_0_a2_i_x2_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_14_0_a2_i_x2_LC_14_20_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un17_address_g0_14_0_a2_i_x2_LC_14_20_4  (
            .in0(N__12301),
            .in1(_gnd_net_),
            .in2(N__12813),
            .in3(N__12659),
            .lcout(\this_vga_signals.N_20_i_i ),
            .ltout(\this_vga_signals.N_20_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_a3_3_LC_14_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_a3_3_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_a3_3_LC_14_20_5 .LUT_INIT=16'b0100101100101101;
    LogicCell40 \this_vga_signals.un17_address_g0_0_a3_3_LC_14_20_5  (
            .in0(N__13454),
            .in1(N__13770),
            .in2(N__11639),
            .in3(N__11636),
            .lcout(\this_vga_signals.g0_0_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_2_2_LC_14_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_2_2_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_2_2_LC_14_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un17_address_g0_2_2_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__12300),
            .in2(_gnd_net_),
            .in3(N__12786),
            .lcout(\this_vga_signals.N_4_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_12_LC_14_22_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_12_LC_14_22_7 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_12_LC_14_22_7 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \this_vram.mem_radreg_12_LC_14_22_7  (
            .in0(N__19995),
            .in1(N__11627),
            .in2(_gnd_net_),
            .in3(N__11576),
            .lcout(\this_vram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17331),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIL305C61_9_LC_14_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIL305C61_9_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIL305C61_9_LC_14_23_0 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIL305C61_9_LC_14_23_0  (
            .in0(N__11540),
            .in1(N__19993),
            .in2(_gnd_net_),
            .in3(N__11525),
            .lcout(M_this_vga_signals_address_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIR6TCF_9_LC_14_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIR6TCF_9_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIR6TCF_9_LC_14_23_2 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIR6TCF_9_LC_14_23_2  (
            .in0(N__19994),
            .in1(N__11405),
            .in2(_gnd_net_),
            .in3(N__12242),
            .lcout(M_this_vga_signals_address_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_17_LC_15_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_17_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_17_LC_15_17_2 .LUT_INIT=16'b1001011101110111;
    LogicCell40 \this_vga_signals.un17_address_g0_17_LC_15_17_2  (
            .in0(N__13450),
            .in1(N__12107),
            .in2(N__13814),
            .in3(N__12485),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIETEJ4_11_LC_15_17_3 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIETEJ4_11_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIETEJ4_11_LC_15_17_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_radreg_RNIETEJ4_11_LC_15_17_3  (
            .in0(N__16977),
            .in1(N__17830),
            .in2(_gnd_net_),
            .in3(N__16999),
            .lcout(),
            .ltout(\this_vram.M_this_vram_read_data_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI0FV6Q_1_11_LC_15_17_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI0FV6Q_1_11_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI0FV6Q_1_11_LC_15_17_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \this_vram.mem_radreg_RNI0FV6Q_1_11_LC_15_17_4  (
            .in0(N__14141),
            .in1(_gnd_net_),
            .in2(N__12101),
            .in3(N__16952),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_6_0_LC_15_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_6_0_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_6_0_LC_15_17_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_6_0_LC_15_17_7  (
            .in0(N__19825),
            .in1(N__13298),
            .in2(N__12071),
            .in3(N__12815),
            .lcout(\this_vga_signals.g0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_5_0_a2_0_LC_15_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_5_0_a2_0_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_5_0_a2_0_LC_15_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_5_0_a2_0_LC_15_18_0  (
            .in0(N__12059),
            .in1(N__12663),
            .in2(N__13820),
            .in3(N__12808),
            .lcout(),
            .ltout(\this_vga_signals.N_3_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_5_LC_15_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_5_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_5_LC_15_18_1 .LUT_INIT=16'b1110010110000101;
    LogicCell40 \this_vga_signals.un17_address_g0_5_LC_15_18_1  (
            .in0(N__12976),
            .in1(N__14050),
            .in2(N__12050),
            .in3(N__12347),
            .lcout(\this_vga_signals.mult1_un89_sum_c5_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_0_0_LC_15_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_0_0_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_0_0_LC_15_18_2 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \this_vga_signals.un17_address_g0_0_0_0_LC_15_18_2  (
            .in0(N__13555),
            .in1(N__12047),
            .in2(N__13818),
            .in3(N__12710),
            .lcout(\this_vga_signals.g0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_a3_2_LC_15_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_a3_2_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_a3_2_LC_15_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_0_a3_2_LC_15_18_3  (
            .in0(N__12033),
            .in1(N__11882),
            .in2(N__12987),
            .in3(N__13556),
            .lcout(\this_vga_signals.g0_0_a3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_13_LC_15_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_13_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_13_LC_15_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_13_LC_15_18_4  (
            .in0(N__12323),
            .in1(N__12662),
            .in2(N__13819),
            .in3(N__12807),
            .lcout(\this_vga_signals.g0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_LC_15_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_LC_15_18_5 .LUT_INIT=16'b0111111111101111;
    LogicCell40 \this_vga_signals.un17_address_g0_LC_15_18_5  (
            .in0(N__12422),
            .in1(N__13798),
            .in2(N__12988),
            .in3(N__12416),
            .lcout(),
            .ltout(\this_vga_signals.N_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_a3_5_LC_15_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_a3_5_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_a3_5_LC_15_18_6 .LUT_INIT=16'b1001101001100101;
    LogicCell40 \this_vga_signals.un17_address_g0_0_a3_5_LC_15_18_6  (
            .in0(N__12410),
            .in1(N__12400),
            .in2(N__12389),
            .in3(N__12386),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_a3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_a3_LC_15_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_a3_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_a3_LC_15_18_7 .LUT_INIT=16'b1011010000101101;
    LogicCell40 \this_vga_signals.un17_address_g0_0_a3_LC_15_18_7  (
            .in0(N__12975),
            .in1(N__14051),
            .in2(N__12380),
            .in3(N__12377),
            .lcout(\this_vga_signals.mult1_un96_sum_axbxc5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_29_LC_15_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_29_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_29_LC_15_19_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vga_signals.un17_address_g0_29_LC_15_19_0  (
            .in0(N__12957),
            .in1(N__12371),
            .in2(_gnd_net_),
            .in3(N__13135),
            .lcout(),
            .ltout(\this_vga_signals.g1_5_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_27_LC_15_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_27_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_27_LC_15_19_1 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_27_LC_15_19_1  (
            .in0(N__12365),
            .in1(N__12356),
            .in2(N__12350),
            .in3(N__12842),
            .lcout(\this_vga_signals.r_N_2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_1_2_LC_15_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_1_2_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_1_2_LC_15_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_1_2_LC_15_19_2  (
            .in0(N__12318),
            .in1(N__12671),
            .in2(N__12341),
            .in3(N__13076),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_12_LC_15_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_12_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_12_LC_15_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un17_address_g0_12_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__13279),
            .in2(N__12326),
            .in3(N__12801),
            .lcout(\this_vga_signals.if_N_3_2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_3_0_a2_1_LC_15_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_3_0_a2_1_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_3_0_a2_1_LC_15_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_3_0_a2_1_LC_15_19_4  (
            .in0(N__12319),
            .in1(N__18356),
            .in2(N__13489),
            .in3(N__13077),
            .lcout(),
            .ltout(\this_vga_signals.g0_3_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_3_0_a2_LC_15_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_3_0_a2_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_3_0_a2_LC_15_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_3_0_a2_LC_15_19_5  (
            .in0(N__12672),
            .in1(N__13280),
            .in2(N__12845),
            .in3(N__12802),
            .lcout(\this_vga_signals.if_N_3_2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_23_LC_15_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_23_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_23_LC_15_19_6 .LUT_INIT=16'b0101011000000110;
    LogicCell40 \this_vga_signals.un17_address_g0_23_LC_15_19_6  (
            .in0(N__13813),
            .in1(N__12482),
            .in2(N__13576),
            .in3(N__12711),
            .lcout(\this_vga_signals.mult1_un82_sum_ac0_7_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_5_0_a2_LC_15_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_5_0_a2_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_5_0_a2_LC_15_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_5_0_a2_LC_15_19_7  (
            .in0(N__12673),
            .in1(N__12836),
            .in2(N__13822),
            .in3(N__12803),
            .lcout(\this_vga_signals.N_3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_37_LC_15_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_37_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_37_LC_15_20_1 .LUT_INIT=16'b0101011000000110;
    LogicCell40 \this_vga_signals.un17_address_g0_37_LC_15_20_1  (
            .in0(N__13774),
            .in1(N__12483),
            .in2(N__13577),
            .in3(N__12712),
            .lcout(\this_vga_signals.mult1_un82_sum_ac0_7_0_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_5_c_RNI8HPEH2_LC_15_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_5_c_RNI8HPEH2_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_5_c_RNI8HPEH2_LC_15_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_5_c_RNI8HPEH2_LC_15_20_2  (
            .in0(N__12689),
            .in1(N__13287),
            .in2(N__13490),
            .in3(N__12676),
            .lcout(),
            .ltout(\this_vga_signals.g1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_5_c_RNICKLJPG_LC_15_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_5_c_RNICKLJPG_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_5_c_RNICKLJPG_LC_15_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_5_c_RNICKLJPG_LC_15_20_3  (
            .in0(N__13564),
            .in1(N__12509),
            .in2(N__12500),
            .in3(N__12497),
            .lcout(),
            .ltout(\this_vga_signals.g1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNI5J0QQK_LC_15_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNI5J0QQK_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNI5J0QQK_LC_15_20_4 .LUT_INIT=16'b0100101111010010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_3_c_RNI5J0QQK_LC_15_20_4  (
            .in0(N__12979),
            .in1(N__13776),
            .in2(N__12488),
            .in3(N__13565),
            .lcout(\this_vga_signals.g1_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_36_LC_15_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_36_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_36_LC_15_20_5 .LUT_INIT=16'b1001011100111111;
    LogicCell40 \this_vga_signals.un17_address_g0_36_LC_15_20_5  (
            .in0(N__13775),
            .in1(N__13482),
            .in2(N__13211),
            .in3(N__12484),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_3_LC_15_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_3_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_3_LC_15_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un17_address_g0_0_3_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__12434),
            .in2(N__12425),
            .in3(N__13563),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_33_LC_15_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_33_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_33_LC_15_20_7 .LUT_INIT=16'b0000111101111000;
    LogicCell40 \this_vga_signals.un17_address_g0_33_LC_15_20_7  (
            .in0(N__13175),
            .in1(N__13163),
            .in2(N__13157),
            .in3(N__13154),
            .lcout(\this_vga_signals.N_3_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_5_0_LC_16_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_5_0_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_5_0_LC_16_17_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un17_address_g0_5_0_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__13777),
            .in2(_gnd_net_),
            .in3(N__13447),
            .lcout(\this_vga_signals.g0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_7_LC_16_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_7_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_7_LC_16_18_2 .LUT_INIT=16'b0011100110011100;
    LogicCell40 \this_vga_signals.un17_address_g0_7_LC_16_18_2  (
            .in0(N__13815),
            .in1(N__13148),
            .in2(N__12989),
            .in3(N__13583),
            .lcout(\this_vga_signals.g0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g1_4_LC_16_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g1_4_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g1_4_LC_16_18_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vga_signals.un17_address_g1_4_LC_16_18_5  (
            .in0(N__12981),
            .in1(N__13142),
            .in2(_gnd_net_),
            .in3(N__13136),
            .lcout(),
            .ltout(\this_vga_signals.g1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_0_0_a2_LC_16_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_0_0_a2_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_0_0_a2_LC_16_18_6 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_0_0_a2_LC_16_18_6  (
            .in0(N__13124),
            .in1(N__13115),
            .in2(N__13109),
            .in3(N__13496),
            .lcout(),
            .ltout(\this_vga_signals.r_N_2_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_10_LC_16_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_10_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_10_LC_16_18_7 .LUT_INIT=16'b1110100000110011;
    LogicCell40 \this_vga_signals.un17_address_g0_10_LC_16_18_7  (
            .in0(N__14049),
            .in1(N__12986),
            .in2(N__13106),
            .in3(N__13103),
            .lcout(\this_vga_signals.mult1_un89_sum_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_5_3_LC_16_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_5_3_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_5_3_LC_16_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_5_3_LC_16_19_1  (
            .in0(N__18357),
            .in1(N__13299),
            .in2(N__13097),
            .in3(N__13085),
            .lcout(),
            .ltout(\this_vga_signals.g0_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_34_LC_16_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_34_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_34_LC_16_19_2 .LUT_INIT=16'b0010110110110100;
    LogicCell40 \this_vga_signals.un17_address_g0_34_LC_16_19_2  (
            .in0(N__13806),
            .in1(N__12982),
            .in2(N__12848),
            .in3(N__13579),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un96_sum_c5_0_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_32_LC_16_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_32_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_32_LC_16_19_3 .LUT_INIT=16'b0101010111101000;
    LogicCell40 \this_vga_signals.un17_address_g0_32_LC_16_19_3  (
            .in0(N__14048),
            .in1(N__14008),
            .in2(N__13991),
            .in3(N__13988),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un96_sum_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNI7M4QI33_LC_16_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNI7M4QI33_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un12_address_un12_address_cry_3_c_RNI7M4QI33_LC_16_19_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un12_address_un12_address_cry_3_c_RNI7M4QI33_LC_16_19_4  (
            .in0(N__13982),
            .in1(_gnd_net_),
            .in2(N__13976),
            .in3(N__13973),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIHKRBFB2_9_LC_16_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIHKRBFB2_9_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIHKRBFB2_9_LC_16_19_5 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIHKRBFB2_9_LC_16_19_5  (
            .in0(N__13964),
            .in1(N__19999),
            .in2(N__13958),
            .in3(N__13955),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_24_LC_16_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_24_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_24_LC_16_19_6 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \this_vga_signals.un17_address_g0_24_LC_16_19_6  (
            .in0(N__13841),
            .in1(N__13829),
            .in2(N__13821),
            .in3(N__13578),
            .lcout(\this_vga_signals.mult1_un82_sum_ac0_7_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un17_address_g0_35_LC_16_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un17_address_g0_35_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un17_address_g0_35_LC_16_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un17_address_g0_35_LC_16_20_3  (
            .in0(N__13487),
            .in1(N__13301),
            .in2(N__13210),
            .in3(N__13190),
            .lcout(\this_vga_signals.if_N_3_2_i_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_1_LC_16_20_4 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_1_LC_16_20_4 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_1_LC_16_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_1_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13169),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17312),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_0_LC_16_20_7 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_0_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_0_LC_16_20_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_0_LC_16_20_7  (
            .in0(N__14122),
            .in1(N__16887),
            .in2(_gnd_net_),
            .in3(N__14105),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17312),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_1_LC_16_21_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_1_LC_16_21_0 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_1_LC_16_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_1_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14093),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17315),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_last_q_LC_16_21_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_last_q_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_edge_detector.M_last_q_LC_16_21_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_last_q_LC_16_21_1  (
            .in0(N__14132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16895),
            .lcout(this_start_data_delay_this_edge_detector_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17315),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_0_LC_16_21_7 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_0_LC_16_21_7 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_0_LC_16_21_7 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_0_LC_16_21_7  (
            .in0(N__14131),
            .in1(N__16894),
            .in2(_gnd_net_),
            .in3(N__14104),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17315),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_4_LC_16_22_2 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_4_LC_16_22_2 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_4_LC_16_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_4_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14087),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17317),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_3_LC_16_22_4 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_3_LC_16_22_4 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_3_LC_16_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_3_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14075),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17317),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_2_LC_16_22_5 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_2_LC_16_22_5 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_2_LC_16_22_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_2_LC_16_22_5  (
            .in0(_gnd_net_),
            .in1(N__14081),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17317),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_6_LC_17_20_0 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_6_LC_17_20_0 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_6_LC_17_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_6_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14069),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17316),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_5_LC_17_20_1 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_5_LC_17_20_1 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_5_LC_17_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_5_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14405),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17316),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_3_LC_17_20_2 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_3_LC_17_20_2 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_3_LC_17_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_3_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14057),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17316),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_2_LC_17_20_5 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_2_LC_17_20_5 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_2_LC_17_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_2_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14063),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17316),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_4_LC_17_20_7 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_4_LC_17_20_7 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_4_LC_17_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_4_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14411),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17316),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_10_LC_17_21_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_10_LC_17_21_0 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_10_LC_17_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_10_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14393),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17319),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_11_LC_17_21_3 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_11_LC_17_21_3 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_11_LC_17_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_11_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14399),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17319),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_9_LC_17_22_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_9_LC_17_22_0 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_9_LC_17_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_9_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14540),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17326),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_6_LC_17_22_2 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_6_LC_17_22_2 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_6_LC_17_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_6_LC_17_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14375),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17326),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_7_LC_17_22_3 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_7_LC_17_22_3 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_7_LC_17_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_7_LC_17_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14387),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17326),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_5_LC_17_22_5 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_5_LC_17_22_5 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_5_LC_17_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_5_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14381),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17326),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIOUPCH9_9_LC_17_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIOUPCH9_9_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIOUPCH9_9_LC_17_23_1 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIOUPCH9_9_LC_17_23_1  (
            .in0(N__20019),
            .in1(N__14369),
            .in2(_gnd_net_),
            .in3(N__14299),
            .lcout(M_this_vga_signals_address_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIETEJ4_0_11_LC_18_17_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIETEJ4_0_11_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIETEJ4_0_11_LC_18_17_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_radreg_RNIETEJ4_0_11_LC_18_17_4  (
            .in0(N__18716),
            .in1(N__17841),
            .in2(_gnd_net_),
            .in3(N__18079),
            .lcout(\this_vram.M_this_vram_read_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIIHGJL_11_LC_18_18_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIIHGJL_11_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIIHGJL_11_LC_18_18_7 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \this_vram.mem_radreg_RNIIHGJL_11_LC_18_18_7  (
            .in0(N__18080),
            .in1(N__17837),
            .in2(N__16951),
            .in3(N__18709),
            .lcout(\this_vram.N_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_12_LC_18_20_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_12_LC_18_20_1 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_12_LC_18_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_12_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14465),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17320),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_13_LC_18_20_2 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_13_LC_18_20_2 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_13_LC_18_20_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_13_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__14459),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17320),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_state_q_s2_0_a3_LC_18_20_6 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_s2_0_a3_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_state_q_s2_0_a3_LC_18_20_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_state_q_s2_0_a3_LC_18_20_6  (
            .in0(N__17503),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16355),
            .lcout(debug_d),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_16_LC_18_21_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_16_LC_18_21_0 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_16_LC_18_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_16_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14423),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17327),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_14_LC_18_21_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_14_LC_18_21_1 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_14_LC_18_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_14_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14435),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17327),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_15_LC_18_21_2 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_15_LC_18_21_2 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_15_LC_18_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_15_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14429),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17327),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_5_LC_18_21_6 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_5_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_5_LC_18_21_6 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_5_LC_18_21_6  (
            .in0(N__14949),
            .in1(N__17567),
            .in2(N__14753),
            .in3(N__16339),
            .lcout(\this_start_data_delay.this_edge_detector.N_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_17_LC_18_22_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_17_LC_18_22_0 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_17_LC_18_22_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_17_LC_18_22_0  (
            .in0(N__14417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17332),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_19_LC_18_22_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_19_LC_18_22_1 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_19_LC_18_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_19_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14552),
            .lcout(M_this_start_data_delay_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17332),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_18_LC_18_22_2 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_18_LC_18_22_2 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_18_LC_18_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_18_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14558),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17332),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_delay.M_pipe_q_8_LC_18_22_6 .C_ON=1'b0;
    defparam \this_start_data_delay.this_delay.M_pipe_q_8_LC_18_22_6 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.this_delay.M_pipe_q_8_LC_18_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_data_delay.this_delay.M_pipe_q_8_LC_18_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14546),
            .lcout(\this_start_data_delay.this_delay.M_pipe_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17332),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_2_LC_18_23_1.C_ON=1'b0;
    defparam M_current_address_q_2_LC_18_23_1.SEQ_MODE=4'b1000;
    defparam M_current_address_q_2_LC_18_23_1.LUT_INIT=16'b1101100011100100;
    LogicCell40 M_current_address_q_2_LC_18_23_1 (
            .in0(N__16343),
            .in1(N__14567),
            .in2(N__14522),
            .in3(N__17500),
            .lcout(M_current_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17338),
            .ce(),
            .sr(N__15464));
    defparam M_current_address_q_5_LC_18_23_6.C_ON=1'b0;
    defparam M_current_address_q_5_LC_18_23_6.SEQ_MODE=4'b1000;
    defparam M_current_address_q_5_LC_18_23_6.LUT_INIT=16'b1101100011100100;
    LogicCell40 M_current_address_q_5_LC_18_23_6 (
            .in0(N__17499),
            .in1(N__14924),
            .in2(N__14534),
            .in3(N__16344),
            .lcout(M_current_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17338),
            .ce(),
            .sr(N__15464));
    defparam M_current_address_q_9_LC_18_24_2.C_ON=1'b0;
    defparam M_current_address_q_9_LC_18_24_2.SEQ_MODE=4'b1000;
    defparam M_current_address_q_9_LC_18_24_2.LUT_INIT=16'b1011100011100010;
    LogicCell40 M_current_address_q_9_LC_18_24_2 (
            .in0(N__14774),
            .in1(N__17486),
            .in2(N__14510),
            .in3(N__16342),
            .lcout(M_current_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17342),
            .ce(),
            .sr(N__15462));
    defparam M_current_address_q_8_LC_18_24_3.C_ON=1'b0;
    defparam M_current_address_q_8_LC_18_24_3.SEQ_MODE=4'b1000;
    defparam M_current_address_q_8_LC_18_24_3.LUT_INIT=16'b1110110101001000;
    LogicCell40 M_current_address_q_8_LC_18_24_3 (
            .in0(N__16341),
            .in1(N__16022),
            .in2(N__17501),
            .in3(N__14909),
            .lcout(M_current_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17342),
            .ce(),
            .sr(N__15462));
    defparam M_current_address_q_4_LC_18_24_4.C_ON=1'b0;
    defparam M_current_address_q_4_LC_18_24_4.SEQ_MODE=4'b1000;
    defparam M_current_address_q_4_LC_18_24_4.LUT_INIT=16'b1011100011100010;
    LogicCell40 M_current_address_q_4_LC_18_24_4 (
            .in0(N__15059),
            .in1(N__17485),
            .in2(N__16370),
            .in3(N__16340),
            .lcout(M_current_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17342),
            .ce(),
            .sr(N__15462));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_2_LC_18_25_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_2_LC_18_25_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_2_LC_18_25_1 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_2_LC_18_25_1  (
            .in0(N__14593),
            .in1(N__17604),
            .in2(N__19036),
            .in3(N__16333),
            .lcout(\this_start_data_delay.this_edge_detector.N_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_9_LC_18_25_3 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_9_LC_18_25_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_9_LC_18_25_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_9_LC_18_25_3  (
            .in0(N__14800),
            .in1(N__17605),
            .in2(N__19037),
            .in3(N__16334),
            .lcout(\this_start_data_delay.this_edge_detector.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_12_LC_19_20_3.C_ON=1'b0;
    defparam M_current_address_q_12_LC_19_20_3.SEQ_MODE=4'b1000;
    defparam M_current_address_q_12_LC_19_20_3.LUT_INIT=16'b1011100011100010;
    LogicCell40 M_current_address_q_12_LC_19_20_3 (
            .in0(N__15131),
            .in1(N__17502),
            .in2(N__14723),
            .in3(N__16351),
            .lcout(M_current_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17328),
            .ce(),
            .sr(N__15466));
    defparam \this_start_address_delay.this_delay.M_pipe_q_9_LC_19_21_1 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_9_LC_19_21_1 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_9_LC_19_21_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_9_LC_19_21_1  (
            .in0(N__14759),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17333),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_8_LC_19_21_3 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_8_LC_19_21_3 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_8_LC_19_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_8_LC_19_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14702),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17333),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_12_LC_19_21_4 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_12_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_12_LC_19_21_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_12_LC_19_21_4  (
            .in0(N__19273),
            .in1(N__17568),
            .in2(N__14752),
            .in3(N__16338),
            .lcout(\this_start_data_delay.this_edge_detector.N_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_7_LC_19_21_5 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_7_LC_19_21_5 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_7_LC_19_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_7_LC_19_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14714),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17333),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_10_LC_19_21_7 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_10_LC_19_21_7 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_10_LC_19_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_10_LC_19_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14696),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17333),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_RNIHDTU_0_LC_19_23_0.C_ON=1'b1;
    defparam M_current_address_q_RNIHDTU_0_LC_19_23_0.SEQ_MODE=4'b0000;
    defparam M_current_address_q_RNIHDTU_0_LC_19_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_current_address_q_RNIHDTU_0_LC_19_23_0 (
            .in0(_gnd_net_),
            .in1(N__15583),
            .in2(N__15116),
            .in3(N__15115),
            .lcout(M_current_address_q_RNIHDTUZ0Z_0),
            .ltout(),
            .carryin(bfn_19_23_0_),
            .carryout(un1_M_current_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_0_c_RNI2QAN_LC_19_23_1.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_0_c_RNI2QAN_LC_19_23_1.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_0_c_RNI2QAN_LC_19_23_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_0_c_RNI2QAN_LC_19_23_1 (
            .in0(_gnd_net_),
            .in1(N__16567),
            .in2(_gnd_net_),
            .in3(N__14690),
            .lcout(un1_M_current_address_q_cry_0_c_RNI2QANZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_0),
            .carryout(un1_M_current_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_1_c_RNI4TBN_LC_19_23_2.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_1_c_RNI4TBN_LC_19_23_2.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_1_c_RNI4TBN_LC_19_23_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_1_c_RNI4TBN_LC_19_23_2 (
            .in0(_gnd_net_),
            .in1(N__14589),
            .in2(_gnd_net_),
            .in3(N__14561),
            .lcout(un1_M_current_address_q_cry_1_c_RNI4TBNZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_1),
            .carryout(un1_M_current_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_2_c_RNI60DN_LC_19_23_3.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_2_c_RNI60DN_LC_19_23_3.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_2_c_RNI60DN_LC_19_23_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_2_c_RNI60DN_LC_19_23_3 (
            .in0(_gnd_net_),
            .in1(N__15160),
            .in2(_gnd_net_),
            .in3(N__15062),
            .lcout(un1_M_current_address_q_cry_2_c_RNI60DNZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_2),
            .carryout(un1_M_current_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_3_c_RNI83EN_LC_19_23_4.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_3_c_RNI83EN_LC_19_23_4.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_3_c_RNI83EN_LC_19_23_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_3_c_RNI83EN_LC_19_23_4 (
            .in0(_gnd_net_),
            .in1(N__16422),
            .in2(_gnd_net_),
            .in3(N__15053),
            .lcout(un1_M_current_address_q_cry_3_c_RNI83ENZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_3),
            .carryout(un1_M_current_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_4_c_RNIA6FN_LC_19_23_5.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_4_c_RNIA6FN_LC_19_23_5.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_4_c_RNIA6FN_LC_19_23_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_4_c_RNIA6FN_LC_19_23_5 (
            .in0(_gnd_net_),
            .in1(N__14950),
            .in2(_gnd_net_),
            .in3(N__14918),
            .lcout(un1_M_current_address_q_cry_4_c_RNIA6FNZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_4),
            .carryout(un1_M_current_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_5_c_RNIC9GN_LC_19_23_6.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_5_c_RNIC9GN_LC_19_23_6.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_5_c_RNIC9GN_LC_19_23_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_5_c_RNIC9GN_LC_19_23_6 (
            .in0(_gnd_net_),
            .in1(N__15289),
            .in2(_gnd_net_),
            .in3(N__14915),
            .lcout(un1_M_current_address_q_cry_5_c_RNIC9GNZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_5),
            .carryout(un1_M_current_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_6_c_RNIECHN_LC_19_23_7.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_6_c_RNIECHN_LC_19_23_7.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_6_c_RNIECHN_LC_19_23_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_6_c_RNIECHN_LC_19_23_7 (
            .in0(_gnd_net_),
            .in1(N__15714),
            .in2(_gnd_net_),
            .in3(N__14912),
            .lcout(un1_M_current_address_q_cry_6_c_RNIECHNZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_6),
            .carryout(un1_M_current_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_7_c_RNIGFIN_LC_19_24_0.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_7_c_RNIGFIN_LC_19_24_0.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_7_c_RNIGFIN_LC_19_24_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_7_c_RNIGFIN_LC_19_24_0 (
            .in0(_gnd_net_),
            .in1(N__16041),
            .in2(_gnd_net_),
            .in3(N__14903),
            .lcout(un1_M_current_address_q_cry_7_c_RNIGFINZ0),
            .ltout(),
            .carryin(bfn_19_24_0_),
            .carryout(un1_M_current_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_8_c_RNIIIJN_LC_19_24_1.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_8_c_RNIIIJN_LC_19_24_1.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_8_c_RNIIIJN_LC_19_24_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_8_c_RNIIIJN_LC_19_24_1 (
            .in0(_gnd_net_),
            .in1(N__14799),
            .in2(_gnd_net_),
            .in3(N__14768),
            .lcout(un1_M_current_address_q_cry_8_c_RNIIIJNZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_8),
            .carryout(un1_M_current_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_9_c_RNIRDIM_LC_19_24_2.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_9_c_RNIRDIM_LC_19_24_2.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_9_c_RNIRDIM_LC_19_24_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_9_c_RNIRDIM_LC_19_24_2 (
            .in0(_gnd_net_),
            .in1(N__15909),
            .in2(_gnd_net_),
            .in3(N__14765),
            .lcout(un1_M_current_address_q_cry_9_c_RNIRDIMZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_9),
            .carryout(un1_M_current_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_10_c_RNI4KKH_LC_19_24_3.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_10_c_RNI4KKH_LC_19_24_3.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_10_c_RNI4KKH_LC_19_24_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_10_c_RNI4KKH_LC_19_24_3 (
            .in0(_gnd_net_),
            .in1(N__19185),
            .in2(_gnd_net_),
            .in3(N__14762),
            .lcout(un1_M_current_address_q_cry_10_c_RNI4KKHZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_10),
            .carryout(un1_M_current_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_11_c_RNI6NLH_LC_19_24_4.C_ON=1'b1;
    defparam un1_M_current_address_q_cry_11_c_RNI6NLH_LC_19_24_4.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_11_c_RNI6NLH_LC_19_24_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_current_address_q_cry_11_c_RNI6NLH_LC_19_24_4 (
            .in0(_gnd_net_),
            .in1(N__19286),
            .in2(_gnd_net_),
            .in3(N__15122),
            .lcout(un1_M_current_address_q_cry_11_c_RNI6NLHZ0),
            .ltout(),
            .carryin(un1_M_current_address_q_cry_11),
            .carryout(un1_M_current_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_current_address_q_cry_12_c_RNI8QMH_LC_19_24_5.C_ON=1'b0;
    defparam un1_M_current_address_q_cry_12_c_RNI8QMH_LC_19_24_5.SEQ_MODE=4'b0000;
    defparam un1_M_current_address_q_cry_12_c_RNI8QMH_LC_19_24_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 un1_M_current_address_q_cry_12_c_RNI8QMH_LC_19_24_5 (
            .in0(N__19082),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15119),
            .lcout(un1_M_current_address_q_cry_12_c_RNI8QMHZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.un1_M_state_q_1_i_LC_19_24_6 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.un1_M_state_q_1_i_LC_19_24_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.un1_M_state_q_1_i_LC_19_24_6 .LUT_INIT=16'b1011101111001100;
    LogicCell40 \this_start_data_delay.this_edge_detector.un1_M_state_q_1_i_LC_19_24_6  (
            .in0(N__17608),
            .in1(N__17484),
            .in2(_gnd_net_),
            .in3(N__16296),
            .lcout(N_177_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_10_LC_19_25_1.C_ON=1'b0;
    defparam M_current_address_q_10_LC_19_25_1.SEQ_MODE=4'b1000;
    defparam M_current_address_q_10_LC_19_25_1.LUT_INIT=16'b1011100011100010;
    LogicCell40 M_current_address_q_10_LC_19_25_1 (
            .in0(N__15101),
            .in1(N__17481),
            .in2(N__15890),
            .in3(N__16335),
            .lcout(M_current_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17354),
            .ce(),
            .sr(N__15463));
    defparam M_current_address_q_1_LC_19_25_2.C_ON=1'b0;
    defparam M_current_address_q_1_LC_19_25_2.SEQ_MODE=4'b1000;
    defparam M_current_address_q_1_LC_19_25_2.LUT_INIT=16'b1101100011100100;
    LogicCell40 M_current_address_q_1_LC_19_25_2 (
            .in0(N__16337),
            .in1(N__15095),
            .in2(N__16541),
            .in3(N__17483),
            .lcout(M_current_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17354),
            .ce(),
            .sr(N__15463));
    defparam M_current_address_q_13_LC_19_25_4.C_ON=1'b0;
    defparam M_current_address_q_13_LC_19_25_4.SEQ_MODE=4'b1000;
    defparam M_current_address_q_13_LC_19_25_4.LUT_INIT=16'b1111100101100000;
    LogicCell40 M_current_address_q_13_LC_19_25_4 (
            .in0(N__16336),
            .in1(N__17482),
            .in2(N__15842),
            .in3(N__15086),
            .lcout(M_current_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17354),
            .ce(),
            .sr(N__15463));
    defparam \this_start_address_delay.this_delay.M_pipe_q_13_LC_20_21_1 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_13_LC_20_21_1 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_13_LC_20_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_13_LC_20_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15080),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17339),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_12_LC_20_21_3 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_12_LC_20_21_3 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_12_LC_20_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_12_LC_20_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15068),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17339),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_11_LC_20_21_5 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_11_LC_20_21_5 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_11_LC_20_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_11_LC_20_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15074),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17339),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_15_LC_20_22_0 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_15_LC_20_22_0 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_15_LC_20_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_15_LC_20_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15548),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17343),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_14_LC_20_22_4 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_14_LC_20_22_4 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_14_LC_20_22_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_14_LC_20_22_4  (
            .in0(_gnd_net_),
            .in1(N__15554),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17343),
            .ce(),
            .sr(_gnd_net_));
    defparam M_current_address_q_0_LC_20_23_0.C_ON=1'b0;
    defparam M_current_address_q_0_LC_20_23_0.SEQ_MODE=4'b1000;
    defparam M_current_address_q_0_LC_20_23_0.LUT_INIT=16'b1101100011100100;
    LogicCell40 M_current_address_q_0_LC_20_23_0 (
            .in0(N__17477),
            .in1(N__15542),
            .in2(N__15563),
            .in3(N__16291),
            .lcout(M_current_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17349),
            .ce(),
            .sr(N__15465));
    defparam M_current_address_q_6_LC_20_23_1.C_ON=1'b0;
    defparam M_current_address_q_6_LC_20_23_1.SEQ_MODE=4'b1000;
    defparam M_current_address_q_6_LC_20_23_1.LUT_INIT=16'b1110110101001000;
    LogicCell40 M_current_address_q_6_LC_20_23_1 (
            .in0(N__16294),
            .in1(N__15269),
            .in2(N__17504),
            .in3(N__15536),
            .lcout(M_current_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17349),
            .ce(),
            .sr(N__15465));
    defparam M_current_address_q_7_LC_20_23_3.C_ON=1'b0;
    defparam M_current_address_q_7_LC_20_23_3.SEQ_MODE=4'b1000;
    defparam M_current_address_q_7_LC_20_23_3.LUT_INIT=16'b1101100011100100;
    LogicCell40 M_current_address_q_7_LC_20_23_3 (
            .in0(N__16295),
            .in1(N__15530),
            .in2(N__15695),
            .in3(N__17480),
            .lcout(M_current_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17349),
            .ce(),
            .sr(N__15465));
    defparam M_current_address_q_11_LC_20_23_4.C_ON=1'b0;
    defparam M_current_address_q_11_LC_20_23_4.SEQ_MODE=4'b1000;
    defparam M_current_address_q_11_LC_20_23_4.LUT_INIT=16'b1101100011100100;
    LogicCell40 M_current_address_q_11_LC_20_23_4 (
            .in0(N__17478),
            .in1(N__15524),
            .in2(N__15881),
            .in3(N__16292),
            .lcout(M_current_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17349),
            .ce(),
            .sr(N__15465));
    defparam M_current_address_q_3_LC_20_23_7.C_ON=1'b0;
    defparam M_current_address_q_3_LC_20_23_7.SEQ_MODE=4'b1000;
    defparam M_current_address_q_3_LC_20_23_7.LUT_INIT=16'b1101100011100100;
    LogicCell40 M_current_address_q_3_LC_20_23_7 (
            .in0(N__16293),
            .in1(N__15518),
            .in2(N__15140),
            .in3(N__17479),
            .lcout(M_current_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17349),
            .ce(),
            .sr(N__15465));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_6_LC_20_24_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_6_LC_20_24_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_6_LC_20_24_0 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_6_LC_20_24_0  (
            .in0(N__15288),
            .in1(N__17613),
            .in2(N__15869),
            .in3(N__16285),
            .lcout(\this_start_data_delay.this_edge_detector.N_216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_3_LC_20_24_6 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_3_LC_20_24_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_3_LC_20_24_6 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_3_LC_20_24_6  (
            .in0(N__15159),
            .in1(N__17614),
            .in2(N__20372),
            .in3(N__16284),
            .lcout(\this_start_data_delay.this_edge_detector.N_213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_8_LC_20_24_7 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_8_LC_20_24_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_8_LC_20_24_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_8_LC_20_24_7  (
            .in0(N__16286),
            .in1(N__16045),
            .in2(N__16835),
            .in3(N__17612),
            .lcout(\this_start_data_delay.this_edge_detector.N_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_10_LC_20_25_4 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_10_LC_20_25_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_10_LC_20_25_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_10_LC_20_25_4  (
            .in0(N__15913),
            .in1(N__17619),
            .in2(N__20368),
            .in3(N__16287),
            .lcout(\this_start_data_delay.this_edge_detector.N_220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_11_LC_20_25_5 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_11_LC_20_25_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_11_LC_20_25_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_11_LC_20_25_5  (
            .in0(N__16288),
            .in1(N__16406),
            .in2(N__17626),
            .in3(N__19203),
            .lcout(\this_start_data_delay.this_edge_detector.N_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_13_LC_20_25_7 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_13_LC_20_25_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_13_LC_20_25_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_13_LC_20_25_7  (
            .in0(N__16289),
            .in1(N__15868),
            .in2(N__17627),
            .in3(N__19081),
            .lcout(\this_start_data_delay.this_edge_detector.N_223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_17_LC_21_22_1 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_17_LC_21_22_1 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_17_LC_21_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_17_LC_21_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15827),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17350),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_en_0_sqmuxa_0_a3_LC_21_22_2 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_en_0_sqmuxa_0_a3_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_en_0_sqmuxa_0_a3_LC_21_22_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_this_vram_write_en_0_sqmuxa_0_a3_LC_21_22_2  (
            .in0(N__17569),
            .in1(N__17453),
            .in2(_gnd_net_),
            .in3(N__16332),
            .lcout(M_this_vram_write_en_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_16_LC_21_22_5 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_16_LC_21_22_5 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_16_LC_21_22_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_16_LC_21_22_5  (
            .in0(_gnd_net_),
            .in1(N__15833),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17350),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_7_LC_21_23_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_7_LC_21_23_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_7_LC_21_23_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_7_LC_21_23_0  (
            .in0(N__16280),
            .in1(N__17624),
            .in2(N__15721),
            .in3(N__17140),
            .lcout(\this_start_data_delay.this_edge_detector.N_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_0_LC_21_23_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_0_LC_21_23_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_0_LC_21_23_1 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_0_LC_21_23_1  (
            .in0(N__17623),
            .in1(N__15582),
            .in2(N__17141),
            .in3(N__16279),
            .lcout(\this_start_data_delay.this_edge_detector.N_210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_18_LC_21_24_2 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_18_LC_21_24_2 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_18_LC_21_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_18_LC_21_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16688),
            .lcout(\this_start_address_delay.this_delay.M_pipe_qZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17361),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.this_delay.M_pipe_q_19_LC_21_24_3 .C_ON=1'b0;
    defparam \this_start_address_delay.this_delay.M_pipe_q_19_LC_21_24_3 .SEQ_MODE=4'b1000;
    defparam \this_start_address_delay.this_delay.M_pipe_q_19_LC_21_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_start_address_delay.this_delay.M_pipe_q_19_LC_21_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16679),
            .lcout(M_this_start_address_delay_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17361),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_ns_1_0__m7_LC_21_24_5.C_ON=1'b0;
    defparam M_state_q_ns_1_0__m7_LC_21_24_5.SEQ_MODE=4'b0000;
    defparam M_state_q_ns_1_0__m7_LC_21_24_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 M_state_q_ns_1_0__m7_LC_21_24_5 (
            .in0(N__19661),
            .in1(N__16841),
            .in2(_gnd_net_),
            .in3(N__16673),
            .lcout(M_state_q_ns_1_0__N_24_mux),
            .ltout(M_state_q_ns_1_0__N_24_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_ns_1_0__m9_LC_21_24_6.C_ON=1'b0;
    defparam M_state_q_ns_1_0__m9_LC_21_24_6.SEQ_MODE=4'b0000;
    defparam M_state_q_ns_1_0__m9_LC_21_24_6.LUT_INIT=16'b0000000001010000;
    LogicCell40 M_state_q_ns_1_0__m9_LC_21_24_6 (
            .in0(N__16169),
            .in1(_gnd_net_),
            .in2(N__16667),
            .in3(N__17451),
            .lcout(),
            .ltout(M_state_q_ns_1_0__N_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_0_LC_21_24_7.C_ON=1'b0;
    defparam M_state_q_0_LC_21_24_7.SEQ_MODE=4'b1000;
    defparam M_state_q_0_LC_21_24_7.LUT_INIT=16'b0001000101010000;
    LogicCell40 M_state_q_0_LC_21_24_7 (
            .in0(N__17740),
            .in1(N__17615),
            .in2(N__16664),
            .in3(N__16290),
            .lcout(M_state_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17361),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_1_LC_21_25_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_1_LC_21_25_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_1_LC_21_25_0 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_1_LC_21_25_0  (
            .in0(N__16566),
            .in1(N__17606),
            .in2(N__16834),
            .in3(N__16281),
            .lcout(\this_start_data_delay.this_edge_detector.N_211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_4_LC_21_25_1 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_4_LC_21_25_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_4_LC_21_25_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_4_LC_21_25_1  (
            .in0(N__16282),
            .in1(N__16432),
            .in2(N__16405),
            .in3(N__17625),
            .lcout(\this_start_data_delay.this_edge_detector.N_214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_ns_1_0__m14_LC_21_25_5.C_ON=1'b0;
    defparam M_state_q_ns_1_0__m14_LC_21_25_5.SEQ_MODE=4'b0000;
    defparam M_state_q_ns_1_0__m14_LC_21_25_5.LUT_INIT=16'b0001000001000000;
    LogicCell40 M_state_q_ns_1_0__m14_LC_21_25_5 (
            .in0(N__16283),
            .in1(N__16190),
            .in2(N__16178),
            .in3(N__16165),
            .lcout(),
            .ltout(M_state_q_ns_1_0__i12_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_1_LC_21_25_6.C_ON=1'b0;
    defparam M_state_q_1_LC_21_25_6.SEQ_MODE=4'b1000;
    defparam M_state_q_1_LC_21_25_6.LUT_INIT=16'b0001000101010000;
    LogicCell40 M_state_q_1_LC_21_25_6 (
            .in0(N__17744),
            .in1(N__17607),
            .in2(N__17507),
            .in3(N__17452),
            .lcout(M_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17365),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_0_LC_21_27_0 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_0_LC_21_27_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_0_LC_21_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_this_vram_write_data_0_LC_21_27_0  (
            .in0(_gnd_net_),
            .in1(N__17136),
            .in2(_gnd_net_),
            .in3(N__20285),
            .lcout(M_this_vram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_22_16_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_22_16_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vram.mem_mem_3_0_wclke_3_LC_22_16_2  (
            .in0(N__19318),
            .in1(N__19243),
            .in2(N__19155),
            .in3(N__20327),
            .lcout(\this_vram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI1GH72_12_LC_22_17_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI1GH72_12_LC_22_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI1GH72_12_LC_22_17_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_radreg_RNI1GH72_12_LC_22_17_6  (
            .in0(N__17993),
            .in1(N__19610),
            .in2(_gnd_net_),
            .in3(N__17894),
            .lcout(\this_vram.mem_N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5OL72_12_LC_22_18_0 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5OL72_12_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5OL72_12_LC_22_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_radreg_RNI5OL72_12_LC_22_18_0  (
            .in0(N__19621),
            .in1(N__19412),
            .in2(_gnd_net_),
            .in3(N__18122),
            .lcout(\this_vram.mem_N_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI4K10H_9_LC_22_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI4K10H_9_LC_22_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI4K10H_9_LC_22_18_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI4K10H_9_LC_22_18_5  (
            .in0(N__17924),
            .in1(N__20006),
            .in2(_gnd_net_),
            .in3(N__17777),
            .lcout(N_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_ns_1_0__m7_5_LC_22_24_2.C_ON=1'b0;
    defparam M_state_q_ns_1_0__m7_5_LC_22_24_2.SEQ_MODE=4'b0000;
    defparam M_state_q_ns_1_0__m7_5_LC_22_24_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_state_q_ns_1_0__m7_5_LC_22_24_2 (
            .in0(N__16922),
            .in1(N__16910),
            .in2(N__16893),
            .in3(N__16853),
            .lcout(M_state_q_ns_1_0__m7Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_1_LC_22_25_3 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_1_LC_22_25_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_1_LC_22_25_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_this_vram_write_data_1_LC_22_25_3  (
            .in0(N__16830),
            .in1(N__20284),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_vram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_23_15_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_23_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_23_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_2_0_RNIU0N11_0_LC_23_15_1  (
            .in0(N__19470),
            .in1(N__16703),
            .in2(_gnd_net_),
            .in3(N__18008),
            .lcout(\this_vram.mem_mem_2_0_RNIU0N11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_23_16_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_23_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_23_16_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vram.mem_mem_0_0_wclke_3_LC_23_16_2  (
            .in0(N__19324),
            .in1(N__19239),
            .in2(N__19156),
            .in3(N__20329),
            .lcout(\this_vram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_23_16_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_23_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_23_16_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vram.mem_mem_2_0_wclke_3_LC_23_16_3  (
            .in0(N__20330),
            .in1(N__19149),
            .in2(N__19244),
            .in3(N__19325),
            .lcout(\this_vram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIMTEJ4_11_LC_23_17_0 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIMTEJ4_11_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIMTEJ4_11_LC_23_17_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_radreg_RNIMTEJ4_11_LC_23_17_0  (
            .in0(N__18806),
            .in1(N__17855),
            .in2(_gnd_net_),
            .in3(N__17848),
            .lcout(M_this_vram_read_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_23_17_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_23_17_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_0_0_RNIQOI11_0_LC_23_17_3  (
            .in0(N__17918),
            .in1(N__17909),
            .in2(_gnd_net_),
            .in3(N__19513),
            .lcout(\this_vram.mem_mem_0_0_RNIQOI11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_1_RNI25P11_0_LC_23_17_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_1_RNI25P11_0_LC_23_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_1_RNI25P11_0_LC_23_17_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_3_1_RNI25P11_0_LC_23_17_6  (
            .in0(N__19514),
            .in1(N__17888),
            .in2(_gnd_net_),
            .in3(N__17870),
            .lcout(),
            .ltout(\this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI9OL72_12_LC_23_17_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI9OL72_12_LC_23_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI9OL72_12_LC_23_17_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vram.mem_radreg_RNI9OL72_12_LC_23_17_7  (
            .in0(_gnd_net_),
            .in1(N__18875),
            .in2(N__17858),
            .in3(N__19619),
            .lcout(\this_vram.mem_N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_23_18_1 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_23_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_23_18_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_23_18_1  (
            .in0(N__18914),
            .in1(N__19562),
            .in2(_gnd_net_),
            .in3(N__17849),
            .lcout(M_this_vram_read_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_23_18_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_23_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_23_18_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vram.mem_mem_1_0_wclke_3_LC_23_18_2  (
            .in0(N__19308),
            .in1(N__19237),
            .in2(N__19142),
            .in3(N__20326),
            .lcout(\this_vram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5OL72_0_12_LC_23_18_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5OL72_0_12_LC_23_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5OL72_0_12_LC_23_18_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_radreg_RNI5OL72_0_12_LC_23_18_6  (
            .in0(N__19529),
            .in1(N__18845),
            .in2(_gnd_net_),
            .in3(N__19622),
            .lcout(\this_vram.mem_N_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_23_22_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_23_22_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_23_22_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_23_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI9M0SU_9_LC_23_31_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI9M0SU_9_LC_23_31_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI9M0SU_9_LC_23_31_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI9M0SU_9_LC_23_31_2  (
            .in0(_gnd_net_),
            .in1(N__20021),
            .in2(_gnd_net_),
            .in3(N__18362),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_15_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_15_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_1_1_RNIUSK11_LC_24_15_0  (
            .in0(N__18176),
            .in1(N__18164),
            .in2(_gnd_net_),
            .in3(N__19473),
            .lcout(\this_vram.mem_mem_1_1_RNIUSKZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_15_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_15_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_15_2  (
            .in0(N__18149),
            .in1(N__19472),
            .in2(_gnd_net_),
            .in3(N__18134),
            .lcout(\this_vram.mem_mem_1_0_RNISSK11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_15_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_2_0_RNIU0N11_LC_24_15_3  (
            .in0(N__18110),
            .in1(N__18095),
            .in2(_gnd_net_),
            .in3(N__19474),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_0_RNIU0NZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_15_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_15_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_15_4  (
            .in0(N__18035),
            .in1(_gnd_net_),
            .in2(N__18083),
            .in3(N__19634),
            .lcout(\this_vram.mem_N_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_15_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_0_0_RNIQOI11_LC_24_15_6  (
            .in0(N__18059),
            .in1(N__18050),
            .in2(_gnd_net_),
            .in3(N__19471),
            .lcout(\this_vram.mem_mem_0_0_RNIQOIZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_16_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_16_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_3_1_RNI25P11_LC_24_16_3  (
            .in0(N__18029),
            .in1(N__19516),
            .in2(_gnd_net_),
            .in3(N__18023),
            .lcout(),
            .ltout(\this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_16_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_16_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_16_4  (
            .in0(N__19633),
            .in1(_gnd_net_),
            .in2(N__18923),
            .in3(N__18920),
            .lcout(\this_vram.mem_N_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_16_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_16_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_16_6  (
            .in0(N__18902),
            .in1(N__18890),
            .in2(_gnd_net_),
            .in3(N__19515),
            .lcout(\this_vram.mem_mem_1_1_RNIUSK11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_17_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_17_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_3_0_RNI05P11_LC_24_17_0  (
            .in0(N__18869),
            .in1(N__19519),
            .in2(_gnd_net_),
            .in3(N__18860),
            .lcout(\this_vram.mem_mem_3_0_RNI05PZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_17_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_17_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_17_2  (
            .in0(N__18839),
            .in1(N__18824),
            .in2(_gnd_net_),
            .in3(N__19518),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5GH72_12_LC_24_17_3 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5GH72_12_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5GH72_12_LC_24_17_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vram.mem_radreg_RNI5GH72_12_LC_24_17_3  (
            .in0(N__19620),
            .in1(_gnd_net_),
            .in2(N__18809),
            .in3(N__18776),
            .lcout(\this_vram.mem_N_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_1_RNISOI11_0_LC_24_17_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_1_RNISOI11_0_LC_24_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_1_RNISOI11_0_LC_24_17_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_0_1_RNISOI11_0_LC_24_17_6  (
            .in0(N__18800),
            .in1(N__19517),
            .in2(_gnd_net_),
            .in3(N__18785),
            .lcout(\this_vram.mem_mem_0_1_RNISOI11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_18_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_18_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_2_1_RNI01N11_LC_24_18_2  (
            .in0(N__19522),
            .in1(N__18770),
            .in2(_gnd_net_),
            .in3(N__18755),
            .lcout(\this_vram.mem_mem_2_1_RNI01NZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_18_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_18_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_0_1_RNISOI11_LC_24_18_3  (
            .in0(N__18740),
            .in1(N__19520),
            .in2(_gnd_net_),
            .in3(N__18725),
            .lcout(),
            .ltout(\this_vram.mem_mem_0_1_RNISOIZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_18_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_18_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_18_4  (
            .in0(N__19643),
            .in1(_gnd_net_),
            .in2(N__19637),
            .in3(N__19632),
            .lcout(\this_vram.mem_N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_18_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_18_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_1_0_RNISSK11_LC_24_18_5  (
            .in0(N__19556),
            .in1(N__19521),
            .in2(_gnd_net_),
            .in3(N__19541),
            .lcout(\this_vram.mem_mem_1_0_RNISSKZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_18_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_18_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_18_6  (
            .in0(N__19523),
            .in1(N__19439),
            .in2(_gnd_net_),
            .in3(N__19424),
            .lcout(\this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_24_19_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_24_19_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vram.mem_mem_4_0_wclke_3_LC_24_19_1  (
            .in0(N__19307),
            .in1(N__19238),
            .in2(N__19157),
            .in3(N__20320),
            .lcout(\this_vram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_23_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_23_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vram.mem_mem_5_0_wclke_3_LC_24_23_1  (
            .in0(N__19315),
            .in1(N__19204),
            .in2(N__19151),
            .in3(N__20317),
            .lcout(\this_vram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_24_24_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_24_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_24_24_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vram.mem_mem_6_0_wclke_3_LC_24_24_7  (
            .in0(N__19316),
            .in1(N__19221),
            .in2(N__19150),
            .in3(N__20318),
            .lcout(\this_vram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_25_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_25_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_25_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vram.mem_mem_7_0_wclke_3_LC_24_25_4  (
            .in0(N__19317),
            .in1(N__19222),
            .in2(N__19112),
            .in3(N__20319),
            .lcout(\this_vram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_2_LC_24_26_7 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_2_LC_24_26_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_2_LC_24_26_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_this_vram_write_data_2_LC_24_26_7  (
            .in0(_gnd_net_),
            .in1(N__19035),
            .in2(_gnd_net_),
            .in3(N__20313),
            .lcout(M_this_vram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_3_LC_24_27_5 .C_ON=1'b0;
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_3_LC_24_27_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.this_edge_detector.M_this_vram_write_data_3_LC_24_27_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.this_edge_detector.M_this_vram_write_data_3_LC_24_27_5  (
            .in0(_gnd_net_),
            .in1(N__20349),
            .in2(_gnd_net_),
            .in3(N__20328),
            .lcout(M_this_vram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI3N285N2_9_LC_24_30_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI3N285N2_9_LC_24_30_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI3N285N2_9_LC_24_30_0 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI3N285N2_9_LC_24_30_0  (
            .in0(N__19864),
            .in1(N__20150),
            .in2(N__20020),
            .in3(N__20135),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIGKVAG41_9_LC_26_30_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIGKVAG41_9_LC_26_30_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIGKVAG41_9_LC_26_30_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIGKVAG41_9_LC_26_30_0  (
            .in0(N__20007),
            .in1(N__19865),
            .in2(_gnd_net_),
            .in3(N__19835),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_state_q_ns_1_0__m7_4_LC_32_21_2.C_ON=1'b0;
    defparam M_state_q_ns_1_0__m7_4_LC_32_21_2.SEQ_MODE=4'b0000;
    defparam M_state_q_ns_1_0__m7_4_LC_32_21_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_state_q_ns_1_0__m7_4_LC_32_21_2 (
            .in0(N__19715),
            .in1(N__19694),
            .in2(N__19682),
            .in3(N__19673),
            .lcout(M_state_q_ns_1_0__m7Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
