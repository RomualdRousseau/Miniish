-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 22 2022 16:14:27

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__22940\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \VCCG0\ : std_logic;
signal \this_vga_signals.N_340_0\ : std_logic;
signal \N_198_i\ : std_logic;
signal rgb_c_0 : std_logic;
signal rgb_c_4 : std_logic;
signal port_nmib_0_i : std_logic;
signal rgb_c_3 : std_logic;
signal rgb_c_5 : std_logic;
signal this_vga_signals_vvisibility_i : std_logic;
signal rgb_c_2 : std_logic;
signal rgb_c_1 : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\ : std_logic;
signal \this_vga_ramdac.i2_mux\ : std_logic;
signal \this_vga_ramdac.N_1764_reto\ : std_logic;
signal \this_vga_ramdac.m16\ : std_logic;
signal \this_vga_ramdac.N_1765_reto\ : std_logic;
signal port_clk_c : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal \this_vga_ramdac.N_24_mux\ : std_logic;
signal \this_vga_ramdac.N_1762_reto\ : std_logic;
signal \this_vga_ramdac.m6\ : std_logic;
signal \this_vga_ramdac.N_1763_reto\ : std_logic;
signal \this_vga_ramdac.m19\ : std_logic;
signal \this_vga_ramdac.N_1766_reto\ : std_logic;
signal \this_vga_signals.M_this_vga_signals_pixel_clk_0_0\ : std_logic;
signal \M_pcounter_q_ret_2_RNIRAOL5\ : std_logic;
signal \M_pcounter_q_ret_2_RNIRAOL5_cascade_\ : std_logic;
signal \this_vga_ramdac.i2_mux_0\ : std_logic;
signal \this_vga_ramdac.N_1767_reto\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m7_0_x4_0\ : std_logic;
signal \this_vga_signals.if_N_9_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.if_m1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.N_2_7_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3\ : std_logic;
signal \this_vga_signals.d_N_11\ : std_logic;
signal \this_vga_signals.d_N_12\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc1\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \this_vga_signals.vaddress_1_0_5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.if_i1_mux_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_6_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.if_m1_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3\ : std_logic;
signal \this_vga_signals.if_m1_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_i\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_i_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0\ : std_logic;
signal \this_vga_signals.if_N_2_1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\ : std_logic;
signal \this_vga_signals.g0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1\ : std_logic;
signal \this_vga_signals.N_5_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0\ : std_logic;
signal \this_vga_signals.g1_2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_2_0_0\ : std_logic;
signal \this_vga_signals.g1_3\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNI8OIBAZ0Z_3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.if_N_8_i_0\ : std_logic;
signal \this_vga_signals.g0_9_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_12_x0\ : std_logic;
signal \this_vga_signals.g0_5_0\ : std_logic;
signal \this_vga_signals.N_6_0_cascade_\ : std_logic;
signal \this_vga_signals.N_5\ : std_logic;
signal \this_vga_signals.d_N_3_i_0_0_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_0_cascade_\ : std_logic;
signal \this_vga_signals.N_2_0\ : std_logic;
signal \this_vga_signals.N_2_0_cascade_\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_3_0\ : std_logic;
signal \this_vga_signals.N_3_0\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_3_1\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_1\ : std_logic;
signal \M_this_vga_signals_address_6\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \this_vga_signals.vaddress_1_0_6\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.N_1_4_1_cascade_\ : std_logic;
signal \this_vga_signals.N_7\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_395_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_5_2_cascade_\ : std_logic;
signal \this_vga_signals.g1_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_1_x1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_1\ : std_logic;
signal \this_vga_signals.N_3_1\ : std_logic;
signal \this_vga_signals.vaddress_1_5\ : std_logic;
signal \this_vga_signals.vaddress_1_6_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_1_0_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3\ : std_logic;
signal \this_vga_signals.g0_12_x1\ : std_logic;
signal \this_vga_signals.g0_0_2_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_0\ : std_logic;
signal \this_vga_signals.g0_0_2\ : std_logic;
signal \this_vga_signals.vaddress_6_5\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_1_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_2_0\ : std_logic;
signal \this_vga_signals.N_236\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_3_2\ : std_logic;
signal \this_vga_signals.N_3_2_1\ : std_logic;
signal \this_vga_signals.N_3_2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb2_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2\ : std_logic;
signal \this_vga_signals.SUM_3_i_0_0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_0\ : std_logic;
signal this_vga_signals_hvisibility_i : std_logic;
signal \this_vga_signals.SUM_3_i_0_0_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\ : std_logic;
signal \M_this_vga_ramdac_en_0\ : std_logic;
signal \this_vga_signals.g0_7_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i_0_1_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_2_3\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i_0_0_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_0_3\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_6_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i\ : std_logic;
signal \this_vga_signals.g1_3_0\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.vaddress_4_0_6\ : std_logic;
signal \this_vga_signals.vaddress_5_0_5\ : std_logic;
signal \this_vga_signals.g2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_1\ : std_logic;
signal \this_vga_signals.g1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_1_0_0\ : std_logic;
signal \this_vga_signals.N_5_i_5_cascade_\ : std_logic;
signal \this_vga_signals.N_20_0\ : std_logic;
signal \this_vga_signals.g1_1_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_0_0\ : std_logic;
signal \this_vga_signals.g0_2_x0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.N_5_i_5\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x2_0_2_0\ : std_logic;
signal \this_vga_signals.if_i4_mux_0_0_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_395\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_1_x0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_1\ : std_logic;
signal \this_vga_signals.g0_2_x1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \this_vga_signals.un4_hsynclt8_0_cascade_\ : std_logic;
signal this_vga_signals_hsync_1_i : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.un3_hsynclt8_0\ : std_logic;
signal \this_vga_signals.un6_vvisibilitylto8_0_cascade_\ : std_logic;
signal \this_vga_signals.un6_vvisibilitylt9_0_cascade_\ : std_logic;
signal \this_vga_signals.vvisibility\ : std_logic;
signal \this_vga_signals.g0_7_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_7_repZ0Z1\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_8_repZ0Z1\ : std_logic;
signal \this_vga_signals.vaddress_2_6\ : std_logic;
signal \this_vga_signals.vaddress_2_5\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_2_0_1_0\ : std_logic;
signal \this_vga_signals.g0_22_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_0_0_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0\ : std_logic;
signal \this_vga_signals.vaddress_5_5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_0_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.vaddress_2_0_6\ : std_logic;
signal \this_vga_signals.g2_1\ : std_logic;
signal \this_vga_signals.if_N_5\ : std_logic;
signal \this_vga_signals.vaddress_4_5\ : std_logic;
signal \this_vga_signals.vaddress_3_6\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0\ : std_logic;
signal \this_vga_signals.vaddress_0_5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_0_cascade_\ : std_logic;
signal \this_vga_signals.g2\ : std_logic;
signal \this_vga_signals.g1\ : std_logic;
signal \this_vga_signals.vaddress_0_6\ : std_logic;
signal \this_vga_signals.g1_0_2\ : std_logic;
signal \this_vga_signals.g0_31_1\ : std_logic;
signal \this_vga_signals.g1_0_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_N_2L1\ : std_logic;
signal \this_vga_signals.N_5_1_0_0\ : std_logic;
signal \this_vga_signals.vsync_1_3\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lto7_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.un2_vsynclt8\ : std_logic;
signal \this_vga_signals.N_340_1\ : std_logic;
signal \this_vga_signals.vsync_1_2\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.vaddress_5_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.vaddress_3_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal \this_vga_signals.N_340_0_g\ : std_logic;
signal \this_vga_signals.N_515_g\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z1\ : std_logic;
signal \this_vga_signals.vaddress_5\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z2\ : std_logic;
signal \this_vga_signals.vaddress_4_6\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lto8_1_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal port_enb_c : std_logic;
signal \this_start_data_delay_M_last_q\ : std_logic;
signal \this_vga_signals.vaddress_ac0_9_0_a0_0\ : std_logic;
signal \this_vga_signals.un6_vvisibilitylt9_0\ : std_logic;
signal \this_vga_signals.vaddress_c2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.g1_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt8_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.un4_lvisibility_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.line_clk_1\ : std_logic;
signal \this_vga_signals.un4_lvisibility_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.g0_0\ : std_logic;
signal \N_206_cascade_\ : std_logic;
signal \N_207\ : std_logic;
signal \M_this_state_q_srsts_0_a2_1_4\ : std_logic;
signal port_dmab_c : std_logic;
signal port_dmab_c_i : std_logic;
signal \M_this_ppu_vga_is_drawing_0\ : std_logic;
signal \this_ppu.M_line_clk_out_0_cascade_\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_5\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_4\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_7_cascade_\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_1\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_2\ : std_logic;
signal \M_this_sprites_address_qZ0Z_4\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_4\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_3\ : std_logic;
signal \M_this_sprites_address_qZ0Z_5\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_5\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_4\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_5\ : std_logic;
signal \M_this_sprites_address_qZ0Z_7\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_7\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_6\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_7\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_8\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_9\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_12\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_8\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_8_cascade_\ : std_logic;
signal \M_this_sprites_address_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_11\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_12\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d7_1_0_cascade_\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d7_1_0\ : std_logic;
signal \this_vga_signals.CO0_cascade_\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_1\ : std_logic;
signal \this_ppu.M_line_clk_out_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \M_counter_q_RNIFKS8_1\ : std_logic;
signal \M_counter_q_RNIFKS8_1_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_d7_0\ : std_logic;
signal \M_this_state_q_nss_0\ : std_logic;
signal \this_pixel_clk.M_counter_q_i_1\ : std_logic;
signal \M_this_state_q_srsts_i_1_2\ : std_logic;
signal port_rw_in : std_logic;
signal \N_171_0_cascade_\ : std_logic;
signal \N_176_0\ : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal \N_153_0\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_2\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_9\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_6\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_6\ : std_logic;
signal \M_this_sprites_address_qZ0Z_6\ : std_logic;
signal \M_this_sprites_address_qZ0Z_9\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_9\ : std_logic;
signal \M_this_sprites_address_qZ0Z_1\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c3_cascade_\ : std_logic;
signal \this_ppu.M_haddress_d8lto6_4\ : std_logic;
signal \this_ppu.un1_M_line_clk_out_ns_1_0\ : std_logic;
signal \M_this_vga_signals_line_clk_0\ : std_logic;
signal \this_ppu.line_clk.M_last_qZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_d8\ : std_logic;
signal \this_vga_signals.M_vcounter_q_249_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNIRO2H5Z0Z_9\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_0\ : std_logic;
signal \this_pixel_clk.M_counter_qZ0Z_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_0\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_0\ : std_logic;
signal \M_this_state_q_srsts_i_a2_1_8_1\ : std_logic;
signal \M_this_state_q_srsts_i_a2_1_7_1_cascade_\ : std_logic;
signal \M_this_state_q_srsts_i_a2_1_9_1\ : std_logic;
signal \M_this_state_q_srsts_i_a2_1_6_1\ : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \bfn_17_23_0_\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \un1_M_this_data_count_q_cry_0\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \un1_M_this_data_count_q_cry_1\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \un1_M_this_data_count_q_cry_2\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \un1_M_this_data_count_q_cry_3\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \un1_M_this_data_count_q_cry_4\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \un1_M_this_data_count_q_cry_5\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \un1_M_this_data_count_q_cry_6\ : std_logic;
signal \un1_M_this_data_count_q_cry_7\ : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \bfn_17_24_0_\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \un1_M_this_data_count_q_cry_8\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \un1_M_this_data_count_q_cry_9\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \un1_M_this_data_count_q_cry_10\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \un1_M_this_data_count_q_cry_11\ : std_logic;
signal \M_this_state_q_RNI20CEZ0Z_0\ : std_logic;
signal \un1_M_this_data_count_q_cry_12\ : std_logic;
signal \un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO\ : std_logic;
signal \un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO\ : std_logic;
signal \bfn_17_25_0_\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c5_cascade_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c5\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c2\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c1\ : std_logic;
signal port_address_in_0 : std_logic;
signal port_address_in_1 : std_logic;
signal \N_218\ : std_logic;
signal \N_204\ : std_logic;
signal \N_202\ : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal \N_233\ : std_logic;
signal \M_this_start_address_delay_out_0\ : std_logic;
signal \M_this_state_q_srsts_i_1_1_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal \this_ppu.N_250_1\ : std_logic;
signal \this_ppu.M_last_q_RNI5NOQ4\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c3\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c5\ : std_logic;
signal \this_ppu.N_258_1\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c5_cascade_\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_13\ : std_logic;
signal \M_this_sprites_address_qZ0Z_2\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_2\ : std_logic;
signal \M_this_ppu_vram_data_3\ : std_logic;
signal \M_this_ppu_sprites_addr_1\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_10\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_10\ : std_logic;
signal \M_this_sprites_address_qZ0Z_10\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal \M_this_sprites_address_q_3_sm0_0\ : std_logic;
signal \M_this_sprites_address_q_3_ns_1_3_cascade_\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_3\ : std_logic;
signal \M_this_sprites_address_qZ0Z_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_3\ : std_logic;
signal \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_3\ : std_logic;
signal \this_sprites_ram_mem_N_102\ : std_logic;
signal \M_this_ppu_vram_data_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_1\ : std_logic;
signal \this_sprites_ram_mem_N_91\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_1\ : std_logic;
signal \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_1\ : std_logic;
signal \M_this_ppu_vram_addr_1\ : std_logic;
signal \bfn_21_17_0_\ : std_logic;
signal \M_this_ppu_vram_addr_2\ : std_logic;
signal \M_this_ppu_sprites_addr_2\ : std_logic;
signal \this_ppu.sprites_addr_cry_1\ : std_logic;
signal \M_this_ppu_vram_addr_3\ : std_logic;
signal \M_this_ppu_sprites_addr_3\ : std_logic;
signal \this_ppu.sprites_addr_cry_2\ : std_logic;
signal \M_this_ppu_vram_addr_4\ : std_logic;
signal \M_this_ppu_sprites_addr_4\ : std_logic;
signal \this_ppu.sprites_addr_cry_3\ : std_logic;
signal \M_this_ppu_vram_addr_5\ : std_logic;
signal \M_this_ppu_sprites_addr_5\ : std_logic;
signal \this_ppu.sprites_addr_cry_4\ : std_logic;
signal \M_this_ppu_vram_addr_6\ : std_logic;
signal \M_this_ppu_sprites_addr_6\ : std_logic;
signal \this_ppu.sprites_addr_cry_5\ : std_logic;
signal \M_this_ppu_vram_addr_7\ : std_logic;
signal \M_this_ppu_sprites_addr_7\ : std_logic;
signal \this_ppu.sprites_addr_cry_6\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_1\ : std_logic;
signal \M_this_ppu_sprites_addr_8\ : std_logic;
signal \this_ppu.sprites_addr_cry_7\ : std_logic;
signal \this_ppu.sprites_addr_cry_8\ : std_logic;
signal \this_ppu.M_vaddress_qZ1Z_2\ : std_logic;
signal \M_this_ppu_sprites_addr_9\ : std_logic;
signal \bfn_21_18_0_\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_3\ : std_logic;
signal \M_this_ppu_sprites_addr_10\ : std_logic;
signal \this_ppu.sprites_addr_cry_9\ : std_logic;
signal \this_ppu.M_vaddress_qZ1Z_4\ : std_logic;
signal \this_ppu.sprites_addr_cry_10\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_5\ : std_logic;
signal \this_ppu.sprites_addr_cry_11\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_6\ : std_logic;
signal \this_ppu.sprites_addr_cry_12\ : std_logic;
signal \M_this_ppu_vram_addr_0\ : std_logic;
signal \M_this_ppu_vram_addr_i_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_1\ : std_logic;
signal \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_1_cascade_\ : std_logic;
signal \this_sprites_ram_mem_N_88\ : std_logic;
signal \this_sprites_ram.mem_WE_14\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_3\ : std_logic;
signal \this_sprites_ram_mem_N_105\ : std_logic;
signal \N_200\ : std_logic;
signal \M_this_ppu_vram_data_2\ : std_logic;
signal \M_this_ppu_vram_en_0\ : std_logic;
signal this_sprites_ram_mem_radreg_11 : std_logic;
signal \M_this_ppu_vram_data_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_3\ : std_logic;
signal \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_3\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal \N_170_0\ : std_logic;
signal \this_sprites_ram.mem_WE_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_2\ : std_logic;
signal \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_2_cascade_\ : std_logic;
signal \this_sprites_ram_mem_N_98\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_0_cascade_\ : std_logic;
signal \this_sprites_ram_mem_N_109\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_0\ : std_logic;
signal \this_sprites_ram_mem_N_112\ : std_logic;
signal \this_sprites_ram.mem_WE_10\ : std_logic;
signal \this_sprites_ram.mem_WE_8\ : std_logic;
signal \this_sprites_ram.mem_WE_12\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_2\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_13\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_2\ : std_logic;
signal \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_2_cascade_\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_12\ : std_logic;
signal \this_sprites_ram_mem_N_95\ : std_logic;
signal \this_sprites_ram.mem_WE_6\ : std_logic;
signal \this_sprites_ram.mem_WE_4\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal \M_this_start_data_delay_out_0\ : std_logic;
signal port_data_c_0 : std_logic;
signal port_data_c_4 : std_logic;
signal \M_this_sprites_ram_write_data_0_sqmuxa_cascade_\ : std_logic;
signal \M_this_sprites_ram_write_data_0_i_0\ : std_logic;
signal port_data_c_3 : std_logic;
signal port_data_c_7 : std_logic;
signal \M_this_sprites_ram_write_data_0_i_3\ : std_logic;
signal port_data_c_2 : std_logic;
signal port_data_c_6 : std_logic;
signal \M_this_sprites_ram_write_data_0_i_2\ : std_logic;
signal port_data_c_1 : std_logic;
signal \un1_M_this_state_q_2_0\ : std_logic;
signal port_data_c_5 : std_logic;
signal \M_this_sprites_ram_write_data_0_sqmuxa\ : std_logic;
signal \M_this_sprites_ram_write_data_0_i_1\ : std_logic;
signal \M_this_sprites_address_qZ0Z_12\ : std_logic;
signal \M_this_sprites_ram_write_en_1_0_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_13\ : std_logic;
signal \M_this_sprites_address_qZ0Z_11\ : std_logic;
signal \this_sprites_ram.mem_WE_2\ : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal \M_this_external_address_qZ0Z_0\ : std_logic;
signal \bfn_30_23_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_external_address_q_cry_0\ : std_logic;
signal \M_this_external_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_external_address_q_cry_1\ : std_logic;
signal \M_this_external_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_external_address_q_cry_2\ : std_logic;
signal \M_this_external_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_external_address_q_cry_3\ : std_logic;
signal \M_this_external_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_external_address_q_cry_4\ : std_logic;
signal \M_this_external_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_5\ : std_logic;
signal \M_this_external_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_external_address_q_cry_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_7\ : std_logic;
signal \M_this_external_address_qZ0Z_8\ : std_logic;
signal \bfn_30_24_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_external_address_q_cry_8\ : std_logic;
signal \M_this_external_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_external_address_q_cry_9\ : std_logic;
signal \M_this_external_address_qZ0Z_11\ : std_logic;
signal \un1_M_this_external_address_q_cry_10\ : std_logic;
signal \M_this_external_address_qZ0Z_12\ : std_logic;
signal \un1_M_this_external_address_q_cry_11\ : std_logic;
signal \M_this_external_address_qZ0Z_13\ : std_logic;
signal \un1_M_this_external_address_q_cry_12\ : std_logic;
signal \M_this_external_address_qZ0Z_14\ : std_logic;
signal \un1_M_this_external_address_q_cry_13\ : std_logic;
signal \M_this_state_qZ0Z_0\ : std_logic;
signal \un1_M_this_external_address_q_cry_14\ : std_logic;
signal \M_this_external_address_qZ0Z_15\ : std_logic;
signal clk_0_c_g : std_logic;
signal \M_this_state_q_nss_g_0\ : std_logic;
signal port_address_in_3 : std_logic;
signal port_address_in_4 : std_logic;
signal port_address_in_5 : std_logic;
signal port_address_in_2 : std_logic;
signal port_address_in_7 : std_logic;
signal \M_this_state_d36_2_0_3_cascade_\ : std_logic;
signal port_address_in_6 : std_logic;
signal \M_this_state_d37_1\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \this_sprites_ram.mem_out_bus0_1\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_0\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ <= \N__19100\&\N__17630\&\N__17771\&\N__17918\&\N__18083\&\N__18242\&\N__18395\&\N__18557\&\N__16985\&\N__16664\&\N__18848\;
    \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ <= \N__16541\&\N__14810\&\N__14030\&\N__13604\&\N__14927\&\N__13742\&\N__13868\&\N__17417\&\N__16817\&\N__14672\&\N__15374\;
    \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21410\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20072\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus0_3\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_2\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ <= \N__19094\&\N__17624\&\N__17765\&\N__17912\&\N__18077\&\N__18236\&\N__18389\&\N__18551\&\N__16979\&\N__16658\&\N__18842\;
    \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ <= \N__16535\&\N__14804\&\N__14024\&\N__13598\&\N__14921\&\N__13736\&\N__13862\&\N__17411\&\N__16811\&\N__14666\&\N__15368\;
    \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19922\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19748\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_1\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_0\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ <= \N__19088\&\N__17618\&\N__17759\&\N__17906\&\N__18071\&\N__18230\&\N__18383\&\N__18545\&\N__16973\&\N__16652\&\N__18836\;
    \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ <= \N__16529\&\N__14798\&\N__14018\&\N__13592\&\N__14915\&\N__13730\&\N__13856\&\N__17405\&\N__16805\&\N__14660\&\N__15362\;
    \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21406\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20068\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_3\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_2\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ <= \N__19082\&\N__17612\&\N__17753\&\N__17900\&\N__18065\&\N__18224\&\N__18377\&\N__18539\&\N__16967\&\N__16646\&\N__18830\;
    \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ <= \N__16523\&\N__14792\&\N__14012\&\N__13586\&\N__14909\&\N__13724\&\N__13850\&\N__17399\&\N__16799\&\N__14654\&\N__15356\;
    \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19918\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19744\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_1\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_0\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ <= \N__19076\&\N__17606\&\N__17747\&\N__17894\&\N__18059\&\N__18218\&\N__18371\&\N__18533\&\N__16961\&\N__16640\&\N__18824\;
    \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ <= \N__16517\&\N__14786\&\N__14006\&\N__13580\&\N__14903\&\N__13718\&\N__13844\&\N__17393\&\N__16793\&\N__14648\&\N__15350\;
    \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21399\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20061\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_3\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_2\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ <= \N__19070\&\N__17600\&\N__17741\&\N__17888\&\N__18053\&\N__18212\&\N__18365\&\N__18527\&\N__16955\&\N__16634\&\N__18818\;
    \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ <= \N__16511\&\N__14780\&\N__14000\&\N__13574\&\N__14897\&\N__13712\&\N__13838\&\N__17387\&\N__16787\&\N__14642\&\N__15344\;
    \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19911\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19736\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_1\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_0\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ <= \N__19064\&\N__17594\&\N__17735\&\N__17882\&\N__18047\&\N__18206\&\N__18359\&\N__18521\&\N__16949\&\N__16628\&\N__18812\;
    \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ <= \N__16505\&\N__14774\&\N__13994\&\N__13568\&\N__14891\&\N__13706\&\N__13832\&\N__17381\&\N__16781\&\N__14636\&\N__15338\;
    \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21390\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20051\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_3\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_2\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ <= \N__19058\&\N__17588\&\N__17729\&\N__17876\&\N__18041\&\N__18200\&\N__18353\&\N__18515\&\N__16943\&\N__16622\&\N__18806\;
    \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ <= \N__16499\&\N__14768\&\N__13988\&\N__13562\&\N__14885\&\N__13700\&\N__13826\&\N__17375\&\N__16775\&\N__14630\&\N__15332\;
    \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19902\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19723\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_1\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_0\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ <= \N__19052\&\N__17582\&\N__17723\&\N__17870\&\N__18035\&\N__18194\&\N__18347\&\N__18509\&\N__16937\&\N__16616\&\N__18800\;
    \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ <= \N__16493\&\N__14762\&\N__13982\&\N__13556\&\N__14879\&\N__13694\&\N__13820\&\N__17369\&\N__16769\&\N__14624\&\N__15326\;
    \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21380\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20038\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_3\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_2\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ <= \N__19046\&\N__17576\&\N__17717\&\N__17864\&\N__18029\&\N__18188\&\N__18341\&\N__18503\&\N__16931\&\N__16610\&\N__18794\;
    \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ <= \N__16487\&\N__14756\&\N__13976\&\N__13550\&\N__14873\&\N__13688\&\N__13814\&\N__17363\&\N__16763\&\N__14618\&\N__15320\;
    \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19888\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19708\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_1\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_0\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ <= \N__19040\&\N__17570\&\N__17711\&\N__17858\&\N__18023\&\N__18182\&\N__18335\&\N__18497\&\N__16925\&\N__16604\&\N__18788\;
    \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ <= \N__16481\&\N__14750\&\N__13970\&\N__13544\&\N__14867\&\N__13682\&\N__13808\&\N__17357\&\N__16757\&\N__14612\&\N__15314\;
    \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21367\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20003\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_3\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_2\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ <= \N__19034\&\N__17564\&\N__17705\&\N__17852\&\N__18017\&\N__18176\&\N__18329\&\N__18491\&\N__16919\&\N__16598\&\N__18782\;
    \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ <= \N__16475\&\N__14744\&\N__13964\&\N__13538\&\N__14861\&\N__13676\&\N__13802\&\N__17351\&\N__16751\&\N__14606\&\N__15308\;
    \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19862\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19694\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_1\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_0\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ <= \N__19028\&\N__17558\&\N__17699\&\N__17846\&\N__18011\&\N__18170\&\N__18323\&\N__18485\&\N__16913\&\N__16592\&\N__18776\;
    \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ <= \N__16469\&\N__14738\&\N__13958\&\N__13532\&\N__14855\&\N__13670\&\N__13796\&\N__17345\&\N__16745\&\N__14600\&\N__15302\;
    \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21376\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20034\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_3\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_2\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ <= \N__19022\&\N__17552\&\N__17693\&\N__17840\&\N__18005\&\N__18164\&\N__18317\&\N__18479\&\N__16907\&\N__16586\&\N__18770\;
    \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ <= \N__16463\&\N__14732\&\N__13952\&\N__13526\&\N__14849\&\N__13664\&\N__13790\&\N__17339\&\N__16739\&\N__14594\&\N__15296\;
    \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19889\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19732\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_1\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_0\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ <= \N__19016\&\N__17546\&\N__17687\&\N__17834\&\N__17999\&\N__18158\&\N__18311\&\N__18473\&\N__16901\&\N__16580\&\N__18764\;
    \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ <= \N__16457\&\N__14726\&\N__13946\&\N__13520\&\N__14843\&\N__13658\&\N__13784\&\N__17333\&\N__16733\&\N__14588\&\N__15290\;
    \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21389\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20050\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_3\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_2\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ <= \N__19010\&\N__17540\&\N__17681\&\N__17828\&\N__17993\&\N__18152\&\N__18305\&\N__18467\&\N__16895\&\N__16574\&\N__18758\;
    \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ <= \N__16451\&\N__14720\&\N__13940\&\N__13514\&\N__14837\&\N__13652\&\N__13778\&\N__17327\&\N__16727\&\N__14582\&\N__15284\;
    \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19901\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19743\&'0'&'0'&'0';
    \M_this_vram_read_data_3\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_vram_read_data_2\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_vram_read_data_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_vram_read_data_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__8381\&\N__8672\&\N__8243\&\N__8231\&\N__8630\&\N__8048\&\N__8036\&\N__8339\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__17966\&\N__18128\&\N__18281\&\N__18443\&\N__18602\&\N__17045\&\N__17114\&\N__18920\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__16676\&\N__19409\&\N__17210\&\N__19229\;

    \this_sprites_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22166\,
            RE => \N__15906\,
            WCLKE => \N__18677\,
            WCLK => \N__22167\,
            WE => \N__15908\
        );

    \this_sprites_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22168\,
            RE => \N__15905\,
            WCLKE => \N__18670\,
            WCLK => \N__22169\,
            WE => \N__15907\
        );

    \this_sprites_ram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22170\,
            RE => \N__15889\,
            WCLKE => \N__19445\,
            WCLK => \N__22171\,
            WE => \N__15903\
        );

    \this_sprites_ram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22172\,
            RE => \N__15888\,
            WCLKE => \N__19441\,
            WCLK => \N__22173\,
            WE => \N__15902\
        );

    \this_sprites_ram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22179\,
            RE => \N__15854\,
            WCLKE => \N__19487\,
            WCLK => \N__22178\,
            WE => \N__15876\
        );

    \this_sprites_ram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22186\,
            RE => \N__15853\,
            WCLKE => \N__19486\,
            WCLK => \N__22187\,
            WE => \N__15875\
        );

    \this_sprites_ram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22199\,
            RE => \N__15799\,
            WCLKE => \N__19459\,
            WCLK => \N__22200\,
            WE => \N__15848\
        );

    \this_sprites_ram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22209\,
            RE => \N__15798\,
            WCLKE => \N__19463\,
            WCLK => \N__22210\,
            WE => \N__15790\
        );

    \this_sprites_ram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22219\,
            RE => \N__15734\,
            WCLKE => \N__20431\,
            WCLK => \N__22220\,
            WE => \N__15786\
        );

    \this_sprites_ram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22225\,
            RE => \N__15733\,
            WCLKE => \N__20435\,
            WCLK => \N__22226\,
            WE => \N__15688\
        );

    \this_sprites_ram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22227\,
            RE => \N__15758\,
            WCLKE => \N__20413\,
            WCLK => \N__22228\,
            WE => \N__15774\
        );

    \this_sprites_ram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22233\,
            RE => \N__15759\,
            WCLKE => \N__20414\,
            WCLK => \N__22234\,
            WE => \N__15840\
        );

    \this_sprites_ram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22235\,
            RE => \N__15829\,
            WCLKE => \N__20989\,
            WCLK => \N__22236\,
            WE => \N__15841\
        );

    \this_sprites_ram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22237\,
            RE => \N__15830\,
            WCLKE => \N__20993\,
            WCLK => \N__22238\,
            WE => \N__15880\
        );

    \this_sprites_ram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22240\,
            RE => \N__15881\,
            WCLKE => \N__19147\,
            WCLK => \N__22241\,
            WE => \N__15883\
        );

    \this_sprites_ram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22243\,
            RE => \N__15882\,
            WCLKE => \N__19151\,
            WCLK => \N__22244\,
            WE => \N__15904\
        );

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22175\,
            RE => \N__15887\,
            WCLKE => \N__19386\,
            WCLK => \N__22174\,
            WE => \N__15849\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__22938\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22940\,
            DIN => \N__22939\,
            DOUT => \N__22938\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22940\,
            PADOUT => \N__22939\,
            PADIN => \N__22938\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22929\,
            DIN => \N__22928\,
            DOUT => \N__22927\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22929\,
            PADOUT => \N__22928\,
            PADIN => \N__22927\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22920\,
            DIN => \N__22919\,
            DOUT => \N__22918\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22920\,
            PADOUT => \N__22919\,
            PADIN => \N__22918\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22911\,
            DIN => \N__22910\,
            DOUT => \N__22909\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22911\,
            PADOUT => \N__22910\,
            PADIN => \N__22909\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__9443\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22902\,
            DIN => \N__22901\,
            DOUT => \N__22900\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22902\,
            PADOUT => \N__22901\,
            PADIN => \N__22900\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10163\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22893\,
            DIN => \N__22892\,
            DOUT => \N__22891\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22893\,
            PADOUT => \N__22892\,
            PADIN => \N__22891\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__20837\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13042\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22884\,
            DIN => \N__22883\,
            DOUT => \N__22882\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22884\,
            PADOUT => \N__22883\,
            PADIN => \N__22882\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__20813\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13052\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22875\,
            DIN => \N__22874\,
            DOUT => \N__22873\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22875\,
            PADOUT => \N__22874\,
            PADIN => \N__22873\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__20789\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13099\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22866\,
            DIN => \N__22865\,
            DOUT => \N__22864\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22866\,
            PADOUT => \N__22865\,
            PADIN => \N__22864\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__20759\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13120\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22857\,
            DIN => \N__22856\,
            DOUT => \N__22855\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22857\,
            PADOUT => \N__22856\,
            PADIN => \N__22855\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__20735\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13035\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22848\,
            DIN => \N__22847\,
            DOUT => \N__22846\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22848\,
            PADOUT => \N__22847\,
            PADIN => \N__22846\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__20717\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13109\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22839\,
            DIN => \N__22838\,
            DOUT => \N__22837\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22839\,
            PADOUT => \N__22838\,
            PADIN => \N__22837\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__21734\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13124\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22830\,
            DIN => \N__22829\,
            DOUT => \N__22828\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22830\,
            PADOUT => \N__22829\,
            PADIN => \N__22828\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__21713\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13142\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22821\,
            DIN => \N__22820\,
            DOUT => \N__22819\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22821\,
            PADOUT => \N__22820\,
            PADIN => \N__22819\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21632\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13068\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22812\,
            DIN => \N__22811\,
            DOUT => \N__22810\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22812\,
            PADOUT => \N__22811\,
            PADIN => \N__22810\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21602\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13129\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22803\,
            DIN => \N__22802\,
            DOUT => \N__22801\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22803\,
            PADOUT => \N__22802\,
            PADIN => \N__22801\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21584\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13102\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22794\,
            DIN => \N__22793\,
            DOUT => \N__22792\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22794\,
            PADOUT => \N__22793\,
            PADIN => \N__22792\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21566\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13110\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22785\,
            DIN => \N__22784\,
            DOUT => \N__22783\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22785\,
            PADOUT => \N__22784\,
            PADIN => \N__22783\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__22532\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13125\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22776\,
            DIN => \N__22775\,
            DOUT => \N__22774\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22776\,
            PADOUT => \N__22775\,
            PADIN => \N__22774\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__22268\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13141\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22767\,
            DIN => \N__22766\,
            DOUT => \N__22765\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22767\,
            PADOUT => \N__22766\,
            PADIN => \N__22765\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21686\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13041\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22758\,
            DIN => \N__22757\,
            DOUT => \N__22756\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22758\,
            PADOUT => \N__22757\,
            PADIN => \N__22756\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21653\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13100\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22749\,
            DIN => \N__22748\,
            DOUT => \N__22747\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22749\,
            PADOUT => \N__22748\,
            PADIN => \N__22747\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22740\,
            DIN => \N__22739\,
            DOUT => \N__22738\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22740\,
            PADOUT => \N__22739\,
            PADIN => \N__22738\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22731\,
            DIN => \N__22730\,
            DOUT => \N__22729\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22731\,
            PADOUT => \N__22730\,
            PADIN => \N__22729\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22722\,
            DIN => \N__22721\,
            DOUT => \N__22720\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22722\,
            PADOUT => \N__22721\,
            PADIN => \N__22720\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22713\,
            DIN => \N__22712\,
            DOUT => \N__22711\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22713\,
            PADOUT => \N__22712\,
            PADIN => \N__22711\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22704\,
            DIN => \N__22703\,
            DOUT => \N__22702\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22704\,
            PADOUT => \N__22703\,
            PADIN => \N__22702\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22695\,
            DIN => \N__22694\,
            DOUT => \N__22693\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22695\,
            PADOUT => \N__22694\,
            PADIN => \N__22693\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22686\,
            DIN => \N__22685\,
            DOUT => \N__22684\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22686\,
            PADOUT => \N__22685\,
            PADIN => \N__22684\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22677\,
            DIN => \N__22676\,
            DOUT => \N__22675\,
            PACKAGEPIN => port_data_wire(7)
        );

    \port_data_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22677\,
            PADOUT => \N__22676\,
            PADIN => \N__22675\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22668\,
            DIN => \N__22667\,
            DOUT => \N__22666\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22668\,
            PADOUT => \N__22667\,
            PADIN => \N__22666\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7643\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22659\,
            DIN => \N__22658\,
            DOUT => \N__22657\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22659\,
            PADOUT => \N__22658\,
            PADIN => \N__22657\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13217\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22650\,
            DIN => \N__22649\,
            DOUT => \N__22648\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22650\,
            PADOUT => \N__22649\,
            PADIN => \N__22648\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22641\,
            DIN => \N__22640\,
            DOUT => \N__22639\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22641\,
            PADOUT => \N__22640\,
            PADIN => \N__22639\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7601\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22632\,
            DIN => \N__22631\,
            DOUT => \N__22630\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__22632\,
            PADOUT => \N__22631\,
            PADIN => \N__22630\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__15797\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13101\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22623\,
            DIN => \N__22622\,
            DOUT => \N__22621\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22623\,
            PADOUT => \N__22622\,
            PADIN => \N__22621\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7637\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22614\,
            DIN => \N__22613\,
            DOUT => \N__22612\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22614\,
            PADOUT => \N__22613\,
            PADIN => \N__22612\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7814\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22605\,
            DIN => \N__22604\,
            DOUT => \N__22603\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22605\,
            PADOUT => \N__22604\,
            PADIN => \N__22603\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7829\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22596\,
            DIN => \N__22595\,
            DOUT => \N__22594\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22596\,
            PADOUT => \N__22595\,
            PADIN => \N__22594\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7589\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22587\,
            DIN => \N__22586\,
            DOUT => \N__22585\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22587\,
            PADOUT => \N__22586\,
            PADIN => \N__22585\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7619\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22578\,
            DIN => \N__22577\,
            DOUT => \N__22576\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22578\,
            PADOUT => \N__22577\,
            PADIN => \N__22576\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7577\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22569\,
            DIN => \N__22568\,
            DOUT => \N__22567\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22569\,
            PADOUT => \N__22568\,
            PADIN => \N__22567\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22560\,
            DIN => \N__22559\,
            DOUT => \N__22558\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22560\,
            PADOUT => \N__22559\,
            PADIN => \N__22558\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7841\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22551\,
            DIN => \N__22550\,
            DOUT => \N__22549\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22551\,
            PADOUT => \N__22550\,
            PADIN => \N__22549\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11210\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__5534\ : IoInMux
    port map (
            O => \N__22532\,
            I => \N__22529\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__22529\,
            I => \N__22526\
        );

    \I__5532\ : Span4Mux_s2_h
    port map (
            O => \N__22526\,
            I => \N__22523\
        );

    \I__5531\ : Sp12to4
    port map (
            O => \N__22523\,
            I => \N__22519\
        );

    \I__5530\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22516\
        );

    \I__5529\ : Odrv12
    port map (
            O => \N__22519\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__22516\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__5527\ : InMux
    port map (
            O => \N__22511\,
            I => \un1_M_this_external_address_q_cry_13\
        );

    \I__5526\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22493\
        );

    \I__5525\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22493\
        );

    \I__5524\ : InMux
    port map (
            O => \N__22506\,
            I => \N__22493\
        );

    \I__5523\ : InMux
    port map (
            O => \N__22505\,
            I => \N__22493\
        );

    \I__5522\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22493\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__22493\,
            I => \N__22479\
        );

    \I__5520\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22472\
        );

    \I__5519\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22472\
        );

    \I__5518\ : InMux
    port map (
            O => \N__22490\,
            I => \N__22472\
        );

    \I__5517\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22463\
        );

    \I__5516\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22463\
        );

    \I__5515\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22463\
        );

    \I__5514\ : InMux
    port map (
            O => \N__22486\,
            I => \N__22463\
        );

    \I__5513\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22454\
        );

    \I__5512\ : InMux
    port map (
            O => \N__22484\,
            I => \N__22454\
        );

    \I__5511\ : InMux
    port map (
            O => \N__22483\,
            I => \N__22454\
        );

    \I__5510\ : InMux
    port map (
            O => \N__22482\,
            I => \N__22454\
        );

    \I__5509\ : Span4Mux_v
    port map (
            O => \N__22479\,
            I => \N__22444\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__22472\,
            I => \N__22439\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__22463\,
            I => \N__22439\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__22454\,
            I => \N__22436\
        );

    \I__5505\ : CascadeMux
    port map (
            O => \N__22453\,
            I => \N__22432\
        );

    \I__5504\ : CascadeMux
    port map (
            O => \N__22452\,
            I => \N__22429\
        );

    \I__5503\ : CascadeMux
    port map (
            O => \N__22451\,
            I => \N__22424\
        );

    \I__5502\ : CascadeMux
    port map (
            O => \N__22450\,
            I => \N__22416\
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__22449\,
            I => \N__22413\
        );

    \I__5500\ : CascadeMux
    port map (
            O => \N__22448\,
            I => \N__22410\
        );

    \I__5499\ : CascadeMux
    port map (
            O => \N__22447\,
            I => \N__22407\
        );

    \I__5498\ : Span4Mux_s1_h
    port map (
            O => \N__22444\,
            I => \N__22400\
        );

    \I__5497\ : Span4Mux_v
    port map (
            O => \N__22439\,
            I => \N__22400\
        );

    \I__5496\ : Span4Mux_v
    port map (
            O => \N__22436\,
            I => \N__22400\
        );

    \I__5495\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22397\
        );

    \I__5494\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22392\
        );

    \I__5493\ : InMux
    port map (
            O => \N__22429\,
            I => \N__22385\
        );

    \I__5492\ : InMux
    port map (
            O => \N__22428\,
            I => \N__22385\
        );

    \I__5491\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22385\
        );

    \I__5490\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22382\
        );

    \I__5489\ : InMux
    port map (
            O => \N__22423\,
            I => \N__22379\
        );

    \I__5488\ : InMux
    port map (
            O => \N__22422\,
            I => \N__22376\
        );

    \I__5487\ : CascadeMux
    port map (
            O => \N__22421\,
            I => \N__22372\
        );

    \I__5486\ : CascadeMux
    port map (
            O => \N__22420\,
            I => \N__22369\
        );

    \I__5485\ : CascadeMux
    port map (
            O => \N__22419\,
            I => \N__22366\
        );

    \I__5484\ : InMux
    port map (
            O => \N__22416\,
            I => \N__22362\
        );

    \I__5483\ : InMux
    port map (
            O => \N__22413\,
            I => \N__22357\
        );

    \I__5482\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22357\
        );

    \I__5481\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22354\
        );

    \I__5480\ : Span4Mux_h
    port map (
            O => \N__22400\,
            I => \N__22351\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__22397\,
            I => \N__22348\
        );

    \I__5478\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22343\
        );

    \I__5477\ : InMux
    port map (
            O => \N__22395\,
            I => \N__22343\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__22392\,
            I => \N__22338\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__22385\,
            I => \N__22338\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22333\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__22379\,
            I => \N__22333\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__22376\,
            I => \N__22330\
        );

    \I__5471\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22327\
        );

    \I__5470\ : InMux
    port map (
            O => \N__22372\,
            I => \N__22324\
        );

    \I__5469\ : InMux
    port map (
            O => \N__22369\,
            I => \N__22321\
        );

    \I__5468\ : InMux
    port map (
            O => \N__22366\,
            I => \N__22316\
        );

    \I__5467\ : InMux
    port map (
            O => \N__22365\,
            I => \N__22316\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__22362\,
            I => \N__22309\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__22357\,
            I => \N__22309\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__22354\,
            I => \N__22309\
        );

    \I__5463\ : Span4Mux_h
    port map (
            O => \N__22351\,
            I => \N__22306\
        );

    \I__5462\ : Span4Mux_h
    port map (
            O => \N__22348\,
            I => \N__22301\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__22343\,
            I => \N__22301\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__22338\,
            I => \N__22296\
        );

    \I__5459\ : Span4Mux_v
    port map (
            O => \N__22333\,
            I => \N__22296\
        );

    \I__5458\ : Span4Mux_h
    port map (
            O => \N__22330\,
            I => \N__22291\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__22327\,
            I => \N__22291\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__22324\,
            I => \N__22278\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__22321\,
            I => \N__22278\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__22316\,
            I => \N__22278\
        );

    \I__5453\ : Span4Mux_v
    port map (
            O => \N__22309\,
            I => \N__22278\
        );

    \I__5452\ : Span4Mux_h
    port map (
            O => \N__22306\,
            I => \N__22278\
        );

    \I__5451\ : Span4Mux_v
    port map (
            O => \N__22301\,
            I => \N__22278\
        );

    \I__5450\ : Odrv4
    port map (
            O => \N__22296\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__22291\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__22278\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__5447\ : InMux
    port map (
            O => \N__22271\,
            I => \un1_M_this_external_address_q_cry_14\
        );

    \I__5446\ : IoInMux
    port map (
            O => \N__22268\,
            I => \N__22265\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__22265\,
            I => \N__22262\
        );

    \I__5444\ : Span4Mux_s2_h
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__5443\ : Sp12to4
    port map (
            O => \N__22259\,
            I => \N__22256\
        );

    \I__5442\ : Span12Mux_v
    port map (
            O => \N__22256\,
            I => \N__22252\
        );

    \I__5441\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22249\
        );

    \I__5440\ : Odrv12
    port map (
            O => \N__22252\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__22249\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__5438\ : ClkMux
    port map (
            O => \N__22244\,
            I => \N__22007\
        );

    \I__5437\ : ClkMux
    port map (
            O => \N__22243\,
            I => \N__22007\
        );

    \I__5436\ : ClkMux
    port map (
            O => \N__22242\,
            I => \N__22007\
        );

    \I__5435\ : ClkMux
    port map (
            O => \N__22241\,
            I => \N__22007\
        );

    \I__5434\ : ClkMux
    port map (
            O => \N__22240\,
            I => \N__22007\
        );

    \I__5433\ : ClkMux
    port map (
            O => \N__22239\,
            I => \N__22007\
        );

    \I__5432\ : ClkMux
    port map (
            O => \N__22238\,
            I => \N__22007\
        );

    \I__5431\ : ClkMux
    port map (
            O => \N__22237\,
            I => \N__22007\
        );

    \I__5430\ : ClkMux
    port map (
            O => \N__22236\,
            I => \N__22007\
        );

    \I__5429\ : ClkMux
    port map (
            O => \N__22235\,
            I => \N__22007\
        );

    \I__5428\ : ClkMux
    port map (
            O => \N__22234\,
            I => \N__22007\
        );

    \I__5427\ : ClkMux
    port map (
            O => \N__22233\,
            I => \N__22007\
        );

    \I__5426\ : ClkMux
    port map (
            O => \N__22232\,
            I => \N__22007\
        );

    \I__5425\ : ClkMux
    port map (
            O => \N__22231\,
            I => \N__22007\
        );

    \I__5424\ : ClkMux
    port map (
            O => \N__22230\,
            I => \N__22007\
        );

    \I__5423\ : ClkMux
    port map (
            O => \N__22229\,
            I => \N__22007\
        );

    \I__5422\ : ClkMux
    port map (
            O => \N__22228\,
            I => \N__22007\
        );

    \I__5421\ : ClkMux
    port map (
            O => \N__22227\,
            I => \N__22007\
        );

    \I__5420\ : ClkMux
    port map (
            O => \N__22226\,
            I => \N__22007\
        );

    \I__5419\ : ClkMux
    port map (
            O => \N__22225\,
            I => \N__22007\
        );

    \I__5418\ : ClkMux
    port map (
            O => \N__22224\,
            I => \N__22007\
        );

    \I__5417\ : ClkMux
    port map (
            O => \N__22223\,
            I => \N__22007\
        );

    \I__5416\ : ClkMux
    port map (
            O => \N__22222\,
            I => \N__22007\
        );

    \I__5415\ : ClkMux
    port map (
            O => \N__22221\,
            I => \N__22007\
        );

    \I__5414\ : ClkMux
    port map (
            O => \N__22220\,
            I => \N__22007\
        );

    \I__5413\ : ClkMux
    port map (
            O => \N__22219\,
            I => \N__22007\
        );

    \I__5412\ : ClkMux
    port map (
            O => \N__22218\,
            I => \N__22007\
        );

    \I__5411\ : ClkMux
    port map (
            O => \N__22217\,
            I => \N__22007\
        );

    \I__5410\ : ClkMux
    port map (
            O => \N__22216\,
            I => \N__22007\
        );

    \I__5409\ : ClkMux
    port map (
            O => \N__22215\,
            I => \N__22007\
        );

    \I__5408\ : ClkMux
    port map (
            O => \N__22214\,
            I => \N__22007\
        );

    \I__5407\ : ClkMux
    port map (
            O => \N__22213\,
            I => \N__22007\
        );

    \I__5406\ : ClkMux
    port map (
            O => \N__22212\,
            I => \N__22007\
        );

    \I__5405\ : ClkMux
    port map (
            O => \N__22211\,
            I => \N__22007\
        );

    \I__5404\ : ClkMux
    port map (
            O => \N__22210\,
            I => \N__22007\
        );

    \I__5403\ : ClkMux
    port map (
            O => \N__22209\,
            I => \N__22007\
        );

    \I__5402\ : ClkMux
    port map (
            O => \N__22208\,
            I => \N__22007\
        );

    \I__5401\ : ClkMux
    port map (
            O => \N__22207\,
            I => \N__22007\
        );

    \I__5400\ : ClkMux
    port map (
            O => \N__22206\,
            I => \N__22007\
        );

    \I__5399\ : ClkMux
    port map (
            O => \N__22205\,
            I => \N__22007\
        );

    \I__5398\ : ClkMux
    port map (
            O => \N__22204\,
            I => \N__22007\
        );

    \I__5397\ : ClkMux
    port map (
            O => \N__22203\,
            I => \N__22007\
        );

    \I__5396\ : ClkMux
    port map (
            O => \N__22202\,
            I => \N__22007\
        );

    \I__5395\ : ClkMux
    port map (
            O => \N__22201\,
            I => \N__22007\
        );

    \I__5394\ : ClkMux
    port map (
            O => \N__22200\,
            I => \N__22007\
        );

    \I__5393\ : ClkMux
    port map (
            O => \N__22199\,
            I => \N__22007\
        );

    \I__5392\ : ClkMux
    port map (
            O => \N__22198\,
            I => \N__22007\
        );

    \I__5391\ : ClkMux
    port map (
            O => \N__22197\,
            I => \N__22007\
        );

    \I__5390\ : ClkMux
    port map (
            O => \N__22196\,
            I => \N__22007\
        );

    \I__5389\ : ClkMux
    port map (
            O => \N__22195\,
            I => \N__22007\
        );

    \I__5388\ : ClkMux
    port map (
            O => \N__22194\,
            I => \N__22007\
        );

    \I__5387\ : ClkMux
    port map (
            O => \N__22193\,
            I => \N__22007\
        );

    \I__5386\ : ClkMux
    port map (
            O => \N__22192\,
            I => \N__22007\
        );

    \I__5385\ : ClkMux
    port map (
            O => \N__22191\,
            I => \N__22007\
        );

    \I__5384\ : ClkMux
    port map (
            O => \N__22190\,
            I => \N__22007\
        );

    \I__5383\ : ClkMux
    port map (
            O => \N__22189\,
            I => \N__22007\
        );

    \I__5382\ : ClkMux
    port map (
            O => \N__22188\,
            I => \N__22007\
        );

    \I__5381\ : ClkMux
    port map (
            O => \N__22187\,
            I => \N__22007\
        );

    \I__5380\ : ClkMux
    port map (
            O => \N__22186\,
            I => \N__22007\
        );

    \I__5379\ : ClkMux
    port map (
            O => \N__22185\,
            I => \N__22007\
        );

    \I__5378\ : ClkMux
    port map (
            O => \N__22184\,
            I => \N__22007\
        );

    \I__5377\ : ClkMux
    port map (
            O => \N__22183\,
            I => \N__22007\
        );

    \I__5376\ : ClkMux
    port map (
            O => \N__22182\,
            I => \N__22007\
        );

    \I__5375\ : ClkMux
    port map (
            O => \N__22181\,
            I => \N__22007\
        );

    \I__5374\ : ClkMux
    port map (
            O => \N__22180\,
            I => \N__22007\
        );

    \I__5373\ : ClkMux
    port map (
            O => \N__22179\,
            I => \N__22007\
        );

    \I__5372\ : ClkMux
    port map (
            O => \N__22178\,
            I => \N__22007\
        );

    \I__5371\ : ClkMux
    port map (
            O => \N__22177\,
            I => \N__22007\
        );

    \I__5370\ : ClkMux
    port map (
            O => \N__22176\,
            I => \N__22007\
        );

    \I__5369\ : ClkMux
    port map (
            O => \N__22175\,
            I => \N__22007\
        );

    \I__5368\ : ClkMux
    port map (
            O => \N__22174\,
            I => \N__22007\
        );

    \I__5367\ : ClkMux
    port map (
            O => \N__22173\,
            I => \N__22007\
        );

    \I__5366\ : ClkMux
    port map (
            O => \N__22172\,
            I => \N__22007\
        );

    \I__5365\ : ClkMux
    port map (
            O => \N__22171\,
            I => \N__22007\
        );

    \I__5364\ : ClkMux
    port map (
            O => \N__22170\,
            I => \N__22007\
        );

    \I__5363\ : ClkMux
    port map (
            O => \N__22169\,
            I => \N__22007\
        );

    \I__5362\ : ClkMux
    port map (
            O => \N__22168\,
            I => \N__22007\
        );

    \I__5361\ : ClkMux
    port map (
            O => \N__22167\,
            I => \N__22007\
        );

    \I__5360\ : ClkMux
    port map (
            O => \N__22166\,
            I => \N__22007\
        );

    \I__5359\ : GlobalMux
    port map (
            O => \N__22007\,
            I => \N__22004\
        );

    \I__5358\ : gio2CtrlBuf
    port map (
            O => \N__22004\,
            I => clk_0_c_g
        );

    \I__5357\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21984\
        );

    \I__5356\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21981\
        );

    \I__5355\ : InMux
    port map (
            O => \N__21999\,
            I => \N__21976\
        );

    \I__5354\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21976\
        );

    \I__5353\ : InMux
    port map (
            O => \N__21997\,
            I => \N__21973\
        );

    \I__5352\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21970\
        );

    \I__5351\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21967\
        );

    \I__5350\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21964\
        );

    \I__5349\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21957\
        );

    \I__5348\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21957\
        );

    \I__5347\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21957\
        );

    \I__5346\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21954\
        );

    \I__5345\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21951\
        );

    \I__5344\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21946\
        );

    \I__5343\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21946\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__21984\,
            I => \N__21934\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__21981\,
            I => \N__21931\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__21976\,
            I => \N__21928\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__21973\,
            I => \N__21925\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__21970\,
            I => \N__21922\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__21967\,
            I => \N__21919\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__21964\,
            I => \N__21916\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__21957\,
            I => \N__21913\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__21954\,
            I => \N__21910\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__21951\,
            I => \N__21907\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__21946\,
            I => \N__21904\
        );

    \I__5331\ : SRMux
    port map (
            O => \N__21945\,
            I => \N__21863\
        );

    \I__5330\ : SRMux
    port map (
            O => \N__21944\,
            I => \N__21863\
        );

    \I__5329\ : SRMux
    port map (
            O => \N__21943\,
            I => \N__21863\
        );

    \I__5328\ : SRMux
    port map (
            O => \N__21942\,
            I => \N__21863\
        );

    \I__5327\ : SRMux
    port map (
            O => \N__21941\,
            I => \N__21863\
        );

    \I__5326\ : SRMux
    port map (
            O => \N__21940\,
            I => \N__21863\
        );

    \I__5325\ : SRMux
    port map (
            O => \N__21939\,
            I => \N__21863\
        );

    \I__5324\ : SRMux
    port map (
            O => \N__21938\,
            I => \N__21863\
        );

    \I__5323\ : SRMux
    port map (
            O => \N__21937\,
            I => \N__21863\
        );

    \I__5322\ : Glb2LocalMux
    port map (
            O => \N__21934\,
            I => \N__21863\
        );

    \I__5321\ : Glb2LocalMux
    port map (
            O => \N__21931\,
            I => \N__21863\
        );

    \I__5320\ : Glb2LocalMux
    port map (
            O => \N__21928\,
            I => \N__21863\
        );

    \I__5319\ : Glb2LocalMux
    port map (
            O => \N__21925\,
            I => \N__21863\
        );

    \I__5318\ : Glb2LocalMux
    port map (
            O => \N__21922\,
            I => \N__21863\
        );

    \I__5317\ : Glb2LocalMux
    port map (
            O => \N__21919\,
            I => \N__21863\
        );

    \I__5316\ : Glb2LocalMux
    port map (
            O => \N__21916\,
            I => \N__21863\
        );

    \I__5315\ : Glb2LocalMux
    port map (
            O => \N__21913\,
            I => \N__21863\
        );

    \I__5314\ : Glb2LocalMux
    port map (
            O => \N__21910\,
            I => \N__21863\
        );

    \I__5313\ : Glb2LocalMux
    port map (
            O => \N__21907\,
            I => \N__21863\
        );

    \I__5312\ : Glb2LocalMux
    port map (
            O => \N__21904\,
            I => \N__21863\
        );

    \I__5311\ : GlobalMux
    port map (
            O => \N__21863\,
            I => \N__21860\
        );

    \I__5310\ : gio2CtrlBuf
    port map (
            O => \N__21860\,
            I => \M_this_state_q_nss_g_0\
        );

    \I__5309\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__5307\ : Span12Mux_v
    port map (
            O => \N__21851\,
            I => \N__21848\
        );

    \I__5306\ : Odrv12
    port map (
            O => \N__21848\,
            I => port_address_in_3
        );

    \I__5305\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__21842\,
            I => port_address_in_4
        );

    \I__5303\ : CascadeMux
    port map (
            O => \N__21839\,
            I => \N__21836\
        );

    \I__5302\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21833\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__21833\,
            I => port_address_in_5
        );

    \I__5300\ : InMux
    port map (
            O => \N__21830\,
            I => \N__21827\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__21827\,
            I => \N__21824\
        );

    \I__5298\ : Span4Mux_s3_h
    port map (
            O => \N__21824\,
            I => \N__21821\
        );

    \I__5297\ : Span4Mux_v
    port map (
            O => \N__21821\,
            I => \N__21818\
        );

    \I__5296\ : Span4Mux_v
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__5295\ : IoSpan4Mux
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__5294\ : IoSpan4Mux
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__21809\,
            I => port_address_in_2
        );

    \I__5292\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__5288\ : Span4Mux_v
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__5287\ : Span4Mux_v
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__21785\,
            I => port_address_in_7
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__21782\,
            I => \M_this_state_d36_2_0_3_cascade_\
        );

    \I__5283\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__5281\ : Span12Mux_v
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__5280\ : Odrv12
    port map (
            O => \N__21770\,
            I => port_address_in_6
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__21767\,
            I => \N__21761\
        );

    \I__5278\ : CascadeMux
    port map (
            O => \N__21766\,
            I => \N__21758\
        );

    \I__5277\ : CascadeMux
    port map (
            O => \N__21765\,
            I => \N__21755\
        );

    \I__5276\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21752\
        );

    \I__5275\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21745\
        );

    \I__5274\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21745\
        );

    \I__5273\ : InMux
    port map (
            O => \N__21755\,
            I => \N__21745\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__21752\,
            I => \N__21740\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__21745\,
            I => \N__21740\
        );

    \I__5270\ : Span12Mux_h
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__5269\ : Odrv12
    port map (
            O => \N__21737\,
            I => \M_this_state_d37_1\
        );

    \I__5268\ : IoInMux
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__5266\ : Span12Mux_s2_h
    port map (
            O => \N__21728\,
            I => \N__21724\
        );

    \I__5265\ : InMux
    port map (
            O => \N__21727\,
            I => \N__21721\
        );

    \I__5264\ : Odrv12
    port map (
            O => \N__21724\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__21721\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__5262\ : InMux
    port map (
            O => \N__21716\,
            I => \un1_M_this_external_address_q_cry_5\
        );

    \I__5261\ : IoInMux
    port map (
            O => \N__21713\,
            I => \N__21710\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__21710\,
            I => \N__21707\
        );

    \I__5259\ : Span4Mux_s2_h
    port map (
            O => \N__21707\,
            I => \N__21704\
        );

    \I__5258\ : Sp12to4
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__5257\ : Span12Mux_v
    port map (
            O => \N__21701\,
            I => \N__21697\
        );

    \I__5256\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21694\
        );

    \I__5255\ : Odrv12
    port map (
            O => \N__21697\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__21694\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__5253\ : InMux
    port map (
            O => \N__21689\,
            I => \un1_M_this_external_address_q_cry_6\
        );

    \I__5252\ : IoInMux
    port map (
            O => \N__21686\,
            I => \N__21683\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__21683\,
            I => \N__21680\
        );

    \I__5250\ : IoSpan4Mux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__5249\ : Span4Mux_s0_v
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__5248\ : Sp12to4
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__5247\ : Span12Mux_v
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__5246\ : Span12Mux_h
    port map (
            O => \N__21668\,
            I => \N__21664\
        );

    \I__5245\ : InMux
    port map (
            O => \N__21667\,
            I => \N__21661\
        );

    \I__5244\ : Odrv12
    port map (
            O => \N__21664\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__21661\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__5242\ : InMux
    port map (
            O => \N__21656\,
            I => \bfn_30_24_0_\
        );

    \I__5241\ : IoInMux
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__5239\ : Span12Mux_s8_v
    port map (
            O => \N__21647\,
            I => \N__21643\
        );

    \I__5238\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21640\
        );

    \I__5237\ : Odrv12
    port map (
            O => \N__21643\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__21640\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__5235\ : InMux
    port map (
            O => \N__21635\,
            I => \un1_M_this_external_address_q_cry_8\
        );

    \I__5234\ : IoInMux
    port map (
            O => \N__21632\,
            I => \N__21629\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__21629\,
            I => \N__21626\
        );

    \I__5232\ : IoSpan4Mux
    port map (
            O => \N__21626\,
            I => \N__21623\
        );

    \I__5231\ : Span4Mux_s2_v
    port map (
            O => \N__21623\,
            I => \N__21620\
        );

    \I__5230\ : Sp12to4
    port map (
            O => \N__21620\,
            I => \N__21617\
        );

    \I__5229\ : Span12Mux_s8_v
    port map (
            O => \N__21617\,
            I => \N__21613\
        );

    \I__5228\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21610\
        );

    \I__5227\ : Odrv12
    port map (
            O => \N__21613\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__21610\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__5225\ : InMux
    port map (
            O => \N__21605\,
            I => \un1_M_this_external_address_q_cry_9\
        );

    \I__5224\ : IoInMux
    port map (
            O => \N__21602\,
            I => \N__21599\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__21599\,
            I => \N__21595\
        );

    \I__5222\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21592\
        );

    \I__5221\ : Odrv12
    port map (
            O => \N__21595\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__21592\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__5219\ : InMux
    port map (
            O => \N__21587\,
            I => \un1_M_this_external_address_q_cry_10\
        );

    \I__5218\ : IoInMux
    port map (
            O => \N__21584\,
            I => \N__21581\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__21581\,
            I => \N__21577\
        );

    \I__5216\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21574\
        );

    \I__5215\ : Odrv4
    port map (
            O => \N__21577\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__21574\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__5213\ : InMux
    port map (
            O => \N__21569\,
            I => \un1_M_this_external_address_q_cry_11\
        );

    \I__5212\ : IoInMux
    port map (
            O => \N__21566\,
            I => \N__21563\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__21563\,
            I => \N__21560\
        );

    \I__5210\ : IoSpan4Mux
    port map (
            O => \N__21560\,
            I => \N__21557\
        );

    \I__5209\ : Sp12to4
    port map (
            O => \N__21557\,
            I => \N__21553\
        );

    \I__5208\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21550\
        );

    \I__5207\ : Odrv12
    port map (
            O => \N__21553\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__21550\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__5205\ : InMux
    port map (
            O => \N__21545\,
            I => \un1_M_this_external_address_q_cry_12\
        );

    \I__5204\ : CascadeMux
    port map (
            O => \N__21542\,
            I => \N__21539\
        );

    \I__5203\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21535\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__21538\,
            I => \N__21532\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__21535\,
            I => \N__21528\
        );

    \I__5200\ : InMux
    port map (
            O => \N__21532\,
            I => \N__21525\
        );

    \I__5199\ : InMux
    port map (
            O => \N__21531\,
            I => \N__21522\
        );

    \I__5198\ : Span4Mux_h
    port map (
            O => \N__21528\,
            I => \N__21519\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__21525\,
            I => \N__21516\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__21522\,
            I => \N__21513\
        );

    \I__5195\ : Span4Mux_v
    port map (
            O => \N__21519\,
            I => \N__21510\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__21516\,
            I => \N__21507\
        );

    \I__5193\ : Span12Mux_h
    port map (
            O => \N__21513\,
            I => \N__21504\
        );

    \I__5192\ : Span4Mux_v
    port map (
            O => \N__21510\,
            I => \N__21501\
        );

    \I__5191\ : Span4Mux_v
    port map (
            O => \N__21507\,
            I => \N__21498\
        );

    \I__5190\ : Odrv12
    port map (
            O => \N__21504\,
            I => port_data_c_1
        );

    \I__5189\ : Odrv4
    port map (
            O => \N__21501\,
            I => port_data_c_1
        );

    \I__5188\ : Odrv4
    port map (
            O => \N__21498\,
            I => port_data_c_1
        );

    \I__5187\ : InMux
    port map (
            O => \N__21491\,
            I => \N__21483\
        );

    \I__5186\ : InMux
    port map (
            O => \N__21490\,
            I => \N__21483\
        );

    \I__5185\ : InMux
    port map (
            O => \N__21489\,
            I => \N__21478\
        );

    \I__5184\ : InMux
    port map (
            O => \N__21488\,
            I => \N__21478\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__21483\,
            I => \un1_M_this_state_q_2_0\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__21478\,
            I => \un1_M_this_state_q_2_0\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__21473\,
            I => \N__21469\
        );

    \I__5180\ : CascadeMux
    port map (
            O => \N__21472\,
            I => \N__21466\
        );

    \I__5179\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21462\
        );

    \I__5178\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21459\
        );

    \I__5177\ : CascadeMux
    port map (
            O => \N__21465\,
            I => \N__21456\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__21462\,
            I => \N__21451\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__21459\,
            I => \N__21451\
        );

    \I__5174\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21448\
        );

    \I__5173\ : Span4Mux_v
    port map (
            O => \N__21451\,
            I => \N__21445\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__21448\,
            I => \N__21442\
        );

    \I__5171\ : Sp12to4
    port map (
            O => \N__21445\,
            I => \N__21439\
        );

    \I__5170\ : Span4Mux_v
    port map (
            O => \N__21442\,
            I => \N__21436\
        );

    \I__5169\ : Span12Mux_h
    port map (
            O => \N__21439\,
            I => \N__21433\
        );

    \I__5168\ : Span4Mux_h
    port map (
            O => \N__21436\,
            I => \N__21430\
        );

    \I__5167\ : Odrv12
    port map (
            O => \N__21433\,
            I => port_data_c_5
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__21430\,
            I => port_data_c_5
        );

    \I__5165\ : InMux
    port map (
            O => \N__21425\,
            I => \N__21418\
        );

    \I__5164\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21418\
        );

    \I__5163\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21415\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__21418\,
            I => \M_this_sprites_ram_write_data_0_sqmuxa\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__21415\,
            I => \M_this_sprites_ram_write_data_0_sqmuxa\
        );

    \I__5160\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__21407\,
            I => \N__21403\
        );

    \I__5158\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21400\
        );

    \I__5157\ : Span4Mux_s2_v
    port map (
            O => \N__21403\,
            I => \N__21394\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__21400\,
            I => \N__21394\
        );

    \I__5155\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21391\
        );

    \I__5154\ : Span4Mux_v
    port map (
            O => \N__21394\,
            I => \N__21384\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__21391\,
            I => \N__21384\
        );

    \I__5152\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21381\
        );

    \I__5151\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21377\
        );

    \I__5150\ : Span4Mux_v
    port map (
            O => \N__21384\,
            I => \N__21371\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__21381\,
            I => \N__21371\
        );

    \I__5148\ : InMux
    port map (
            O => \N__21380\,
            I => \N__21368\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__21377\,
            I => \N__21364\
        );

    \I__5146\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21361\
        );

    \I__5145\ : Span4Mux_v
    port map (
            O => \N__21371\,
            I => \N__21356\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__21368\,
            I => \N__21356\
        );

    \I__5143\ : InMux
    port map (
            O => \N__21367\,
            I => \N__21353\
        );

    \I__5142\ : Span4Mux_v
    port map (
            O => \N__21364\,
            I => \N__21348\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__21361\,
            I => \N__21348\
        );

    \I__5140\ : Span4Mux_v
    port map (
            O => \N__21356\,
            I => \N__21343\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__21353\,
            I => \N__21343\
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__21348\,
            I => \M_this_sprites_ram_write_data_0_i_1\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__21343\,
            I => \M_this_sprites_ram_write_data_0_i_1\
        );

    \I__5136\ : InMux
    port map (
            O => \N__21338\,
            I => \N__21335\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__21335\,
            I => \N__21332\
        );

    \I__5134\ : Span4Mux_v
    port map (
            O => \N__21332\,
            I => \N__21328\
        );

    \I__5133\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21321\
        );

    \I__5132\ : Span4Mux_v
    port map (
            O => \N__21328\,
            I => \N__21317\
        );

    \I__5131\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21310\
        );

    \I__5130\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21310\
        );

    \I__5129\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21310\
        );

    \I__5128\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21307\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__21321\,
            I => \N__21304\
        );

    \I__5126\ : InMux
    port map (
            O => \N__21320\,
            I => \N__21301\
        );

    \I__5125\ : Span4Mux_v
    port map (
            O => \N__21317\,
            I => \N__21297\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__21310\,
            I => \N__21292\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21292\
        );

    \I__5122\ : Span4Mux_v
    port map (
            O => \N__21304\,
            I => \N__21289\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__21301\,
            I => \N__21286\
        );

    \I__5120\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21283\
        );

    \I__5119\ : Sp12to4
    port map (
            O => \N__21297\,
            I => \N__21270\
        );

    \I__5118\ : Span12Mux_v
    port map (
            O => \N__21292\,
            I => \N__21270\
        );

    \I__5117\ : Sp12to4
    port map (
            O => \N__21289\,
            I => \N__21270\
        );

    \I__5116\ : Span12Mux_s8_h
    port map (
            O => \N__21286\,
            I => \N__21270\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__21283\,
            I => \N__21270\
        );

    \I__5114\ : InMux
    port map (
            O => \N__21282\,
            I => \N__21265\
        );

    \I__5113\ : InMux
    port map (
            O => \N__21281\,
            I => \N__21265\
        );

    \I__5112\ : Odrv12
    port map (
            O => \N__21270\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__21265\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__5110\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21250\
        );

    \I__5109\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21250\
        );

    \I__5108\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21250\
        );

    \I__5107\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21244\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__21250\,
            I => \N__21241\
        );

    \I__5105\ : InMux
    port map (
            O => \N__21249\,
            I => \N__21238\
        );

    \I__5104\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21235\
        );

    \I__5103\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21231\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__21244\,
            I => \N__21228\
        );

    \I__5101\ : Span4Mux_h
    port map (
            O => \N__21241\,
            I => \N__21225\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21238\,
            I => \N__21222\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__21235\,
            I => \N__21219\
        );

    \I__5098\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21216\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__21231\,
            I => \N__21213\
        );

    \I__5096\ : Sp12to4
    port map (
            O => \N__21228\,
            I => \N__21210\
        );

    \I__5095\ : Span4Mux_v
    port map (
            O => \N__21225\,
            I => \N__21205\
        );

    \I__5094\ : Span4Mux_h
    port map (
            O => \N__21222\,
            I => \N__21205\
        );

    \I__5093\ : Span4Mux_v
    port map (
            O => \N__21219\,
            I => \N__21202\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__21216\,
            I => \N__21199\
        );

    \I__5091\ : Span4Mux_h
    port map (
            O => \N__21213\,
            I => \N__21196\
        );

    \I__5090\ : Odrv12
    port map (
            O => \N__21210\,
            I => \M_this_sprites_ram_write_en_1_0_0\
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__21205\,
            I => \M_this_sprites_ram_write_en_1_0_0\
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__21202\,
            I => \M_this_sprites_ram_write_en_1_0_0\
        );

    \I__5087\ : Odrv4
    port map (
            O => \N__21199\,
            I => \M_this_sprites_ram_write_en_1_0_0\
        );

    \I__5086\ : Odrv4
    port map (
            O => \N__21196\,
            I => \M_this_sprites_ram_write_en_1_0_0\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__21185\,
            I => \N__21179\
        );

    \I__5084\ : CascadeMux
    port map (
            O => \N__21184\,
            I => \N__21176\
        );

    \I__5083\ : CascadeMux
    port map (
            O => \N__21183\,
            I => \N__21172\
        );

    \I__5082\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21165\
        );

    \I__5081\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21165\
        );

    \I__5080\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21165\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__21175\,
            I => \N__21162\
        );

    \I__5078\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21157\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__21165\,
            I => \N__21153\
        );

    \I__5076\ : InMux
    port map (
            O => \N__21162\,
            I => \N__21150\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__21161\,
            I => \N__21147\
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__21160\,
            I => \N__21144\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__21157\,
            I => \N__21141\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__21156\,
            I => \N__21138\
        );

    \I__5071\ : Span4Mux_v
    port map (
            O => \N__21153\,
            I => \N__21133\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__21150\,
            I => \N__21133\
        );

    \I__5069\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21130\
        );

    \I__5068\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21127\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__21141\,
            I => \N__21124\
        );

    \I__5066\ : InMux
    port map (
            O => \N__21138\,
            I => \N__21121\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__21133\,
            I => \N__21116\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__21130\,
            I => \N__21116\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__21127\,
            I => \N__21113\
        );

    \I__5062\ : Span4Mux_v
    port map (
            O => \N__21124\,
            I => \N__21110\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__21121\,
            I => \N__21107\
        );

    \I__5060\ : Span4Mux_v
    port map (
            O => \N__21116\,
            I => \N__21101\
        );

    \I__5059\ : Span4Mux_v
    port map (
            O => \N__21113\,
            I => \N__21101\
        );

    \I__5058\ : Span4Mux_v
    port map (
            O => \N__21110\,
            I => \N__21096\
        );

    \I__5057\ : Span4Mux_v
    port map (
            O => \N__21107\,
            I => \N__21096\
        );

    \I__5056\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21093\
        );

    \I__5055\ : Sp12to4
    port map (
            O => \N__21101\,
            I => \N__21085\
        );

    \I__5054\ : Sp12to4
    port map (
            O => \N__21096\,
            I => \N__21085\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21093\,
            I => \N__21085\
        );

    \I__5052\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21082\
        );

    \I__5051\ : Odrv12
    port map (
            O => \N__21085\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__21082\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__5049\ : CascadeMux
    port map (
            O => \N__21077\,
            I => \N__21073\
        );

    \I__5048\ : InMux
    port map (
            O => \N__21076\,
            I => \N__21068\
        );

    \I__5047\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21061\
        );

    \I__5046\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21061\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21061\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__21068\,
            I => \N__21057\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__21061\,
            I => \N__21054\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21060\,
            I => \N__21051\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__21057\,
            I => \N__21047\
        );

    \I__5040\ : Span4Mux_v
    port map (
            O => \N__21054\,
            I => \N__21042\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__21051\,
            I => \N__21042\
        );

    \I__5038\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21039\
        );

    \I__5037\ : Span4Mux_v
    port map (
            O => \N__21047\,
            I => \N__21036\
        );

    \I__5036\ : Span4Mux_v
    port map (
            O => \N__21042\,
            I => \N__21031\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__21039\,
            I => \N__21031\
        );

    \I__5034\ : Span4Mux_v
    port map (
            O => \N__21036\,
            I => \N__21026\
        );

    \I__5033\ : Span4Mux_v
    port map (
            O => \N__21031\,
            I => \N__21023\
        );

    \I__5032\ : InMux
    port map (
            O => \N__21030\,
            I => \N__21020\
        );

    \I__5031\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21017\
        );

    \I__5030\ : Sp12to4
    port map (
            O => \N__21026\,
            I => \N__21006\
        );

    \I__5029\ : Sp12to4
    port map (
            O => \N__21023\,
            I => \N__21006\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__21020\,
            I => \N__21006\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__21017\,
            I => \N__21006\
        );

    \I__5026\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21003\
        );

    \I__5025\ : InMux
    port map (
            O => \N__21015\,
            I => \N__21000\
        );

    \I__5024\ : Odrv12
    port map (
            O => \N__21006\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__21003\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__21000\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__5021\ : CEMux
    port map (
            O => \N__20993\,
            I => \N__20990\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__20990\,
            I => \N__20986\
        );

    \I__5019\ : CEMux
    port map (
            O => \N__20989\,
            I => \N__20983\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__20986\,
            I => \N__20978\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__20983\,
            I => \N__20978\
        );

    \I__5016\ : Odrv4
    port map (
            O => \N__20978\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__5015\ : CascadeMux
    port map (
            O => \N__20975\,
            I => \N__20970\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__20974\,
            I => \N__20966\
        );

    \I__5013\ : CascadeMux
    port map (
            O => \N__20973\,
            I => \N__20963\
        );

    \I__5012\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20955\
        );

    \I__5011\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20949\
        );

    \I__5010\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20946\
        );

    \I__5009\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20943\
        );

    \I__5008\ : InMux
    port map (
            O => \N__20962\,
            I => \N__20938\
        );

    \I__5007\ : InMux
    port map (
            O => \N__20961\,
            I => \N__20938\
        );

    \I__5006\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20931\
        );

    \I__5005\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20931\
        );

    \I__5004\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20931\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__20955\,
            I => \N__20919\
        );

    \I__5002\ : InMux
    port map (
            O => \N__20954\,
            I => \N__20916\
        );

    \I__5001\ : InMux
    port map (
            O => \N__20953\,
            I => \N__20913\
        );

    \I__5000\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20910\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__20949\,
            I => \N__20907\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__20946\,
            I => \N__20904\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__20943\,
            I => \N__20897\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__20938\,
            I => \N__20897\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__20931\,
            I => \N__20897\
        );

    \I__4994\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20888\
        );

    \I__4993\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20888\
        );

    \I__4992\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20888\
        );

    \I__4991\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20888\
        );

    \I__4990\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20879\
        );

    \I__4989\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20879\
        );

    \I__4988\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20879\
        );

    \I__4987\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20879\
        );

    \I__4986\ : InMux
    port map (
            O => \N__20922\,
            I => \N__20876\
        );

    \I__4985\ : Span4Mux_h
    port map (
            O => \N__20919\,
            I => \N__20873\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__20916\,
            I => \N__20868\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__20913\,
            I => \N__20868\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__20910\,
            I => \N__20861\
        );

    \I__4981\ : Sp12to4
    port map (
            O => \N__20907\,
            I => \N__20861\
        );

    \I__4980\ : Span12Mux_s2_h
    port map (
            O => \N__20904\,
            I => \N__20861\
        );

    \I__4979\ : Span4Mux_v
    port map (
            O => \N__20897\,
            I => \N__20854\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__20888\,
            I => \N__20854\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20854\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__20876\,
            I => \N__20851\
        );

    \I__4975\ : Span4Mux_h
    port map (
            O => \N__20873\,
            I => \N__20846\
        );

    \I__4974\ : Span4Mux_h
    port map (
            O => \N__20868\,
            I => \N__20846\
        );

    \I__4973\ : Odrv12
    port map (
            O => \N__20861\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4972\ : Odrv4
    port map (
            O => \N__20854\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4971\ : Odrv12
    port map (
            O => \N__20851\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__20846\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4969\ : IoInMux
    port map (
            O => \N__20837\,
            I => \N__20834\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__4967\ : Span4Mux_s1_v
    port map (
            O => \N__20831\,
            I => \N__20828\
        );

    \I__4966\ : Sp12to4
    port map (
            O => \N__20828\,
            I => \N__20825\
        );

    \I__4965\ : Span12Mux_h
    port map (
            O => \N__20825\,
            I => \N__20821\
        );

    \I__4964\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20818\
        );

    \I__4963\ : Odrv12
    port map (
            O => \N__20821\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__20818\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__4961\ : IoInMux
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__4959\ : IoSpan4Mux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__4958\ : Sp12to4
    port map (
            O => \N__20804\,
            I => \N__20800\
        );

    \I__4957\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20797\
        );

    \I__4956\ : Odrv12
    port map (
            O => \N__20800\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__20797\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__4954\ : InMux
    port map (
            O => \N__20792\,
            I => \un1_M_this_external_address_q_cry_0\
        );

    \I__4953\ : IoInMux
    port map (
            O => \N__20789\,
            I => \N__20786\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__20786\,
            I => \N__20783\
        );

    \I__4951\ : IoSpan4Mux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__4950\ : IoSpan4Mux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__4949\ : Span4Mux_s2_v
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__4948\ : Span4Mux_v
    port map (
            O => \N__20774\,
            I => \N__20770\
        );

    \I__4947\ : InMux
    port map (
            O => \N__20773\,
            I => \N__20767\
        );

    \I__4946\ : Odrv4
    port map (
            O => \N__20770\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__20767\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__4944\ : InMux
    port map (
            O => \N__20762\,
            I => \un1_M_this_external_address_q_cry_1\
        );

    \I__4943\ : IoInMux
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__4941\ : Span4Mux_s2_h
    port map (
            O => \N__20753\,
            I => \N__20750\
        );

    \I__4940\ : Span4Mux_v
    port map (
            O => \N__20750\,
            I => \N__20746\
        );

    \I__4939\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20743\
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__20746\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__20743\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__4936\ : InMux
    port map (
            O => \N__20738\,
            I => \un1_M_this_external_address_q_cry_2\
        );

    \I__4935\ : IoInMux
    port map (
            O => \N__20735\,
            I => \N__20732\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__20732\,
            I => \N__20728\
        );

    \I__4933\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20725\
        );

    \I__4932\ : Odrv4
    port map (
            O => \N__20728\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__20725\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__4930\ : InMux
    port map (
            O => \N__20720\,
            I => \un1_M_this_external_address_q_cry_3\
        );

    \I__4929\ : IoInMux
    port map (
            O => \N__20717\,
            I => \N__20714\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__4927\ : Span4Mux_s2_h
    port map (
            O => \N__20711\,
            I => \N__20707\
        );

    \I__4926\ : InMux
    port map (
            O => \N__20710\,
            I => \N__20704\
        );

    \I__4925\ : Odrv4
    port map (
            O => \N__20707\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__20704\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__4923\ : InMux
    port map (
            O => \N__20699\,
            I => \un1_M_this_external_address_q_cry_4\
        );

    \I__4922\ : InMux
    port map (
            O => \N__20696\,
            I => \N__20693\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__20693\,
            I => \N__20690\
        );

    \I__4920\ : Sp12to4
    port map (
            O => \N__20690\,
            I => \N__20687\
        );

    \I__4919\ : Odrv12
    port map (
            O => \N__20687\,
            I => \this_sprites_ram.mem_out_bus5_2\
        );

    \I__4918\ : CascadeMux
    port map (
            O => \N__20684\,
            I => \N__20679\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__20683\,
            I => \N__20675\
        );

    \I__4916\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20667\
        );

    \I__4915\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20667\
        );

    \I__4914\ : CascadeMux
    port map (
            O => \N__20678\,
            I => \N__20664\
        );

    \I__4913\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20661\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__20674\,
            I => \N__20658\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__20673\,
            I => \N__20654\
        );

    \I__4910\ : CascadeMux
    port map (
            O => \N__20672\,
            I => \N__20651\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__20667\,
            I => \N__20648\
        );

    \I__4908\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20645\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__20661\,
            I => \N__20642\
        );

    \I__4906\ : InMux
    port map (
            O => \N__20658\,
            I => \N__20639\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__20657\,
            I => \N__20636\
        );

    \I__4904\ : InMux
    port map (
            O => \N__20654\,
            I => \N__20633\
        );

    \I__4903\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20630\
        );

    \I__4902\ : Span4Mux_v
    port map (
            O => \N__20648\,
            I => \N__20625\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__20645\,
            I => \N__20625\
        );

    \I__4900\ : Span4Mux_v
    port map (
            O => \N__20642\,
            I => \N__20620\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__20639\,
            I => \N__20620\
        );

    \I__4898\ : InMux
    port map (
            O => \N__20636\,
            I => \N__20617\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__20633\,
            I => \N__20614\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__20630\,
            I => \N__20611\
        );

    \I__4895\ : Span4Mux_v
    port map (
            O => \N__20625\,
            I => \N__20608\
        );

    \I__4894\ : Span4Mux_v
    port map (
            O => \N__20620\,
            I => \N__20605\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__20617\,
            I => \N__20602\
        );

    \I__4892\ : Span12Mux_s11_h
    port map (
            O => \N__20614\,
            I => \N__20597\
        );

    \I__4891\ : Sp12to4
    port map (
            O => \N__20611\,
            I => \N__20597\
        );

    \I__4890\ : Odrv4
    port map (
            O => \N__20608\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__20605\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__4888\ : Odrv4
    port map (
            O => \N__20602\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__4887\ : Odrv12
    port map (
            O => \N__20597\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__4886\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20585\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__20585\,
            I => \N__20582\
        );

    \I__4884\ : Span4Mux_v
    port map (
            O => \N__20582\,
            I => \N__20579\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__20579\,
            I => \this_sprites_ram.mem_out_bus1_2\
        );

    \I__4882\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20573\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__20573\,
            I => \N__20570\
        );

    \I__4880\ : Sp12to4
    port map (
            O => \N__20570\,
            I => \N__20567\
        );

    \I__4879\ : Span12Mux_v
    port map (
            O => \N__20567\,
            I => \N__20564\
        );

    \I__4878\ : Odrv12
    port map (
            O => \N__20564\,
            I => \this_sprites_ram.mem_out_bus7_2\
        );

    \I__4877\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20558\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__20558\,
            I => \this_sprites_ram.mem_out_bus3_2\
        );

    \I__4875\ : CascadeMux
    port map (
            O => \N__20555\,
            I => \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_2_cascade_\
        );

    \I__4874\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20537\
        );

    \I__4873\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20537\
        );

    \I__4872\ : InMux
    port map (
            O => \N__20550\,
            I => \N__20537\
        );

    \I__4871\ : InMux
    port map (
            O => \N__20549\,
            I => \N__20537\
        );

    \I__4870\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20525\
        );

    \I__4869\ : InMux
    port map (
            O => \N__20547\,
            I => \N__20525\
        );

    \I__4868\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20522\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__20537\,
            I => \N__20519\
        );

    \I__4866\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20514\
        );

    \I__4865\ : InMux
    port map (
            O => \N__20535\,
            I => \N__20514\
        );

    \I__4864\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20511\
        );

    \I__4863\ : InMux
    port map (
            O => \N__20533\,
            I => \N__20506\
        );

    \I__4862\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20506\
        );

    \I__4861\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20503\
        );

    \I__4860\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20500\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__20525\,
            I => \N__20497\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__20522\,
            I => \N__20488\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__20519\,
            I => \N__20488\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__20514\,
            I => \N__20488\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__20511\,
            I => \N__20481\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__20506\,
            I => \N__20481\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__20503\,
            I => \N__20481\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__20500\,
            I => \N__20476\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__20497\,
            I => \N__20476\
        );

    \I__4850\ : InMux
    port map (
            O => \N__20496\,
            I => \N__20473\
        );

    \I__4849\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20470\
        );

    \I__4848\ : Span4Mux_v
    port map (
            O => \N__20488\,
            I => \N__20467\
        );

    \I__4847\ : Span4Mux_h
    port map (
            O => \N__20481\,
            I => \N__20464\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__20476\,
            I => \N__20459\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__20473\,
            I => \N__20459\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__20470\,
            I => \N__20456\
        );

    \I__4843\ : Odrv4
    port map (
            O => \N__20467\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4842\ : Odrv4
    port map (
            O => \N__20464\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__20459\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4840\ : Odrv12
    port map (
            O => \N__20456\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4839\ : InMux
    port map (
            O => \N__20447\,
            I => \N__20444\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__20444\,
            I => \N__20441\
        );

    \I__4837\ : Span4Mux_v
    port map (
            O => \N__20441\,
            I => \N__20438\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__20438\,
            I => \this_sprites_ram_mem_N_95\
        );

    \I__4835\ : CEMux
    port map (
            O => \N__20435\,
            I => \N__20432\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__20432\,
            I => \N__20428\
        );

    \I__4833\ : CEMux
    port map (
            O => \N__20431\,
            I => \N__20425\
        );

    \I__4832\ : Span4Mux_h
    port map (
            O => \N__20428\,
            I => \N__20422\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__20425\,
            I => \N__20419\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__20422\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__4829\ : Odrv12
    port map (
            O => \N__20419\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__4828\ : CEMux
    port map (
            O => \N__20414\,
            I => \N__20410\
        );

    \I__4827\ : CEMux
    port map (
            O => \N__20413\,
            I => \N__20407\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__20410\,
            I => \N__20404\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__20407\,
            I => \N__20401\
        );

    \I__4824\ : Span4Mux_h
    port map (
            O => \N__20404\,
            I => \N__20398\
        );

    \I__4823\ : Span4Mux_h
    port map (
            O => \N__20401\,
            I => \N__20395\
        );

    \I__4822\ : Odrv4
    port map (
            O => \N__20398\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__4821\ : Odrv4
    port map (
            O => \N__20395\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__4820\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20384\
        );

    \I__4819\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20381\
        );

    \I__4818\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20378\
        );

    \I__4817\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20374\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__20384\,
            I => \N__20370\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__20381\,
            I => \N__20365\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__20378\,
            I => \N__20365\
        );

    \I__4813\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20362\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__20374\,
            I => \N__20359\
        );

    \I__4811\ : InMux
    port map (
            O => \N__20373\,
            I => \N__20356\
        );

    \I__4810\ : Span4Mux_h
    port map (
            O => \N__20370\,
            I => \N__20353\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__20365\,
            I => \N__20350\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__20362\,
            I => \N__20343\
        );

    \I__4807\ : Span12Mux_s8_h
    port map (
            O => \N__20359\,
            I => \N__20343\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__20356\,
            I => \N__20343\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__20353\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4804\ : Odrv4
    port map (
            O => \N__20350\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4803\ : Odrv12
    port map (
            O => \N__20343\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__20336\,
            I => \N__20332\
        );

    \I__4801\ : InMux
    port map (
            O => \N__20335\,
            I => \N__20328\
        );

    \I__4800\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20318\
        );

    \I__4799\ : InMux
    port map (
            O => \N__20331\,
            I => \N__20315\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__20328\,
            I => \N__20312\
        );

    \I__4797\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20309\
        );

    \I__4796\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20306\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20303\
        );

    \I__4794\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20298\
        );

    \I__4793\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20298\
        );

    \I__4792\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20295\
        );

    \I__4791\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20292\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__20318\,
            I => \N__20283\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__20315\,
            I => \N__20270\
        );

    \I__4788\ : Span4Mux_v
    port map (
            O => \N__20312\,
            I => \N__20270\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__20309\,
            I => \N__20270\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__20306\,
            I => \N__20270\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__20303\,
            I => \N__20270\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__20298\,
            I => \N__20263\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__20295\,
            I => \N__20263\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__20292\,
            I => \N__20263\
        );

    \I__4781\ : InMux
    port map (
            O => \N__20291\,
            I => \N__20259\
        );

    \I__4780\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20251\
        );

    \I__4779\ : InMux
    port map (
            O => \N__20289\,
            I => \N__20244\
        );

    \I__4778\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20244\
        );

    \I__4777\ : InMux
    port map (
            O => \N__20287\,
            I => \N__20244\
        );

    \I__4776\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20241\
        );

    \I__4775\ : Span4Mux_v
    port map (
            O => \N__20283\,
            I => \N__20238\
        );

    \I__4774\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20235\
        );

    \I__4773\ : InMux
    port map (
            O => \N__20281\,
            I => \N__20232\
        );

    \I__4772\ : Span4Mux_v
    port map (
            O => \N__20270\,
            I => \N__20227\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__20263\,
            I => \N__20227\
        );

    \I__4770\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20224\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__20259\,
            I => \N__20221\
        );

    \I__4768\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20216\
        );

    \I__4767\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20216\
        );

    \I__4766\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20213\
        );

    \I__4765\ : InMux
    port map (
            O => \N__20255\,
            I => \N__20208\
        );

    \I__4764\ : InMux
    port map (
            O => \N__20254\,
            I => \N__20208\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__20251\,
            I => \N__20205\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__20244\,
            I => \N__20202\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__20241\,
            I => \N__20185\
        );

    \I__4760\ : Sp12to4
    port map (
            O => \N__20238\,
            I => \N__20185\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__20235\,
            I => \N__20185\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__20232\,
            I => \N__20185\
        );

    \I__4757\ : Sp12to4
    port map (
            O => \N__20227\,
            I => \N__20185\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__20224\,
            I => \N__20185\
        );

    \I__4755\ : Sp12to4
    port map (
            O => \N__20221\,
            I => \N__20185\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__20216\,
            I => \N__20185\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__20213\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__20208\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__20205\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4750\ : Odrv4
    port map (
            O => \N__20202\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4749\ : Odrv12
    port map (
            O => \N__20185\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__20174\,
            I => \N__20170\
        );

    \I__4747\ : InMux
    port map (
            O => \N__20173\,
            I => \N__20167\
        );

    \I__4746\ : InMux
    port map (
            O => \N__20170\,
            I => \N__20164\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__20167\,
            I => \N__20160\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__20164\,
            I => \N__20157\
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__20163\,
            I => \N__20154\
        );

    \I__4742\ : Span4Mux_v
    port map (
            O => \N__20160\,
            I => \N__20151\
        );

    \I__4741\ : Span4Mux_v
    port map (
            O => \N__20157\,
            I => \N__20148\
        );

    \I__4740\ : InMux
    port map (
            O => \N__20154\,
            I => \N__20145\
        );

    \I__4739\ : Sp12to4
    port map (
            O => \N__20151\,
            I => \N__20142\
        );

    \I__4738\ : Span4Mux_h
    port map (
            O => \N__20148\,
            I => \N__20137\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__20145\,
            I => \N__20137\
        );

    \I__4736\ : Span12Mux_h
    port map (
            O => \N__20142\,
            I => \N__20134\
        );

    \I__4735\ : Span4Mux_h
    port map (
            O => \N__20137\,
            I => \N__20131\
        );

    \I__4734\ : Span12Mux_v
    port map (
            O => \N__20134\,
            I => \N__20128\
        );

    \I__4733\ : Sp12to4
    port map (
            O => \N__20131\,
            I => \N__20125\
        );

    \I__4732\ : Odrv12
    port map (
            O => \N__20128\,
            I => port_data_c_0
        );

    \I__4731\ : Odrv12
    port map (
            O => \N__20125\,
            I => port_data_c_0
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__20120\,
            I => \N__20115\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__20119\,
            I => \N__20112\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20109\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20115\,
            I => \N__20106\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20112\,
            I => \N__20103\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__20109\,
            I => \N__20100\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__20106\,
            I => \N__20095\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__20103\,
            I => \N__20095\
        );

    \I__4722\ : Span4Mux_v
    port map (
            O => \N__20100\,
            I => \N__20092\
        );

    \I__4721\ : Span12Mux_v
    port map (
            O => \N__20095\,
            I => \N__20089\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__20092\,
            I => \N__20086\
        );

    \I__4719\ : Span12Mux_h
    port map (
            O => \N__20089\,
            I => \N__20083\
        );

    \I__4718\ : IoSpan4Mux
    port map (
            O => \N__20086\,
            I => \N__20080\
        );

    \I__4717\ : Odrv12
    port map (
            O => \N__20083\,
            I => port_data_c_4
        );

    \I__4716\ : Odrv4
    port map (
            O => \N__20080\,
            I => port_data_c_4
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__20075\,
            I => \M_this_sprites_ram_write_data_0_sqmuxa_cascade_\
        );

    \I__4714\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20069\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__20069\,
            I => \N__20065\
        );

    \I__4712\ : InMux
    port map (
            O => \N__20068\,
            I => \N__20062\
        );

    \I__4711\ : Span4Mux_h
    port map (
            O => \N__20065\,
            I => \N__20058\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__20062\,
            I => \N__20055\
        );

    \I__4709\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20052\
        );

    \I__4708\ : Span4Mux_v
    port map (
            O => \N__20058\,
            I => \N__20045\
        );

    \I__4707\ : Span4Mux_h
    port map (
            O => \N__20055\,
            I => \N__20045\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__20052\,
            I => \N__20042\
        );

    \I__4705\ : InMux
    port map (
            O => \N__20051\,
            I => \N__20039\
        );

    \I__4704\ : InMux
    port map (
            O => \N__20050\,
            I => \N__20035\
        );

    \I__4703\ : Span4Mux_v
    port map (
            O => \N__20045\,
            I => \N__20029\
        );

    \I__4702\ : Span4Mux_h
    port map (
            O => \N__20042\,
            I => \N__20029\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__20039\,
            I => \N__20026\
        );

    \I__4700\ : InMux
    port map (
            O => \N__20038\,
            I => \N__20023\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__20035\,
            I => \N__20020\
        );

    \I__4698\ : InMux
    port map (
            O => \N__20034\,
            I => \N__20017\
        );

    \I__4697\ : Span4Mux_v
    port map (
            O => \N__20029\,
            I => \N__20012\
        );

    \I__4696\ : Span4Mux_h
    port map (
            O => \N__20026\,
            I => \N__20012\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__20023\,
            I => \N__20009\
        );

    \I__4694\ : Span4Mux_v
    port map (
            O => \N__20020\,
            I => \N__20004\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__20017\,
            I => \N__20004\
        );

    \I__4692\ : Span4Mux_v
    port map (
            O => \N__20012\,
            I => \N__19998\
        );

    \I__4691\ : Span4Mux_h
    port map (
            O => \N__20009\,
            I => \N__19998\
        );

    \I__4690\ : Span4Mux_v
    port map (
            O => \N__20004\,
            I => \N__19995\
        );

    \I__4689\ : InMux
    port map (
            O => \N__20003\,
            I => \N__19992\
        );

    \I__4688\ : Odrv4
    port map (
            O => \N__19998\,
            I => \M_this_sprites_ram_write_data_0_i_0\
        );

    \I__4687\ : Odrv4
    port map (
            O => \N__19995\,
            I => \M_this_sprites_ram_write_data_0_i_0\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__19992\,
            I => \M_this_sprites_ram_write_data_0_i_0\
        );

    \I__4685\ : CascadeMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__4684\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19979\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__19979\,
            I => \N__19975\
        );

    \I__4682\ : InMux
    port map (
            O => \N__19978\,
            I => \N__19972\
        );

    \I__4681\ : Span4Mux_v
    port map (
            O => \N__19975\,
            I => \N__19968\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__19972\,
            I => \N__19965\
        );

    \I__4679\ : InMux
    port map (
            O => \N__19971\,
            I => \N__19962\
        );

    \I__4678\ : Span4Mux_h
    port map (
            O => \N__19968\,
            I => \N__19957\
        );

    \I__4677\ : Span4Mux_v
    port map (
            O => \N__19965\,
            I => \N__19957\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__19962\,
            I => \N__19954\
        );

    \I__4675\ : Span4Mux_v
    port map (
            O => \N__19957\,
            I => \N__19951\
        );

    \I__4674\ : Span12Mux_h
    port map (
            O => \N__19954\,
            I => \N__19948\
        );

    \I__4673\ : Span4Mux_h
    port map (
            O => \N__19951\,
            I => \N__19945\
        );

    \I__4672\ : Odrv12
    port map (
            O => \N__19948\,
            I => port_data_c_3
        );

    \I__4671\ : Odrv4
    port map (
            O => \N__19945\,
            I => port_data_c_3
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__4669\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__4667\ : Span12Mux_h
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__4666\ : Span12Mux_v
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__4665\ : Odrv12
    port map (
            O => \N__19925\,
            I => port_data_c_7
        );

    \I__4664\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19915\
        );

    \I__4662\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19912\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__19915\,
            I => \N__19906\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__19912\,
            I => \N__19906\
        );

    \I__4659\ : InMux
    port map (
            O => \N__19911\,
            I => \N__19903\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__19906\,
            I => \N__19896\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__19903\,
            I => \N__19896\
        );

    \I__4656\ : InMux
    port map (
            O => \N__19902\,
            I => \N__19893\
        );

    \I__4655\ : InMux
    port map (
            O => \N__19901\,
            I => \N__19890\
        );

    \I__4654\ : Span4Mux_v
    port map (
            O => \N__19896\,
            I => \N__19883\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__19893\,
            I => \N__19883\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__19890\,
            I => \N__19880\
        );

    \I__4651\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19877\
        );

    \I__4650\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19874\
        );

    \I__4649\ : Span4Mux_v
    port map (
            O => \N__19883\,
            I => \N__19871\
        );

    \I__4648\ : Span4Mux_s3_v
    port map (
            O => \N__19880\,
            I => \N__19866\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19866\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__19874\,
            I => \N__19863\
        );

    \I__4645\ : Span4Mux_v
    port map (
            O => \N__19871\,
            I => \N__19857\
        );

    \I__4644\ : Span4Mux_v
    port map (
            O => \N__19866\,
            I => \N__19857\
        );

    \I__4643\ : Span4Mux_h
    port map (
            O => \N__19863\,
            I => \N__19854\
        );

    \I__4642\ : InMux
    port map (
            O => \N__19862\,
            I => \N__19851\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__19857\,
            I => \M_this_sprites_ram_write_data_0_i_3\
        );

    \I__4640\ : Odrv4
    port map (
            O => \N__19854\,
            I => \M_this_sprites_ram_write_data_0_i_3\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__19851\,
            I => \M_this_sprites_ram_write_data_0_i_3\
        );

    \I__4638\ : CascadeMux
    port map (
            O => \N__19844\,
            I => \N__19840\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__19843\,
            I => \N__19837\
        );

    \I__4636\ : InMux
    port map (
            O => \N__19840\,
            I => \N__19834\
        );

    \I__4635\ : InMux
    port map (
            O => \N__19837\,
            I => \N__19831\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__19834\,
            I => \N__19828\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__19831\,
            I => \N__19824\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__19828\,
            I => \N__19821\
        );

    \I__4631\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19818\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__19824\,
            I => \N__19815\
        );

    \I__4629\ : Span4Mux_h
    port map (
            O => \N__19821\,
            I => \N__19810\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__19818\,
            I => \N__19810\
        );

    \I__4627\ : Sp12to4
    port map (
            O => \N__19815\,
            I => \N__19807\
        );

    \I__4626\ : Span4Mux_h
    port map (
            O => \N__19810\,
            I => \N__19804\
        );

    \I__4625\ : Span12Mux_h
    port map (
            O => \N__19807\,
            I => \N__19799\
        );

    \I__4624\ : Sp12to4
    port map (
            O => \N__19804\,
            I => \N__19799\
        );

    \I__4623\ : Odrv12
    port map (
            O => \N__19799\,
            I => port_data_c_2
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__19796\,
            I => \N__19792\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__19795\,
            I => \N__19789\
        );

    \I__4620\ : InMux
    port map (
            O => \N__19792\,
            I => \N__19785\
        );

    \I__4619\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19782\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__19788\,
            I => \N__19779\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__19785\,
            I => \N__19776\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__19782\,
            I => \N__19773\
        );

    \I__4615\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19770\
        );

    \I__4614\ : Span12Mux_v
    port map (
            O => \N__19776\,
            I => \N__19767\
        );

    \I__4613\ : Span12Mux_h
    port map (
            O => \N__19773\,
            I => \N__19764\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__19770\,
            I => \N__19761\
        );

    \I__4611\ : Span12Mux_h
    port map (
            O => \N__19767\,
            I => \N__19756\
        );

    \I__4610\ : Span12Mux_v
    port map (
            O => \N__19764\,
            I => \N__19756\
        );

    \I__4609\ : Span12Mux_v
    port map (
            O => \N__19761\,
            I => \N__19753\
        );

    \I__4608\ : Odrv12
    port map (
            O => \N__19756\,
            I => port_data_c_6
        );

    \I__4607\ : Odrv12
    port map (
            O => \N__19753\,
            I => port_data_c_6
        );

    \I__4606\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__19745\,
            I => \N__19740\
        );

    \I__4604\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19737\
        );

    \I__4603\ : InMux
    port map (
            O => \N__19743\,
            I => \N__19733\
        );

    \I__4602\ : Span4Mux_v
    port map (
            O => \N__19740\,
            I => \N__19727\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__19737\,
            I => \N__19727\
        );

    \I__4600\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19724\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__19733\,
            I => \N__19720\
        );

    \I__4598\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19717\
        );

    \I__4597\ : Span4Mux_v
    port map (
            O => \N__19727\,
            I => \N__19712\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__19724\,
            I => \N__19712\
        );

    \I__4595\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19709\
        );

    \I__4594\ : Span4Mux_s3_v
    port map (
            O => \N__19720\,
            I => \N__19703\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19703\
        );

    \I__4592\ : Span4Mux_v
    port map (
            O => \N__19712\,
            I => \N__19698\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__19709\,
            I => \N__19698\
        );

    \I__4590\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19695\
        );

    \I__4589\ : Span4Mux_v
    port map (
            O => \N__19703\,
            I => \N__19691\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__19698\,
            I => \N__19686\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__19695\,
            I => \N__19686\
        );

    \I__4586\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19683\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__19691\,
            I => \M_this_sprites_ram_write_data_0_i_2\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__19686\,
            I => \M_this_sprites_ram_write_data_0_i_2\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__19683\,
            I => \M_this_sprites_ram_write_data_0_i_2\
        );

    \I__4582\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__4580\ : Span4Mux_v
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__4579\ : Span4Mux_v
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__4578\ : Odrv4
    port map (
            O => \N__19664\,
            I => \this_sprites_ram.mem_out_bus4_2\
        );

    \I__4577\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__4575\ : Span4Mux_v
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__4574\ : Odrv4
    port map (
            O => \N__19652\,
            I => \this_sprites_ram.mem_out_bus0_2\
        );

    \I__4573\ : InMux
    port map (
            O => \N__19649\,
            I => \N__19646\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__4571\ : Span4Mux_h
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__4570\ : Sp12to4
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__4569\ : Span12Mux_v
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__4568\ : Odrv12
    port map (
            O => \N__19634\,
            I => \this_sprites_ram.mem_out_bus6_2\
        );

    \I__4567\ : InMux
    port map (
            O => \N__19631\,
            I => \N__19628\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__19628\,
            I => \N__19625\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__19625\,
            I => \this_sprites_ram.mem_out_bus2_2\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__19622\,
            I => \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_2_cascade_\
        );

    \I__4563\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__19616\,
            I => \this_sprites_ram_mem_N_98\
        );

    \I__4561\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__4559\ : Span4Mux_v
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__4558\ : Span4Mux_v
    port map (
            O => \N__19604\,
            I => \N__19601\
        );

    \I__4557\ : Odrv4
    port map (
            O => \N__19601\,
            I => \this_sprites_ram.mem_out_bus5_0\
        );

    \I__4556\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__4554\ : Span4Mux_v
    port map (
            O => \N__19592\,
            I => \N__19589\
        );

    \I__4553\ : Odrv4
    port map (
            O => \N__19589\,
            I => \this_sprites_ram.mem_out_bus1_0\
        );

    \I__4552\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19583\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__19583\,
            I => \N__19580\
        );

    \I__4550\ : Odrv4
    port map (
            O => \N__19580\,
            I => \this_sprites_ram.mem_out_bus3_0\
        );

    \I__4549\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19574\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__19574\,
            I => \N__19571\
        );

    \I__4547\ : Span4Mux_v
    port map (
            O => \N__19571\,
            I => \N__19568\
        );

    \I__4546\ : Sp12to4
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__4545\ : Span12Mux_v
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__4544\ : Odrv12
    port map (
            O => \N__19562\,
            I => \this_sprites_ram.mem_out_bus7_0\
        );

    \I__4543\ : CascadeMux
    port map (
            O => \N__19559\,
            I => \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_0_cascade_\
        );

    \I__4542\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__19553\,
            I => \this_sprites_ram_mem_N_109\
        );

    \I__4540\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__19547\,
            I => \N__19544\
        );

    \I__4538\ : Span4Mux_v
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__4537\ : Span4Mux_v
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__4536\ : Odrv4
    port map (
            O => \N__19538\,
            I => \this_sprites_ram.mem_out_bus0_0\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__4534\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19529\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__19529\,
            I => \N__19526\
        );

    \I__4532\ : Span4Mux_v
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__4531\ : Span4Mux_h
    port map (
            O => \N__19523\,
            I => \N__19520\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__19520\,
            I => \this_sprites_ram.mem_out_bus4_0\
        );

    \I__4529\ : InMux
    port map (
            O => \N__19517\,
            I => \N__19514\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__4527\ : Sp12to4
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__4526\ : Span12Mux_v
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__4525\ : Odrv12
    port map (
            O => \N__19505\,
            I => \this_sprites_ram.mem_out_bus6_0\
        );

    \I__4524\ : CascadeMux
    port map (
            O => \N__19502\,
            I => \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_0_cascade_\
        );

    \I__4523\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__19496\,
            I => \this_sprites_ram.mem_out_bus2_0\
        );

    \I__4521\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__19490\,
            I => \this_sprites_ram_mem_N_112\
        );

    \I__4519\ : CEMux
    port map (
            O => \N__19487\,
            I => \N__19483\
        );

    \I__4518\ : CEMux
    port map (
            O => \N__19486\,
            I => \N__19480\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__19483\,
            I => \N__19477\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__19480\,
            I => \N__19474\
        );

    \I__4515\ : Span12Mux_s8_h
    port map (
            O => \N__19477\,
            I => \N__19471\
        );

    \I__4514\ : Span4Mux_h
    port map (
            O => \N__19474\,
            I => \N__19468\
        );

    \I__4513\ : Odrv12
    port map (
            O => \N__19471\,
            I => \this_sprites_ram.mem_WE_10\
        );

    \I__4512\ : Odrv4
    port map (
            O => \N__19468\,
            I => \this_sprites_ram.mem_WE_10\
        );

    \I__4511\ : CEMux
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__19460\,
            I => \N__19456\
        );

    \I__4509\ : CEMux
    port map (
            O => \N__19459\,
            I => \N__19453\
        );

    \I__4508\ : Span4Mux_v
    port map (
            O => \N__19456\,
            I => \N__19448\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__19453\,
            I => \N__19448\
        );

    \I__4506\ : Odrv4
    port map (
            O => \N__19448\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__4505\ : CEMux
    port map (
            O => \N__19445\,
            I => \N__19442\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__19442\,
            I => \N__19438\
        );

    \I__4503\ : CEMux
    port map (
            O => \N__19441\,
            I => \N__19435\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__19438\,
            I => \N__19430\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19435\,
            I => \N__19430\
        );

    \I__4500\ : Span4Mux_v
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__4499\ : Span4Mux_h
    port map (
            O => \N__19427\,
            I => \N__19424\
        );

    \I__4498\ : Odrv4
    port map (
            O => \N__19424\,
            I => \this_sprites_ram.mem_WE_12\
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__19421\,
            I => \N__19418\
        );

    \I__4496\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__19415\,
            I => \N__19412\
        );

    \I__4494\ : Odrv12
    port map (
            O => \N__19412\,
            I => \N_200\
        );

    \I__4493\ : InMux
    port map (
            O => \N__19409\,
            I => \N__19406\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__19406\,
            I => \N__19403\
        );

    \I__4491\ : Span4Mux_v
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__4490\ : Sp12to4
    port map (
            O => \N__19400\,
            I => \N__19397\
        );

    \I__4489\ : Span12Mux_h
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__4488\ : Odrv12
    port map (
            O => \N__19394\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__4487\ : InMux
    port map (
            O => \N__19391\,
            I => \N__19388\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__19388\,
            I => \N__19382\
        );

    \I__4485\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19379\
        );

    \I__4484\ : CEMux
    port map (
            O => \N__19386\,
            I => \N__19375\
        );

    \I__4483\ : CascadeMux
    port map (
            O => \N__19385\,
            I => \N__19369\
        );

    \I__4482\ : Span4Mux_v
    port map (
            O => \N__19382\,
            I => \N__19362\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__19379\,
            I => \N__19362\
        );

    \I__4480\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19359\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__19375\,
            I => \N__19356\
        );

    \I__4478\ : InMux
    port map (
            O => \N__19374\,
            I => \N__19353\
        );

    \I__4477\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19350\
        );

    \I__4476\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19347\
        );

    \I__4475\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19344\
        );

    \I__4474\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19341\
        );

    \I__4473\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19338\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__19362\,
            I => \N__19333\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__19359\,
            I => \N__19333\
        );

    \I__4470\ : Sp12to4
    port map (
            O => \N__19356\,
            I => \N__19330\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__19353\,
            I => \N__19327\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__19350\,
            I => \N__19322\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__19347\,
            I => \N__19322\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__19344\,
            I => \N__19319\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__19341\,
            I => \N__19314\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__19338\,
            I => \N__19314\
        );

    \I__4463\ : Span4Mux_v
    port map (
            O => \N__19333\,
            I => \N__19311\
        );

    \I__4462\ : Span12Mux_v
    port map (
            O => \N__19330\,
            I => \N__19306\
        );

    \I__4461\ : Span12Mux_v
    port map (
            O => \N__19327\,
            I => \N__19306\
        );

    \I__4460\ : Span4Mux_h
    port map (
            O => \N__19322\,
            I => \N__19303\
        );

    \I__4459\ : Span4Mux_h
    port map (
            O => \N__19319\,
            I => \N__19298\
        );

    \I__4458\ : Span4Mux_h
    port map (
            O => \N__19314\,
            I => \N__19298\
        );

    \I__4457\ : Odrv4
    port map (
            O => \N__19311\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4456\ : Odrv12
    port map (
            O => \N__19306\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__19303\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__19298\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__4452\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19282\
        );

    \I__4451\ : CascadeMux
    port map (
            O => \N__19285\,
            I => \N__19279\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__19282\,
            I => \N__19275\
        );

    \I__4449\ : InMux
    port map (
            O => \N__19279\,
            I => \N__19272\
        );

    \I__4448\ : CascadeMux
    port map (
            O => \N__19278\,
            I => \N__19269\
        );

    \I__4447\ : Span4Mux_h
    port map (
            O => \N__19275\,
            I => \N__19265\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__19272\,
            I => \N__19262\
        );

    \I__4445\ : InMux
    port map (
            O => \N__19269\,
            I => \N__19259\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__19268\,
            I => \N__19256\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__19265\,
            I => \N__19253\
        );

    \I__4442\ : Span4Mux_h
    port map (
            O => \N__19262\,
            I => \N__19248\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__19259\,
            I => \N__19248\
        );

    \I__4440\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19245\
        );

    \I__4439\ : Span4Mux_v
    port map (
            O => \N__19253\,
            I => \N__19242\
        );

    \I__4438\ : Span4Mux_v
    port map (
            O => \N__19248\,
            I => \N__19239\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__19245\,
            I => \N__19236\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__19242\,
            I => this_sprites_ram_mem_radreg_11
        );

    \I__4435\ : Odrv4
    port map (
            O => \N__19239\,
            I => this_sprites_ram_mem_radreg_11
        );

    \I__4434\ : Odrv12
    port map (
            O => \N__19236\,
            I => this_sprites_ram_mem_radreg_11
        );

    \I__4433\ : InMux
    port map (
            O => \N__19229\,
            I => \N__19226\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__4431\ : Span12Mux_h
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__4430\ : Odrv12
    port map (
            O => \N__19220\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__4429\ : InMux
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__19214\,
            I => \N__19211\
        );

    \I__4427\ : Span4Mux_h
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__4426\ : Odrv4
    port map (
            O => \N__19208\,
            I => \this_sprites_ram.mem_out_bus4_3\
        );

    \I__4425\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__4423\ : Span12Mux_h
    port map (
            O => \N__19199\,
            I => \N__19196\
        );

    \I__4422\ : Span12Mux_v
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__4421\ : Odrv12
    port map (
            O => \N__19193\,
            I => \this_sprites_ram.mem_out_bus0_3\
        );

    \I__4420\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__19187\,
            I => \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_3\
        );

    \I__4418\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19179\
        );

    \I__4417\ : InMux
    port map (
            O => \N__19183\,
            I => \N__19174\
        );

    \I__4416\ : InMux
    port map (
            O => \N__19182\,
            I => \N__19174\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__19179\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__19174\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4413\ : InMux
    port map (
            O => \N__19169\,
            I => \N__19166\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__19166\,
            I => \N__19162\
        );

    \I__4411\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19159\
        );

    \I__4410\ : Span4Mux_h
    port map (
            O => \N__19162\,
            I => \N__19156\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__19159\,
            I => \N_170_0\
        );

    \I__4408\ : Odrv4
    port map (
            O => \N__19156\,
            I => \N_170_0\
        );

    \I__4407\ : CEMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__19148\,
            I => \N__19144\
        );

    \I__4405\ : CEMux
    port map (
            O => \N__19147\,
            I => \N__19141\
        );

    \I__4404\ : Span4Mux_h
    port map (
            O => \N__19144\,
            I => \N__19136\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19141\,
            I => \N__19136\
        );

    \I__4402\ : Span4Mux_v
    port map (
            O => \N__19136\,
            I => \N__19133\
        );

    \I__4401\ : Span4Mux_v
    port map (
            O => \N__19133\,
            I => \N__19130\
        );

    \I__4400\ : Odrv4
    port map (
            O => \N__19130\,
            I => \this_sprites_ram.mem_WE_0\
        );

    \I__4399\ : InMux
    port map (
            O => \N__19127\,
            I => \N__19121\
        );

    \I__4398\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19118\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19125\,
            I => \N__19115\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19124\,
            I => \N__19112\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__19121\,
            I => \N__19105\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__19118\,
            I => \N__19105\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__19115\,
            I => \N__19105\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__19112\,
            I => \this_ppu.M_vaddress_qZ0Z_3\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__19105\,
            I => \this_ppu.M_vaddress_qZ0Z_3\
        );

    \I__4390\ : CascadeMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__4389\ : CascadeBuf
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__4388\ : CascadeMux
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__4387\ : CascadeBuf
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__19088\,
            I => \N__19085\
        );

    \I__4385\ : CascadeBuf
    port map (
            O => \N__19085\,
            I => \N__19082\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__4383\ : CascadeBuf
    port map (
            O => \N__19079\,
            I => \N__19076\
        );

    \I__4382\ : CascadeMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__4381\ : CascadeBuf
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__4379\ : CascadeBuf
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__4377\ : CascadeBuf
    port map (
            O => \N__19061\,
            I => \N__19058\
        );

    \I__4376\ : CascadeMux
    port map (
            O => \N__19058\,
            I => \N__19055\
        );

    \I__4375\ : CascadeBuf
    port map (
            O => \N__19055\,
            I => \N__19052\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__19052\,
            I => \N__19049\
        );

    \I__4373\ : CascadeBuf
    port map (
            O => \N__19049\,
            I => \N__19046\
        );

    \I__4372\ : CascadeMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__4371\ : CascadeBuf
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__4370\ : CascadeMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__4369\ : CascadeBuf
    port map (
            O => \N__19037\,
            I => \N__19034\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__19034\,
            I => \N__19031\
        );

    \I__4367\ : CascadeBuf
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__4366\ : CascadeMux
    port map (
            O => \N__19028\,
            I => \N__19025\
        );

    \I__4365\ : CascadeBuf
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__4363\ : CascadeBuf
    port map (
            O => \N__19019\,
            I => \N__19016\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__19016\,
            I => \N__19013\
        );

    \I__4361\ : CascadeBuf
    port map (
            O => \N__19013\,
            I => \N__19010\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__19010\,
            I => \N__19007\
        );

    \I__4359\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19004\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__4357\ : Span12Mux_s11_h
    port map (
            O => \N__19001\,
            I => \N__18998\
        );

    \I__4356\ : Span12Mux_v
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__4355\ : Odrv12
    port map (
            O => \N__18995\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__4354\ : InMux
    port map (
            O => \N__18992\,
            I => \this_ppu.sprites_addr_cry_9\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__18989\,
            I => \N__18985\
        );

    \I__4352\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18982\
        );

    \I__4351\ : InMux
    port map (
            O => \N__18985\,
            I => \N__18978\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__18982\,
            I => \N__18975\
        );

    \I__4349\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18972\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__18978\,
            I => \this_ppu.M_vaddress_qZ1Z_4\
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__18975\,
            I => \this_ppu.M_vaddress_qZ1Z_4\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__18972\,
            I => \this_ppu.M_vaddress_qZ1Z_4\
        );

    \I__4345\ : InMux
    port map (
            O => \N__18965\,
            I => \this_ppu.sprites_addr_cry_10\
        );

    \I__4344\ : InMux
    port map (
            O => \N__18962\,
            I => \N__18955\
        );

    \I__4343\ : InMux
    port map (
            O => \N__18961\,
            I => \N__18955\
        );

    \I__4342\ : InMux
    port map (
            O => \N__18960\,
            I => \N__18952\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__18955\,
            I => \N__18947\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__18952\,
            I => \N__18947\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__18947\,
            I => \this_ppu.M_vaddress_qZ0Z_5\
        );

    \I__4338\ : InMux
    port map (
            O => \N__18944\,
            I => \this_ppu.sprites_addr_cry_11\
        );

    \I__4337\ : CascadeMux
    port map (
            O => \N__18941\,
            I => \N__18938\
        );

    \I__4336\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18934\
        );

    \I__4335\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18931\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__18934\,
            I => \N__18926\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__18931\,
            I => \N__18926\
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__18926\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__4331\ : InMux
    port map (
            O => \N__18923\,
            I => \this_ppu.sprites_addr_cry_12\
        );

    \I__4330\ : CascadeMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__4329\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__18911\,
            I => \N__18907\
        );

    \I__4326\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18904\
        );

    \I__4325\ : Sp12to4
    port map (
            O => \N__18907\,
            I => \N__18897\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__18904\,
            I => \N__18891\
        );

    \I__4323\ : InMux
    port map (
            O => \N__18903\,
            I => \N__18888\
        );

    \I__4322\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18885\
        );

    \I__4321\ : InMux
    port map (
            O => \N__18901\,
            I => \N__18880\
        );

    \I__4320\ : InMux
    port map (
            O => \N__18900\,
            I => \N__18880\
        );

    \I__4319\ : Span12Mux_v
    port map (
            O => \N__18897\,
            I => \N__18877\
        );

    \I__4318\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18872\
        );

    \I__4317\ : InMux
    port map (
            O => \N__18895\,
            I => \N__18872\
        );

    \I__4316\ : InMux
    port map (
            O => \N__18894\,
            I => \N__18869\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__18891\,
            I => \N__18862\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__18888\,
            I => \N__18862\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__18885\,
            I => \N__18862\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__18880\,
            I => \N__18859\
        );

    \I__4311\ : Odrv12
    port map (
            O => \N__18877\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__18872\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__18869\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__4308\ : Odrv4
    port map (
            O => \N__18862\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__4307\ : Odrv4
    port map (
            O => \N__18859\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__18848\,
            I => \N__18845\
        );

    \I__4305\ : CascadeBuf
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__18842\,
            I => \N__18839\
        );

    \I__4303\ : CascadeBuf
    port map (
            O => \N__18839\,
            I => \N__18836\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__4301\ : CascadeBuf
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__4299\ : CascadeBuf
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__4297\ : CascadeBuf
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__4296\ : CascadeMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__4295\ : CascadeBuf
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__4293\ : CascadeBuf
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__4291\ : CascadeBuf
    port map (
            O => \N__18803\,
            I => \N__18800\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__4289\ : CascadeBuf
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__4287\ : CascadeBuf
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__4285\ : CascadeBuf
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__4284\ : CascadeMux
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__4283\ : CascadeBuf
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__4281\ : CascadeBuf
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__18770\,
            I => \N__18767\
        );

    \I__4279\ : CascadeBuf
    port map (
            O => \N__18767\,
            I => \N__18764\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__4277\ : CascadeBuf
    port map (
            O => \N__18761\,
            I => \N__18758\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__4275\ : InMux
    port map (
            O => \N__18755\,
            I => \N__18752\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__4273\ : Span12Mux_v
    port map (
            O => \N__18749\,
            I => \N__18746\
        );

    \I__4272\ : Odrv12
    port map (
            O => \N__18746\,
            I => \M_this_ppu_vram_addr_i_0\
        );

    \I__4271\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18740\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__4269\ : Span12Mux_h
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__4268\ : Odrv12
    port map (
            O => \N__18734\,
            I => \this_sprites_ram.mem_out_bus5_1\
        );

    \I__4267\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18728\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__18728\,
            I => \N__18725\
        );

    \I__4265\ : Span4Mux_v
    port map (
            O => \N__18725\,
            I => \N__18722\
        );

    \I__4264\ : Span4Mux_v
    port map (
            O => \N__18722\,
            I => \N__18719\
        );

    \I__4263\ : Odrv4
    port map (
            O => \N__18719\,
            I => \this_sprites_ram.mem_out_bus1_1\
        );

    \I__4262\ : InMux
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__18713\,
            I => \N__18710\
        );

    \I__4260\ : Span4Mux_h
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__4259\ : Span4Mux_v
    port map (
            O => \N__18707\,
            I => \N__18704\
        );

    \I__4258\ : Span4Mux_v
    port map (
            O => \N__18704\,
            I => \N__18701\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__18701\,
            I => \N__18698\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__18698\,
            I => \this_sprites_ram.mem_out_bus7_1\
        );

    \I__4255\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__18689\,
            I => \this_sprites_ram.mem_out_bus3_1\
        );

    \I__4252\ : CascadeMux
    port map (
            O => \N__18686\,
            I => \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_1_cascade_\
        );

    \I__4251\ : InMux
    port map (
            O => \N__18683\,
            I => \N__18680\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__18680\,
            I => \this_sprites_ram_mem_N_88\
        );

    \I__4249\ : CEMux
    port map (
            O => \N__18677\,
            I => \N__18674\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__4247\ : Span4Mux_s3_v
    port map (
            O => \N__18671\,
            I => \N__18667\
        );

    \I__4246\ : CEMux
    port map (
            O => \N__18670\,
            I => \N__18664\
        );

    \I__4245\ : Span4Mux_h
    port map (
            O => \N__18667\,
            I => \N__18659\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__18664\,
            I => \N__18659\
        );

    \I__4243\ : Span4Mux_h
    port map (
            O => \N__18659\,
            I => \N__18656\
        );

    \I__4242\ : Span4Mux_v
    port map (
            O => \N__18656\,
            I => \N__18653\
        );

    \I__4241\ : Span4Mux_v
    port map (
            O => \N__18653\,
            I => \N__18650\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__18650\,
            I => \this_sprites_ram.mem_WE_14\
        );

    \I__4239\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18644\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__18644\,
            I => \N__18641\
        );

    \I__4237\ : Span4Mux_v
    port map (
            O => \N__18641\,
            I => \N__18638\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__18638\,
            I => \this_sprites_ram.mem_out_bus2_3\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__18635\,
            I => \N__18632\
        );

    \I__4234\ : InMux
    port map (
            O => \N__18632\,
            I => \N__18629\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__18629\,
            I => \N__18626\
        );

    \I__4232\ : Span12Mux_h
    port map (
            O => \N__18626\,
            I => \N__18623\
        );

    \I__4231\ : Span12Mux_v
    port map (
            O => \N__18623\,
            I => \N__18620\
        );

    \I__4230\ : Odrv12
    port map (
            O => \N__18620\,
            I => \this_sprites_ram.mem_out_bus6_3\
        );

    \I__4229\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__18614\,
            I => \N__18611\
        );

    \I__4227\ : Span4Mux_h
    port map (
            O => \N__18611\,
            I => \N__18608\
        );

    \I__4226\ : Odrv4
    port map (
            O => \N__18608\,
            I => \this_sprites_ram_mem_N_105\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18605\,
            I => \this_ppu.sprites_addr_cry_1\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__18602\,
            I => \N__18599\
        );

    \I__4223\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__18596\,
            I => \N__18592\
        );

    \I__4221\ : InMux
    port map (
            O => \N__18595\,
            I => \N__18587\
        );

    \I__4220\ : Span12Mux_v
    port map (
            O => \N__18592\,
            I => \N__18582\
        );

    \I__4219\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18579\
        );

    \I__4218\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18576\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__18587\,
            I => \N__18573\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18586\,
            I => \N__18568\
        );

    \I__4215\ : InMux
    port map (
            O => \N__18585\,
            I => \N__18568\
        );

    \I__4214\ : Odrv12
    port map (
            O => \N__18582\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__18579\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__18576\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__4211\ : Odrv12
    port map (
            O => \N__18573\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__18568\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__4208\ : CascadeBuf
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__4206\ : CascadeBuf
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__4204\ : CascadeBuf
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__4202\ : CascadeBuf
    port map (
            O => \N__18536\,
            I => \N__18533\
        );

    \I__4201\ : CascadeMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__4200\ : CascadeBuf
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__4198\ : CascadeBuf
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__4196\ : CascadeBuf
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__4194\ : CascadeBuf
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__4192\ : CascadeBuf
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__4190\ : CascadeBuf
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__4189\ : CascadeMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__4188\ : CascadeBuf
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__18491\,
            I => \N__18488\
        );

    \I__4186\ : CascadeBuf
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__4185\ : CascadeMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__4184\ : CascadeBuf
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__4182\ : CascadeBuf
    port map (
            O => \N__18476\,
            I => \N__18473\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__4180\ : CascadeBuf
    port map (
            O => \N__18470\,
            I => \N__18467\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__4178\ : InMux
    port map (
            O => \N__18464\,
            I => \N__18461\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__18458\,
            I => \N__18455\
        );

    \I__4175\ : Span4Mux_h
    port map (
            O => \N__18455\,
            I => \N__18452\
        );

    \I__4174\ : Sp12to4
    port map (
            O => \N__18452\,
            I => \N__18449\
        );

    \I__4173\ : Odrv12
    port map (
            O => \N__18449\,
            I => \M_this_ppu_sprites_addr_3\
        );

    \I__4172\ : InMux
    port map (
            O => \N__18446\,
            I => \this_ppu.sprites_addr_cry_2\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__4170\ : InMux
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__4168\ : Sp12to4
    port map (
            O => \N__18434\,
            I => \N__18427\
        );

    \I__4167\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18424\
        );

    \I__4166\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18421\
        );

    \I__4165\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18418\
        );

    \I__4164\ : CascadeMux
    port map (
            O => \N__18430\,
            I => \N__18415\
        );

    \I__4163\ : Span12Mux_h
    port map (
            O => \N__18427\,
            I => \N__18412\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__18424\,
            I => \N__18405\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__18421\,
            I => \N__18405\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__18418\,
            I => \N__18405\
        );

    \I__4159\ : InMux
    port map (
            O => \N__18415\,
            I => \N__18402\
        );

    \I__4158\ : Odrv12
    port map (
            O => \N__18412\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__4157\ : Odrv12
    port map (
            O => \N__18405\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__18402\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__4155\ : CascadeMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__4154\ : CascadeBuf
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__4152\ : CascadeBuf
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__4151\ : CascadeMux
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__4150\ : CascadeBuf
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__4148\ : CascadeBuf
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__18371\,
            I => \N__18368\
        );

    \I__4146\ : CascadeBuf
    port map (
            O => \N__18368\,
            I => \N__18365\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__18365\,
            I => \N__18362\
        );

    \I__4144\ : CascadeBuf
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__18359\,
            I => \N__18356\
        );

    \I__4142\ : CascadeBuf
    port map (
            O => \N__18356\,
            I => \N__18353\
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__18353\,
            I => \N__18350\
        );

    \I__4140\ : CascadeBuf
    port map (
            O => \N__18350\,
            I => \N__18347\
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__18347\,
            I => \N__18344\
        );

    \I__4138\ : CascadeBuf
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__18341\,
            I => \N__18338\
        );

    \I__4136\ : CascadeBuf
    port map (
            O => \N__18338\,
            I => \N__18335\
        );

    \I__4135\ : CascadeMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__4134\ : CascadeBuf
    port map (
            O => \N__18332\,
            I => \N__18329\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__4132\ : CascadeBuf
    port map (
            O => \N__18326\,
            I => \N__18323\
        );

    \I__4131\ : CascadeMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__4130\ : CascadeBuf
    port map (
            O => \N__18320\,
            I => \N__18317\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__18317\,
            I => \N__18314\
        );

    \I__4128\ : CascadeBuf
    port map (
            O => \N__18314\,
            I => \N__18311\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__18311\,
            I => \N__18308\
        );

    \I__4126\ : CascadeBuf
    port map (
            O => \N__18308\,
            I => \N__18305\
        );

    \I__4125\ : CascadeMux
    port map (
            O => \N__18305\,
            I => \N__18302\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18299\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__4122\ : Span4Mux_s3_v
    port map (
            O => \N__18296\,
            I => \N__18293\
        );

    \I__4121\ : Span4Mux_h
    port map (
            O => \N__18293\,
            I => \N__18290\
        );

    \I__4120\ : Sp12to4
    port map (
            O => \N__18290\,
            I => \N__18287\
        );

    \I__4119\ : Odrv12
    port map (
            O => \N__18287\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__4118\ : InMux
    port map (
            O => \N__18284\,
            I => \this_ppu.sprites_addr_cry_3\
        );

    \I__4117\ : CascadeMux
    port map (
            O => \N__18281\,
            I => \N__18278\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18275\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__18275\,
            I => \N__18271\
        );

    \I__4114\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18266\
        );

    \I__4113\ : Span12Mux_h
    port map (
            O => \N__18271\,
            I => \N__18262\
        );

    \I__4112\ : InMux
    port map (
            O => \N__18270\,
            I => \N__18257\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18269\,
            I => \N__18257\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__18266\,
            I => \N__18254\
        );

    \I__4109\ : InMux
    port map (
            O => \N__18265\,
            I => \N__18251\
        );

    \I__4108\ : Odrv12
    port map (
            O => \N__18262\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__18257\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__18254\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18251\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__18242\,
            I => \N__18239\
        );

    \I__4103\ : CascadeBuf
    port map (
            O => \N__18239\,
            I => \N__18236\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__4101\ : CascadeBuf
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__18230\,
            I => \N__18227\
        );

    \I__4099\ : CascadeBuf
    port map (
            O => \N__18227\,
            I => \N__18224\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__18224\,
            I => \N__18221\
        );

    \I__4097\ : CascadeBuf
    port map (
            O => \N__18221\,
            I => \N__18218\
        );

    \I__4096\ : CascadeMux
    port map (
            O => \N__18218\,
            I => \N__18215\
        );

    \I__4095\ : CascadeBuf
    port map (
            O => \N__18215\,
            I => \N__18212\
        );

    \I__4094\ : CascadeMux
    port map (
            O => \N__18212\,
            I => \N__18209\
        );

    \I__4093\ : CascadeBuf
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__4092\ : CascadeMux
    port map (
            O => \N__18206\,
            I => \N__18203\
        );

    \I__4091\ : CascadeBuf
    port map (
            O => \N__18203\,
            I => \N__18200\
        );

    \I__4090\ : CascadeMux
    port map (
            O => \N__18200\,
            I => \N__18197\
        );

    \I__4089\ : CascadeBuf
    port map (
            O => \N__18197\,
            I => \N__18194\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__18194\,
            I => \N__18191\
        );

    \I__4087\ : CascadeBuf
    port map (
            O => \N__18191\,
            I => \N__18188\
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__4085\ : CascadeBuf
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__4083\ : CascadeBuf
    port map (
            O => \N__18179\,
            I => \N__18176\
        );

    \I__4082\ : CascadeMux
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__4081\ : CascadeBuf
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__18170\,
            I => \N__18167\
        );

    \I__4079\ : CascadeBuf
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__4078\ : CascadeMux
    port map (
            O => \N__18164\,
            I => \N__18161\
        );

    \I__4077\ : CascadeBuf
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__18158\,
            I => \N__18155\
        );

    \I__4075\ : CascadeBuf
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__4073\ : InMux
    port map (
            O => \N__18149\,
            I => \N__18146\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__18146\,
            I => \N__18143\
        );

    \I__4071\ : Sp12to4
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__4070\ : Span12Mux_s3_v
    port map (
            O => \N__18140\,
            I => \N__18137\
        );

    \I__4069\ : Span12Mux_v
    port map (
            O => \N__18137\,
            I => \N__18134\
        );

    \I__4068\ : Odrv12
    port map (
            O => \N__18134\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__4067\ : InMux
    port map (
            O => \N__18131\,
            I => \this_ppu.sprites_addr_cry_4\
        );

    \I__4066\ : CascadeMux
    port map (
            O => \N__18128\,
            I => \N__18125\
        );

    \I__4065\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__18122\,
            I => \N__18119\
        );

    \I__4063\ : Span4Mux_h
    port map (
            O => \N__18119\,
            I => \N__18116\
        );

    \I__4062\ : Sp12to4
    port map (
            O => \N__18116\,
            I => \N__18110\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__18115\,
            I => \N__18107\
        );

    \I__4060\ : InMux
    port map (
            O => \N__18114\,
            I => \N__18104\
        );

    \I__4059\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18101\
        );

    \I__4058\ : Span12Mux_v
    port map (
            O => \N__18110\,
            I => \N__18098\
        );

    \I__4057\ : InMux
    port map (
            O => \N__18107\,
            I => \N__18095\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__18104\,
            I => \N__18090\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__18101\,
            I => \N__18090\
        );

    \I__4054\ : Odrv12
    port map (
            O => \N__18098\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__18095\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__18090\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__4051\ : CascadeMux
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__4050\ : CascadeBuf
    port map (
            O => \N__18080\,
            I => \N__18077\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__18077\,
            I => \N__18074\
        );

    \I__4048\ : CascadeBuf
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__4047\ : CascadeMux
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__4046\ : CascadeBuf
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__4044\ : CascadeBuf
    port map (
            O => \N__18062\,
            I => \N__18059\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__18059\,
            I => \N__18056\
        );

    \I__4042\ : CascadeBuf
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__18053\,
            I => \N__18050\
        );

    \I__4040\ : CascadeBuf
    port map (
            O => \N__18050\,
            I => \N__18047\
        );

    \I__4039\ : CascadeMux
    port map (
            O => \N__18047\,
            I => \N__18044\
        );

    \I__4038\ : CascadeBuf
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__4036\ : CascadeBuf
    port map (
            O => \N__18038\,
            I => \N__18035\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__18035\,
            I => \N__18032\
        );

    \I__4034\ : CascadeBuf
    port map (
            O => \N__18032\,
            I => \N__18029\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__18029\,
            I => \N__18026\
        );

    \I__4032\ : CascadeBuf
    port map (
            O => \N__18026\,
            I => \N__18023\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__18023\,
            I => \N__18020\
        );

    \I__4030\ : CascadeBuf
    port map (
            O => \N__18020\,
            I => \N__18017\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__18017\,
            I => \N__18014\
        );

    \I__4028\ : CascadeBuf
    port map (
            O => \N__18014\,
            I => \N__18011\
        );

    \I__4027\ : CascadeMux
    port map (
            O => \N__18011\,
            I => \N__18008\
        );

    \I__4026\ : CascadeBuf
    port map (
            O => \N__18008\,
            I => \N__18005\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__18005\,
            I => \N__18002\
        );

    \I__4024\ : CascadeBuf
    port map (
            O => \N__18002\,
            I => \N__17999\
        );

    \I__4023\ : CascadeMux
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__4022\ : CascadeBuf
    port map (
            O => \N__17996\,
            I => \N__17993\
        );

    \I__4021\ : CascadeMux
    port map (
            O => \N__17993\,
            I => \N__17990\
        );

    \I__4020\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__17987\,
            I => \N__17984\
        );

    \I__4018\ : Span4Mux_v
    port map (
            O => \N__17984\,
            I => \N__17981\
        );

    \I__4017\ : Span4Mux_h
    port map (
            O => \N__17981\,
            I => \N__17978\
        );

    \I__4016\ : Span4Mux_v
    port map (
            O => \N__17978\,
            I => \N__17975\
        );

    \I__4015\ : Span4Mux_v
    port map (
            O => \N__17975\,
            I => \N__17972\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__17972\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__4013\ : InMux
    port map (
            O => \N__17969\,
            I => \this_ppu.sprites_addr_cry_5\
        );

    \I__4012\ : CascadeMux
    port map (
            O => \N__17966\,
            I => \N__17963\
        );

    \I__4011\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17960\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__17960\,
            I => \N__17956\
        );

    \I__4009\ : InMux
    port map (
            O => \N__17959\,
            I => \N__17953\
        );

    \I__4008\ : Span4Mux_h
    port map (
            O => \N__17956\,
            I => \N__17950\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__17953\,
            I => \N__17947\
        );

    \I__4006\ : Span4Mux_v
    port map (
            O => \N__17950\,
            I => \N__17944\
        );

    \I__4005\ : Span4Mux_h
    port map (
            O => \N__17947\,
            I => \N__17940\
        );

    \I__4004\ : Span4Mux_h
    port map (
            O => \N__17944\,
            I => \N__17936\
        );

    \I__4003\ : InMux
    port map (
            O => \N__17943\,
            I => \N__17933\
        );

    \I__4002\ : Span4Mux_h
    port map (
            O => \N__17940\,
            I => \N__17930\
        );

    \I__4001\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17927\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__17936\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__17933\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__3998\ : Odrv4
    port map (
            O => \N__17930\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__17927\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__3996\ : CascadeMux
    port map (
            O => \N__17918\,
            I => \N__17915\
        );

    \I__3995\ : CascadeBuf
    port map (
            O => \N__17915\,
            I => \N__17912\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__17912\,
            I => \N__17909\
        );

    \I__3993\ : CascadeBuf
    port map (
            O => \N__17909\,
            I => \N__17906\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__17906\,
            I => \N__17903\
        );

    \I__3991\ : CascadeBuf
    port map (
            O => \N__17903\,
            I => \N__17900\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__3989\ : CascadeBuf
    port map (
            O => \N__17897\,
            I => \N__17894\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__17894\,
            I => \N__17891\
        );

    \I__3987\ : CascadeBuf
    port map (
            O => \N__17891\,
            I => \N__17888\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__17888\,
            I => \N__17885\
        );

    \I__3985\ : CascadeBuf
    port map (
            O => \N__17885\,
            I => \N__17882\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__17882\,
            I => \N__17879\
        );

    \I__3983\ : CascadeBuf
    port map (
            O => \N__17879\,
            I => \N__17876\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__17876\,
            I => \N__17873\
        );

    \I__3981\ : CascadeBuf
    port map (
            O => \N__17873\,
            I => \N__17870\
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__17870\,
            I => \N__17867\
        );

    \I__3979\ : CascadeBuf
    port map (
            O => \N__17867\,
            I => \N__17864\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__17864\,
            I => \N__17861\
        );

    \I__3977\ : CascadeBuf
    port map (
            O => \N__17861\,
            I => \N__17858\
        );

    \I__3976\ : CascadeMux
    port map (
            O => \N__17858\,
            I => \N__17855\
        );

    \I__3975\ : CascadeBuf
    port map (
            O => \N__17855\,
            I => \N__17852\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__17852\,
            I => \N__17849\
        );

    \I__3973\ : CascadeBuf
    port map (
            O => \N__17849\,
            I => \N__17846\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__3971\ : CascadeBuf
    port map (
            O => \N__17843\,
            I => \N__17840\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__17840\,
            I => \N__17837\
        );

    \I__3969\ : CascadeBuf
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__3968\ : CascadeMux
    port map (
            O => \N__17834\,
            I => \N__17831\
        );

    \I__3967\ : CascadeBuf
    port map (
            O => \N__17831\,
            I => \N__17828\
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__17828\,
            I => \N__17825\
        );

    \I__3965\ : InMux
    port map (
            O => \N__17825\,
            I => \N__17822\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__17822\,
            I => \N__17819\
        );

    \I__3963\ : Span4Mux_v
    port map (
            O => \N__17819\,
            I => \N__17816\
        );

    \I__3962\ : Span4Mux_h
    port map (
            O => \N__17816\,
            I => \N__17813\
        );

    \I__3961\ : Span4Mux_v
    port map (
            O => \N__17813\,
            I => \N__17810\
        );

    \I__3960\ : Span4Mux_v
    port map (
            O => \N__17810\,
            I => \N__17807\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__17807\,
            I => \M_this_ppu_sprites_addr_7\
        );

    \I__3958\ : InMux
    port map (
            O => \N__17804\,
            I => \this_ppu.sprites_addr_cry_6\
        );

    \I__3957\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17798\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__17798\,
            I => \N__17793\
        );

    \I__3955\ : InMux
    port map (
            O => \N__17797\,
            I => \N__17789\
        );

    \I__3954\ : InMux
    port map (
            O => \N__17796\,
            I => \N__17786\
        );

    \I__3953\ : Span4Mux_v
    port map (
            O => \N__17793\,
            I => \N__17783\
        );

    \I__3952\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17780\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__17789\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__17786\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__17783\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__17780\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__17771\,
            I => \N__17768\
        );

    \I__3946\ : CascadeBuf
    port map (
            O => \N__17768\,
            I => \N__17765\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__17765\,
            I => \N__17762\
        );

    \I__3944\ : CascadeBuf
    port map (
            O => \N__17762\,
            I => \N__17759\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__17759\,
            I => \N__17756\
        );

    \I__3942\ : CascadeBuf
    port map (
            O => \N__17756\,
            I => \N__17753\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__17753\,
            I => \N__17750\
        );

    \I__3940\ : CascadeBuf
    port map (
            O => \N__17750\,
            I => \N__17747\
        );

    \I__3939\ : CascadeMux
    port map (
            O => \N__17747\,
            I => \N__17744\
        );

    \I__3938\ : CascadeBuf
    port map (
            O => \N__17744\,
            I => \N__17741\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__17741\,
            I => \N__17738\
        );

    \I__3936\ : CascadeBuf
    port map (
            O => \N__17738\,
            I => \N__17735\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__17735\,
            I => \N__17732\
        );

    \I__3934\ : CascadeBuf
    port map (
            O => \N__17732\,
            I => \N__17729\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__17729\,
            I => \N__17726\
        );

    \I__3932\ : CascadeBuf
    port map (
            O => \N__17726\,
            I => \N__17723\
        );

    \I__3931\ : CascadeMux
    port map (
            O => \N__17723\,
            I => \N__17720\
        );

    \I__3930\ : CascadeBuf
    port map (
            O => \N__17720\,
            I => \N__17717\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__3928\ : CascadeBuf
    port map (
            O => \N__17714\,
            I => \N__17711\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__17711\,
            I => \N__17708\
        );

    \I__3926\ : CascadeBuf
    port map (
            O => \N__17708\,
            I => \N__17705\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__17705\,
            I => \N__17702\
        );

    \I__3924\ : CascadeBuf
    port map (
            O => \N__17702\,
            I => \N__17699\
        );

    \I__3923\ : CascadeMux
    port map (
            O => \N__17699\,
            I => \N__17696\
        );

    \I__3922\ : CascadeBuf
    port map (
            O => \N__17696\,
            I => \N__17693\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__17693\,
            I => \N__17690\
        );

    \I__3920\ : CascadeBuf
    port map (
            O => \N__17690\,
            I => \N__17687\
        );

    \I__3919\ : CascadeMux
    port map (
            O => \N__17687\,
            I => \N__17684\
        );

    \I__3918\ : CascadeBuf
    port map (
            O => \N__17684\,
            I => \N__17681\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__17681\,
            I => \N__17678\
        );

    \I__3916\ : InMux
    port map (
            O => \N__17678\,
            I => \N__17675\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__17675\,
            I => \N__17672\
        );

    \I__3914\ : Span4Mux_v
    port map (
            O => \N__17672\,
            I => \N__17669\
        );

    \I__3913\ : Span4Mux_h
    port map (
            O => \N__17669\,
            I => \N__17666\
        );

    \I__3912\ : Span4Mux_v
    port map (
            O => \N__17666\,
            I => \N__17663\
        );

    \I__3911\ : Span4Mux_v
    port map (
            O => \N__17663\,
            I => \N__17660\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__17660\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__3909\ : InMux
    port map (
            O => \N__17657\,
            I => \this_ppu.sprites_addr_cry_7\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__17654\,
            I => \N__17650\
        );

    \I__3907\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17647\
        );

    \I__3906\ : InMux
    port map (
            O => \N__17650\,
            I => \N__17643\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__17647\,
            I => \N__17640\
        );

    \I__3904\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17637\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__17643\,
            I => \this_ppu.M_vaddress_qZ1Z_2\
        );

    \I__3902\ : Odrv12
    port map (
            O => \N__17640\,
            I => \this_ppu.M_vaddress_qZ1Z_2\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__17637\,
            I => \this_ppu.M_vaddress_qZ1Z_2\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__17630\,
            I => \N__17627\
        );

    \I__3899\ : CascadeBuf
    port map (
            O => \N__17627\,
            I => \N__17624\
        );

    \I__3898\ : CascadeMux
    port map (
            O => \N__17624\,
            I => \N__17621\
        );

    \I__3897\ : CascadeBuf
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__17618\,
            I => \N__17615\
        );

    \I__3895\ : CascadeBuf
    port map (
            O => \N__17615\,
            I => \N__17612\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__17612\,
            I => \N__17609\
        );

    \I__3893\ : CascadeBuf
    port map (
            O => \N__17609\,
            I => \N__17606\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__17606\,
            I => \N__17603\
        );

    \I__3891\ : CascadeBuf
    port map (
            O => \N__17603\,
            I => \N__17600\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__17600\,
            I => \N__17597\
        );

    \I__3889\ : CascadeBuf
    port map (
            O => \N__17597\,
            I => \N__17594\
        );

    \I__3888\ : CascadeMux
    port map (
            O => \N__17594\,
            I => \N__17591\
        );

    \I__3887\ : CascadeBuf
    port map (
            O => \N__17591\,
            I => \N__17588\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__17588\,
            I => \N__17585\
        );

    \I__3885\ : CascadeBuf
    port map (
            O => \N__17585\,
            I => \N__17582\
        );

    \I__3884\ : CascadeMux
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__3883\ : CascadeBuf
    port map (
            O => \N__17579\,
            I => \N__17576\
        );

    \I__3882\ : CascadeMux
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__3881\ : CascadeBuf
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__3879\ : CascadeBuf
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__3878\ : CascadeMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__3877\ : CascadeBuf
    port map (
            O => \N__17561\,
            I => \N__17558\
        );

    \I__3876\ : CascadeMux
    port map (
            O => \N__17558\,
            I => \N__17555\
        );

    \I__3875\ : CascadeBuf
    port map (
            O => \N__17555\,
            I => \N__17552\
        );

    \I__3874\ : CascadeMux
    port map (
            O => \N__17552\,
            I => \N__17549\
        );

    \I__3873\ : CascadeBuf
    port map (
            O => \N__17549\,
            I => \N__17546\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__3871\ : CascadeBuf
    port map (
            O => \N__17543\,
            I => \N__17540\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__3869\ : InMux
    port map (
            O => \N__17537\,
            I => \N__17534\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__17534\,
            I => \N__17531\
        );

    \I__3867\ : Span4Mux_s2_v
    port map (
            O => \N__17531\,
            I => \N__17528\
        );

    \I__3866\ : Span4Mux_v
    port map (
            O => \N__17528\,
            I => \N__17525\
        );

    \I__3865\ : Span4Mux_v
    port map (
            O => \N__17525\,
            I => \N__17522\
        );

    \I__3864\ : Span4Mux_v
    port map (
            O => \N__17522\,
            I => \N__17519\
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__17519\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__3862\ : InMux
    port map (
            O => \N__17516\,
            I => \bfn_21_18_0_\
        );

    \I__3861\ : InMux
    port map (
            O => \N__17513\,
            I => \N__17499\
        );

    \I__3860\ : InMux
    port map (
            O => \N__17512\,
            I => \N__17499\
        );

    \I__3859\ : InMux
    port map (
            O => \N__17511\,
            I => \N__17496\
        );

    \I__3858\ : InMux
    port map (
            O => \N__17510\,
            I => \N__17491\
        );

    \I__3857\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17484\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17508\,
            I => \N__17484\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17484\
        );

    \I__3854\ : InMux
    port map (
            O => \N__17506\,
            I => \N__17479\
        );

    \I__3853\ : InMux
    port map (
            O => \N__17505\,
            I => \N__17474\
        );

    \I__3852\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17474\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__17499\,
            I => \N__17469\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__17496\,
            I => \N__17469\
        );

    \I__3849\ : InMux
    port map (
            O => \N__17495\,
            I => \N__17464\
        );

    \I__3848\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17464\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__17491\,
            I => \N__17459\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__17484\,
            I => \N__17459\
        );

    \I__3845\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17454\
        );

    \I__3844\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17454\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17479\,
            I => \N__17451\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__17474\,
            I => \N__17448\
        );

    \I__3841\ : Span4Mux_v
    port map (
            O => \N__17469\,
            I => \N__17439\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__17464\,
            I => \N__17439\
        );

    \I__3839\ : Span4Mux_v
    port map (
            O => \N__17459\,
            I => \N__17439\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__17454\,
            I => \N__17439\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__17451\,
            I => \M_this_sprites_address_q_3_sm0_0\
        );

    \I__3836\ : Odrv4
    port map (
            O => \N__17448\,
            I => \M_this_sprites_address_q_3_sm0_0\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__17439\,
            I => \M_this_sprites_address_q_3_sm0_0\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__17432\,
            I => \M_this_sprites_address_q_3_ns_1_3_cascade_\
        );

    \I__3833\ : InMux
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__17426\,
            I => \N__17423\
        );

    \I__3831\ : Span12Mux_s10_v
    port map (
            O => \N__17423\,
            I => \N__17420\
        );

    \I__3830\ : Odrv12
    port map (
            O => \N__17420\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_3\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__17417\,
            I => \N__17414\
        );

    \I__3828\ : CascadeBuf
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__3826\ : CascadeBuf
    port map (
            O => \N__17408\,
            I => \N__17405\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__17405\,
            I => \N__17402\
        );

    \I__3824\ : CascadeBuf
    port map (
            O => \N__17402\,
            I => \N__17399\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3822\ : CascadeBuf
    port map (
            O => \N__17396\,
            I => \N__17393\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__17393\,
            I => \N__17390\
        );

    \I__3820\ : CascadeBuf
    port map (
            O => \N__17390\,
            I => \N__17387\
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__17387\,
            I => \N__17384\
        );

    \I__3818\ : CascadeBuf
    port map (
            O => \N__17384\,
            I => \N__17381\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__17381\,
            I => \N__17378\
        );

    \I__3816\ : CascadeBuf
    port map (
            O => \N__17378\,
            I => \N__17375\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__17375\,
            I => \N__17372\
        );

    \I__3814\ : CascadeBuf
    port map (
            O => \N__17372\,
            I => \N__17369\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__17369\,
            I => \N__17366\
        );

    \I__3812\ : CascadeBuf
    port map (
            O => \N__17366\,
            I => \N__17363\
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__17363\,
            I => \N__17360\
        );

    \I__3810\ : CascadeBuf
    port map (
            O => \N__17360\,
            I => \N__17357\
        );

    \I__3809\ : CascadeMux
    port map (
            O => \N__17357\,
            I => \N__17354\
        );

    \I__3808\ : CascadeBuf
    port map (
            O => \N__17354\,
            I => \N__17351\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__17351\,
            I => \N__17348\
        );

    \I__3806\ : CascadeBuf
    port map (
            O => \N__17348\,
            I => \N__17345\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__17345\,
            I => \N__17342\
        );

    \I__3804\ : CascadeBuf
    port map (
            O => \N__17342\,
            I => \N__17339\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__17339\,
            I => \N__17336\
        );

    \I__3802\ : CascadeBuf
    port map (
            O => \N__17336\,
            I => \N__17333\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__17333\,
            I => \N__17330\
        );

    \I__3800\ : CascadeBuf
    port map (
            O => \N__17330\,
            I => \N__17327\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17324\,
            I => \N__17320\
        );

    \I__3797\ : InMux
    port map (
            O => \N__17323\,
            I => \N__17317\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__17320\,
            I => \N__17314\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__17317\,
            I => \N__17310\
        );

    \I__3794\ : Span4Mux_s2_v
    port map (
            O => \N__17314\,
            I => \N__17307\
        );

    \I__3793\ : CascadeMux
    port map (
            O => \N__17313\,
            I => \N__17304\
        );

    \I__3792\ : Span4Mux_h
    port map (
            O => \N__17310\,
            I => \N__17301\
        );

    \I__3791\ : Span4Mux_h
    port map (
            O => \N__17307\,
            I => \N__17298\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17295\
        );

    \I__3789\ : Span4Mux_h
    port map (
            O => \N__17301\,
            I => \N__17290\
        );

    \I__3788\ : Span4Mux_v
    port map (
            O => \N__17298\,
            I => \N__17290\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__17295\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__17290\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__3785\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17282\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__17282\,
            I => \N__17279\
        );

    \I__3783\ : Span4Mux_v
    port map (
            O => \N__17279\,
            I => \N__17276\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__17276\,
            I => \N__17273\
        );

    \I__3781\ : Sp12to4
    port map (
            O => \N__17273\,
            I => \N__17270\
        );

    \I__3780\ : Odrv12
    port map (
            O => \N__17270\,
            I => \this_sprites_ram.mem_out_bus5_3\
        );

    \I__3779\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__17264\,
            I => \N__17261\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__17261\,
            I => \N__17258\
        );

    \I__3776\ : Odrv4
    port map (
            O => \N__17258\,
            I => \this_sprites_ram.mem_out_bus1_3\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17255\,
            I => \N__17252\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__17252\,
            I => \N__17249\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__17249\,
            I => \N__17246\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__17246\,
            I => \N__17243\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__17243\,
            I => \this_sprites_ram.mem_out_bus3_3\
        );

    \I__3770\ : CascadeMux
    port map (
            O => \N__17240\,
            I => \N__17237\
        );

    \I__3769\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17234\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__17234\,
            I => \N__17231\
        );

    \I__3767\ : Span12Mux_h
    port map (
            O => \N__17231\,
            I => \N__17228\
        );

    \I__3766\ : Span12Mux_v
    port map (
            O => \N__17228\,
            I => \N__17225\
        );

    \I__3765\ : Odrv12
    port map (
            O => \N__17225\,
            I => \this_sprites_ram.mem_out_bus7_3\
        );

    \I__3764\ : InMux
    port map (
            O => \N__17222\,
            I => \N__17219\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__17219\,
            I => \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_3\
        );

    \I__3762\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17213\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__17213\,
            I => \this_sprites_ram_mem_N_102\
        );

    \I__3760\ : InMux
    port map (
            O => \N__17210\,
            I => \N__17207\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__17207\,
            I => \N__17204\
        );

    \I__3758\ : Span4Mux_v
    port map (
            O => \N__17204\,
            I => \N__17201\
        );

    \I__3757\ : Span4Mux_h
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__3756\ : Sp12to4
    port map (
            O => \N__17198\,
            I => \N__17195\
        );

    \I__3755\ : Odrv12
    port map (
            O => \N__17195\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__3754\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__17189\,
            I => \N__17186\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__17186\,
            I => \N__17183\
        );

    \I__3751\ : Span4Mux_h
    port map (
            O => \N__17183\,
            I => \N__17180\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__17180\,
            I => \this_sprites_ram.mem_out_bus2_1\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__17177\,
            I => \N__17174\
        );

    \I__3748\ : InMux
    port map (
            O => \N__17174\,
            I => \N__17171\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__17171\,
            I => \N__17168\
        );

    \I__3746\ : Span4Mux_v
    port map (
            O => \N__17168\,
            I => \N__17165\
        );

    \I__3745\ : Span4Mux_v
    port map (
            O => \N__17165\,
            I => \N__17162\
        );

    \I__3744\ : Span4Mux_h
    port map (
            O => \N__17162\,
            I => \N__17159\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__17159\,
            I => \this_sprites_ram.mem_out_bus6_1\
        );

    \I__3742\ : InMux
    port map (
            O => \N__17156\,
            I => \N__17153\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__17153\,
            I => \this_sprites_ram_mem_N_91\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17150\,
            I => \N__17147\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__17147\,
            I => \N__17144\
        );

    \I__3738\ : Span4Mux_h
    port map (
            O => \N__17144\,
            I => \N__17141\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__17141\,
            I => \this_sprites_ram.mem_out_bus4_1\
        );

    \I__3736\ : InMux
    port map (
            O => \N__17138\,
            I => \N__17135\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__17135\,
            I => \N__17132\
        );

    \I__3734\ : Span4Mux_h
    port map (
            O => \N__17132\,
            I => \N__17129\
        );

    \I__3733\ : Sp12to4
    port map (
            O => \N__17129\,
            I => \N__17126\
        );

    \I__3732\ : Span12Mux_v
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__3731\ : Odrv12
    port map (
            O => \N__17123\,
            I => \this_sprites_ram.mem_out_bus0_1\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17117\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17117\,
            I => \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_1\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__17114\,
            I => \N__17111\
        );

    \I__3727\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17108\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__17108\,
            I => \N__17104\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__17107\,
            I => \N__17101\
        );

    \I__3724\ : Span4Mux_v
    port map (
            O => \N__17104\,
            I => \N__17096\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17093\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17090\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__17099\,
            I => \N__17087\
        );

    \I__3720\ : Sp12to4
    port map (
            O => \N__17096\,
            I => \N__17082\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__17093\,
            I => \N__17076\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__17090\,
            I => \N__17076\
        );

    \I__3717\ : InMux
    port map (
            O => \N__17087\,
            I => \N__17073\
        );

    \I__3716\ : InMux
    port map (
            O => \N__17086\,
            I => \N__17070\
        );

    \I__3715\ : InMux
    port map (
            O => \N__17085\,
            I => \N__17067\
        );

    \I__3714\ : Span12Mux_h
    port map (
            O => \N__17082\,
            I => \N__17064\
        );

    \I__3713\ : InMux
    port map (
            O => \N__17081\,
            I => \N__17061\
        );

    \I__3712\ : Span4Mux_h
    port map (
            O => \N__17076\,
            I => \N__17056\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__17073\,
            I => \N__17056\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__17070\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__17067\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__3708\ : Odrv12
    port map (
            O => \N__17064\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__17061\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__17056\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__3704\ : InMux
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__17039\,
            I => \N__17036\
        );

    \I__3702\ : Span4Mux_v
    port map (
            O => \N__17036\,
            I => \N__17032\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__17035\,
            I => \N__17028\
        );

    \I__3700\ : Sp12to4
    port map (
            O => \N__17032\,
            I => \N__17022\
        );

    \I__3699\ : InMux
    port map (
            O => \N__17031\,
            I => \N__17018\
        );

    \I__3698\ : InMux
    port map (
            O => \N__17028\,
            I => \N__17013\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17013\
        );

    \I__3696\ : InMux
    port map (
            O => \N__17026\,
            I => \N__17010\
        );

    \I__3695\ : InMux
    port map (
            O => \N__17025\,
            I => \N__17007\
        );

    \I__3694\ : Span12Mux_h
    port map (
            O => \N__17022\,
            I => \N__17004\
        );

    \I__3693\ : InMux
    port map (
            O => \N__17021\,
            I => \N__17001\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__17018\,
            I => \N__16998\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__17013\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__17010\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__17007\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__3688\ : Odrv12
    port map (
            O => \N__17004\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__17001\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__16998\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__16985\,
            I => \N__16982\
        );

    \I__3684\ : CascadeBuf
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__16979\,
            I => \N__16976\
        );

    \I__3682\ : CascadeBuf
    port map (
            O => \N__16976\,
            I => \N__16973\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__16973\,
            I => \N__16970\
        );

    \I__3680\ : CascadeBuf
    port map (
            O => \N__16970\,
            I => \N__16967\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__16967\,
            I => \N__16964\
        );

    \I__3678\ : CascadeBuf
    port map (
            O => \N__16964\,
            I => \N__16961\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__16961\,
            I => \N__16958\
        );

    \I__3676\ : CascadeBuf
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__16955\,
            I => \N__16952\
        );

    \I__3674\ : CascadeBuf
    port map (
            O => \N__16952\,
            I => \N__16949\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__16949\,
            I => \N__16946\
        );

    \I__3672\ : CascadeBuf
    port map (
            O => \N__16946\,
            I => \N__16943\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__16943\,
            I => \N__16940\
        );

    \I__3670\ : CascadeBuf
    port map (
            O => \N__16940\,
            I => \N__16937\
        );

    \I__3669\ : CascadeMux
    port map (
            O => \N__16937\,
            I => \N__16934\
        );

    \I__3668\ : CascadeBuf
    port map (
            O => \N__16934\,
            I => \N__16931\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__3666\ : CascadeBuf
    port map (
            O => \N__16928\,
            I => \N__16925\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__16925\,
            I => \N__16922\
        );

    \I__3664\ : CascadeBuf
    port map (
            O => \N__16922\,
            I => \N__16919\
        );

    \I__3663\ : CascadeMux
    port map (
            O => \N__16919\,
            I => \N__16916\
        );

    \I__3662\ : CascadeBuf
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__16913\,
            I => \N__16910\
        );

    \I__3660\ : CascadeBuf
    port map (
            O => \N__16910\,
            I => \N__16907\
        );

    \I__3659\ : CascadeMux
    port map (
            O => \N__16907\,
            I => \N__16904\
        );

    \I__3658\ : CascadeBuf
    port map (
            O => \N__16904\,
            I => \N__16901\
        );

    \I__3657\ : CascadeMux
    port map (
            O => \N__16901\,
            I => \N__16898\
        );

    \I__3656\ : CascadeBuf
    port map (
            O => \N__16898\,
            I => \N__16895\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__16895\,
            I => \N__16892\
        );

    \I__3654\ : InMux
    port map (
            O => \N__16892\,
            I => \N__16889\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__16889\,
            I => \N__16886\
        );

    \I__3652\ : Span4Mux_v
    port map (
            O => \N__16886\,
            I => \N__16883\
        );

    \I__3651\ : Span4Mux_h
    port map (
            O => \N__16883\,
            I => \N__16880\
        );

    \I__3650\ : Sp12to4
    port map (
            O => \N__16880\,
            I => \N__16877\
        );

    \I__3649\ : Odrv12
    port map (
            O => \N__16877\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__3648\ : InMux
    port map (
            O => \N__16874\,
            I => \N__16871\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__16871\,
            I => \this_ppu.un1_M_vaddress_q_c5\
        );

    \I__3646\ : InMux
    port map (
            O => \N__16868\,
            I => \N__16856\
        );

    \I__3645\ : InMux
    port map (
            O => \N__16867\,
            I => \N__16856\
        );

    \I__3644\ : InMux
    port map (
            O => \N__16866\,
            I => \N__16856\
        );

    \I__3643\ : InMux
    port map (
            O => \N__16865\,
            I => \N__16851\
        );

    \I__3642\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16851\
        );

    \I__3641\ : InMux
    port map (
            O => \N__16863\,
            I => \N__16847\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__16856\,
            I => \N__16842\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__16851\,
            I => \N__16842\
        );

    \I__3638\ : InMux
    port map (
            O => \N__16850\,
            I => \N__16839\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__16847\,
            I => \N__16832\
        );

    \I__3636\ : Span4Mux_h
    port map (
            O => \N__16842\,
            I => \N__16832\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__16839\,
            I => \N__16832\
        );

    \I__3634\ : Odrv4
    port map (
            O => \N__16832\,
            I => \this_ppu.N_258_1\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__16829\,
            I => \this_ppu.un1_M_vaddress_q_c5_cascade_\
        );

    \I__3632\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16823\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__16823\,
            I => \N__16820\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__16820\,
            I => \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_13\
        );

    \I__3629\ : CascadeMux
    port map (
            O => \N__16817\,
            I => \N__16814\
        );

    \I__3628\ : CascadeBuf
    port map (
            O => \N__16814\,
            I => \N__16811\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__16811\,
            I => \N__16808\
        );

    \I__3626\ : CascadeBuf
    port map (
            O => \N__16808\,
            I => \N__16805\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__16805\,
            I => \N__16802\
        );

    \I__3624\ : CascadeBuf
    port map (
            O => \N__16802\,
            I => \N__16799\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__16799\,
            I => \N__16796\
        );

    \I__3622\ : CascadeBuf
    port map (
            O => \N__16796\,
            I => \N__16793\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__16793\,
            I => \N__16790\
        );

    \I__3620\ : CascadeBuf
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__16787\,
            I => \N__16784\
        );

    \I__3618\ : CascadeBuf
    port map (
            O => \N__16784\,
            I => \N__16781\
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__16781\,
            I => \N__16778\
        );

    \I__3616\ : CascadeBuf
    port map (
            O => \N__16778\,
            I => \N__16775\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__16775\,
            I => \N__16772\
        );

    \I__3614\ : CascadeBuf
    port map (
            O => \N__16772\,
            I => \N__16769\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__16769\,
            I => \N__16766\
        );

    \I__3612\ : CascadeBuf
    port map (
            O => \N__16766\,
            I => \N__16763\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__3610\ : CascadeBuf
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__16757\,
            I => \N__16754\
        );

    \I__3608\ : CascadeBuf
    port map (
            O => \N__16754\,
            I => \N__16751\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__16751\,
            I => \N__16748\
        );

    \I__3606\ : CascadeBuf
    port map (
            O => \N__16748\,
            I => \N__16745\
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__3604\ : CascadeBuf
    port map (
            O => \N__16742\,
            I => \N__16739\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__16739\,
            I => \N__16736\
        );

    \I__3602\ : CascadeBuf
    port map (
            O => \N__16736\,
            I => \N__16733\
        );

    \I__3601\ : CascadeMux
    port map (
            O => \N__16733\,
            I => \N__16730\
        );

    \I__3600\ : CascadeBuf
    port map (
            O => \N__16730\,
            I => \N__16727\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__16727\,
            I => \N__16723\
        );

    \I__3598\ : InMux
    port map (
            O => \N__16726\,
            I => \N__16720\
        );

    \I__3597\ : InMux
    port map (
            O => \N__16723\,
            I => \N__16717\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__16720\,
            I => \N__16713\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__16717\,
            I => \N__16710\
        );

    \I__3594\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16707\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__16713\,
            I => \N__16704\
        );

    \I__3592\ : Span12Mux_h
    port map (
            O => \N__16710\,
            I => \N__16701\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__16707\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__16704\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__3589\ : Odrv12
    port map (
            O => \N__16701\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__16694\,
            I => \N__16691\
        );

    \I__3587\ : InMux
    port map (
            O => \N__16691\,
            I => \N__16688\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__16688\,
            I => \N__16685\
        );

    \I__3585\ : Span4Mux_v
    port map (
            O => \N__16685\,
            I => \N__16682\
        );

    \I__3584\ : Span4Mux_h
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__16679\,
            I => \M_this_sprites_address_q_3_ns_1_2\
        );

    \I__3582\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__3580\ : Span12Mux_h
    port map (
            O => \N__16670\,
            I => \N__16667\
        );

    \I__3579\ : Odrv12
    port map (
            O => \N__16667\,
            I => \M_this_ppu_vram_data_3\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__3577\ : CascadeBuf
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__3576\ : CascadeMux
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__3575\ : CascadeBuf
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3573\ : CascadeBuf
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__16646\,
            I => \N__16643\
        );

    \I__3571\ : CascadeBuf
    port map (
            O => \N__16643\,
            I => \N__16640\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__16640\,
            I => \N__16637\
        );

    \I__3569\ : CascadeBuf
    port map (
            O => \N__16637\,
            I => \N__16634\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__16634\,
            I => \N__16631\
        );

    \I__3567\ : CascadeBuf
    port map (
            O => \N__16631\,
            I => \N__16628\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__16628\,
            I => \N__16625\
        );

    \I__3565\ : CascadeBuf
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__16622\,
            I => \N__16619\
        );

    \I__3563\ : CascadeBuf
    port map (
            O => \N__16619\,
            I => \N__16616\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__16616\,
            I => \N__16613\
        );

    \I__3561\ : CascadeBuf
    port map (
            O => \N__16613\,
            I => \N__16610\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__16610\,
            I => \N__16607\
        );

    \I__3559\ : CascadeBuf
    port map (
            O => \N__16607\,
            I => \N__16604\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__16604\,
            I => \N__16601\
        );

    \I__3557\ : CascadeBuf
    port map (
            O => \N__16601\,
            I => \N__16598\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__3555\ : CascadeBuf
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__3553\ : CascadeBuf
    port map (
            O => \N__16589\,
            I => \N__16586\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__16586\,
            I => \N__16583\
        );

    \I__3551\ : CascadeBuf
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__3549\ : CascadeBuf
    port map (
            O => \N__16577\,
            I => \N__16574\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__3547\ : InMux
    port map (
            O => \N__16571\,
            I => \N__16568\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__16568\,
            I => \N__16565\
        );

    \I__3545\ : Span12Mux_s3_v
    port map (
            O => \N__16565\,
            I => \N__16562\
        );

    \I__3544\ : Span12Mux_v
    port map (
            O => \N__16562\,
            I => \N__16559\
        );

    \I__3543\ : Odrv12
    port map (
            O => \N__16559\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__3542\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16553\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__16553\,
            I => \M_this_sprites_address_q_3_ns_1_10\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16550\,
            I => \N__16547\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__16547\,
            I => \N__16544\
        );

    \I__3538\ : Odrv12
    port map (
            O => \N__16544\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_10\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__16541\,
            I => \N__16538\
        );

    \I__3536\ : CascadeBuf
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__16535\,
            I => \N__16532\
        );

    \I__3534\ : CascadeBuf
    port map (
            O => \N__16532\,
            I => \N__16529\
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__16529\,
            I => \N__16526\
        );

    \I__3532\ : CascadeBuf
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__3530\ : CascadeBuf
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__3528\ : CascadeBuf
    port map (
            O => \N__16514\,
            I => \N__16511\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__16511\,
            I => \N__16508\
        );

    \I__3526\ : CascadeBuf
    port map (
            O => \N__16508\,
            I => \N__16505\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__3524\ : CascadeBuf
    port map (
            O => \N__16502\,
            I => \N__16499\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__16499\,
            I => \N__16496\
        );

    \I__3522\ : CascadeBuf
    port map (
            O => \N__16496\,
            I => \N__16493\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__16493\,
            I => \N__16490\
        );

    \I__3520\ : CascadeBuf
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__16487\,
            I => \N__16484\
        );

    \I__3518\ : CascadeBuf
    port map (
            O => \N__16484\,
            I => \N__16481\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__16481\,
            I => \N__16478\
        );

    \I__3516\ : CascadeBuf
    port map (
            O => \N__16478\,
            I => \N__16475\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__16475\,
            I => \N__16472\
        );

    \I__3514\ : CascadeBuf
    port map (
            O => \N__16472\,
            I => \N__16469\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__16469\,
            I => \N__16466\
        );

    \I__3512\ : CascadeBuf
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__16463\,
            I => \N__16460\
        );

    \I__3510\ : CascadeBuf
    port map (
            O => \N__16460\,
            I => \N__16457\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__16457\,
            I => \N__16454\
        );

    \I__3508\ : CascadeBuf
    port map (
            O => \N__16454\,
            I => \N__16451\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__3506\ : InMux
    port map (
            O => \N__16448\,
            I => \N__16445\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__16445\,
            I => \N__16441\
        );

    \I__3504\ : InMux
    port map (
            O => \N__16444\,
            I => \N__16438\
        );

    \I__3503\ : Sp12to4
    port map (
            O => \N__16441\,
            I => \N__16434\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__16438\,
            I => \N__16431\
        );

    \I__3501\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16428\
        );

    \I__3500\ : Span12Mux_h
    port map (
            O => \N__16434\,
            I => \N__16425\
        );

    \I__3499\ : Odrv12
    port map (
            O => \N__16431\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__16428\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__3497\ : Odrv12
    port map (
            O => \N__16425\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__3496\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16405\
        );

    \I__3495\ : InMux
    port map (
            O => \N__16417\,
            I => \N__16405\
        );

    \I__3494\ : InMux
    port map (
            O => \N__16416\,
            I => \N__16401\
        );

    \I__3493\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16397\
        );

    \I__3492\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16393\
        );

    \I__3491\ : InMux
    port map (
            O => \N__16413\,
            I => \N__16390\
        );

    \I__3490\ : InMux
    port map (
            O => \N__16412\,
            I => \N__16387\
        );

    \I__3489\ : InMux
    port map (
            O => \N__16411\,
            I => \N__16382\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16410\,
            I => \N__16379\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__16405\,
            I => \N__16376\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__16404\,
            I => \N__16372\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__16401\,
            I => \N__16368\
        );

    \I__3484\ : InMux
    port map (
            O => \N__16400\,
            I => \N__16365\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__16397\,
            I => \N__16362\
        );

    \I__3482\ : InMux
    port map (
            O => \N__16396\,
            I => \N__16359\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__16393\,
            I => \N__16354\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__16390\,
            I => \N__16354\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__16387\,
            I => \N__16351\
        );

    \I__3478\ : InMux
    port map (
            O => \N__16386\,
            I => \N__16348\
        );

    \I__3477\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16345\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__16382\,
            I => \N__16338\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__16379\,
            I => \N__16338\
        );

    \I__3474\ : Span4Mux_v
    port map (
            O => \N__16376\,
            I => \N__16338\
        );

    \I__3473\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16335\
        );

    \I__3472\ : InMux
    port map (
            O => \N__16372\,
            I => \N__16332\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16329\
        );

    \I__3470\ : Span4Mux_v
    port map (
            O => \N__16368\,
            I => \N__16324\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__16365\,
            I => \N__16324\
        );

    \I__3468\ : Span4Mux_v
    port map (
            O => \N__16362\,
            I => \N__16313\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__16359\,
            I => \N__16313\
        );

    \I__3466\ : Span4Mux_v
    port map (
            O => \N__16354\,
            I => \N__16313\
        );

    \I__3465\ : Span4Mux_v
    port map (
            O => \N__16351\,
            I => \N__16313\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__16348\,
            I => \N__16313\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__16345\,
            I => \N__16310\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__16338\,
            I => \N__16305\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__16335\,
            I => \N__16305\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__16332\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__16329\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3458\ : Odrv4
    port map (
            O => \N__16324\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__16313\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__16310\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3455\ : Odrv4
    port map (
            O => \N__16305\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__3454\ : InMux
    port map (
            O => \N__16292\,
            I => \N__16289\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__16289\,
            I => \N_202\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16280\
        );

    \I__3451\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16280\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__16280\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__3449\ : InMux
    port map (
            O => \N__16277\,
            I => \N__16272\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16276\,
            I => \N__16269\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16275\,
            I => \N__16266\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__16272\,
            I => \N__16263\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__16269\,
            I => \N_233\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__16266\,
            I => \N_233\
        );

    \I__3443\ : Odrv4
    port map (
            O => \N__16263\,
            I => \N_233\
        );

    \I__3442\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16253\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__16253\,
            I => \N__16250\
        );

    \I__3440\ : Span4Mux_h
    port map (
            O => \N__16250\,
            I => \N__16244\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__16249\,
            I => \N__16241\
        );

    \I__3438\ : InMux
    port map (
            O => \N__16248\,
            I => \N__16236\
        );

    \I__3437\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16236\
        );

    \I__3436\ : Span4Mux_h
    port map (
            O => \N__16244\,
            I => \N__16233\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16230\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__16236\,
            I => \N__16227\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__16233\,
            I => \M_this_start_address_delay_out_0\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__16230\,
            I => \M_this_start_address_delay_out_0\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__16227\,
            I => \M_this_start_address_delay_out_0\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__16220\,
            I => \M_this_state_q_srsts_i_1_1_cascade_\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16210\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16205\
        );

    \I__3427\ : InMux
    port map (
            O => \N__16215\,
            I => \N__16205\
        );

    \I__3426\ : InMux
    port map (
            O => \N__16214\,
            I => \N__16201\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16198\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__16210\,
            I => \N__16193\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__16205\,
            I => \N__16193\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16204\,
            I => \N__16190\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__16201\,
            I => \N__16185\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__16198\,
            I => \N__16185\
        );

    \I__3419\ : Span4Mux_h
    port map (
            O => \N__16193\,
            I => \N__16182\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__16190\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__3417\ : Odrv12
    port map (
            O => \N__16185\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__16182\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__16175\,
            I => \N__16171\
        );

    \I__3414\ : InMux
    port map (
            O => \N__16174\,
            I => \N__16167\
        );

    \I__3413\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16162\
        );

    \I__3412\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16162\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__16167\,
            I => \N__16153\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__16162\,
            I => \N__16153\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16161\,
            I => \N__16144\
        );

    \I__3408\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16144\
        );

    \I__3407\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16144\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16158\,
            I => \N__16144\
        );

    \I__3405\ : Span4Mux_h
    port map (
            O => \N__16153\,
            I => \N__16141\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__16144\,
            I => \N__16138\
        );

    \I__3403\ : Odrv4
    port map (
            O => \N__16141\,
            I => \this_ppu.N_250_1\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__16138\,
            I => \this_ppu.N_250_1\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16133\,
            I => \N__16124\
        );

    \I__3400\ : InMux
    port map (
            O => \N__16132\,
            I => \N__16124\
        );

    \I__3399\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16124\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__16124\,
            I => \N__16121\
        );

    \I__3397\ : Span4Mux_h
    port map (
            O => \N__16121\,
            I => \N__16116\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16120\,
            I => \N__16113\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16110\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__16116\,
            I => \this_ppu.M_last_q_RNI5NOQ4\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__16113\,
            I => \this_ppu.M_last_q_RNI5NOQ4\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__16110\,
            I => \this_ppu.M_last_q_RNI5NOQ4\
        );

    \I__3391\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16098\
        );

    \I__3390\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16093\
        );

    \I__3389\ : InMux
    port map (
            O => \N__16101\,
            I => \N__16093\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__16098\,
            I => \this_ppu.un1_M_vaddress_q_c3\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__16093\,
            I => \this_ppu.un1_M_vaddress_q_c3\
        );

    \I__3386\ : InMux
    port map (
            O => \N__16088\,
            I => \N__16085\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__16085\,
            I => \this_ppu.un1_M_haddress_q_c5\
        );

    \I__3384\ : InMux
    port map (
            O => \N__16082\,
            I => \N__16076\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16076\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__16076\,
            I => \this_ppu.un1_M_haddress_q_c2\
        );

    \I__3381\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16068\
        );

    \I__3380\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16065\
        );

    \I__3379\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16062\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__16068\,
            I => \this_ppu.un1_M_vaddress_q_c1\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__16065\,
            I => \this_ppu.un1_M_vaddress_q_c1\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16062\,
            I => \this_ppu.un1_M_vaddress_q_c1\
        );

    \I__3375\ : InMux
    port map (
            O => \N__16055\,
            I => \N__16046\
        );

    \I__3374\ : InMux
    port map (
            O => \N__16054\,
            I => \N__16046\
        );

    \I__3373\ : InMux
    port map (
            O => \N__16053\,
            I => \N__16046\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__16046\,
            I => \N__16042\
        );

    \I__3371\ : InMux
    port map (
            O => \N__16045\,
            I => \N__16039\
        );

    \I__3370\ : Span4Mux_v
    port map (
            O => \N__16042\,
            I => \N__16036\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__16039\,
            I => \N__16033\
        );

    \I__3368\ : Span4Mux_v
    port map (
            O => \N__16036\,
            I => \N__16030\
        );

    \I__3367\ : Sp12to4
    port map (
            O => \N__16033\,
            I => \N__16027\
        );

    \I__3366\ : IoSpan4Mux
    port map (
            O => \N__16030\,
            I => \N__16024\
        );

    \I__3365\ : Odrv12
    port map (
            O => \N__16027\,
            I => port_address_in_0
        );

    \I__3364\ : Odrv4
    port map (
            O => \N__16024\,
            I => port_address_in_0
        );

    \I__3363\ : InMux
    port map (
            O => \N__16019\,
            I => \N__16013\
        );

    \I__3362\ : InMux
    port map (
            O => \N__16018\,
            I => \N__16006\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16017\,
            I => \N__16006\
        );

    \I__3360\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16006\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__16013\,
            I => \N__16003\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__16006\,
            I => \N__16000\
        );

    \I__3357\ : Span4Mux_v
    port map (
            O => \N__16003\,
            I => \N__15997\
        );

    \I__3356\ : Span4Mux_v
    port map (
            O => \N__16000\,
            I => \N__15994\
        );

    \I__3355\ : Sp12to4
    port map (
            O => \N__15997\,
            I => \N__15991\
        );

    \I__3354\ : Sp12to4
    port map (
            O => \N__15994\,
            I => \N__15988\
        );

    \I__3353\ : Span12Mux_h
    port map (
            O => \N__15991\,
            I => \N__15985\
        );

    \I__3352\ : Span12Mux_h
    port map (
            O => \N__15988\,
            I => \N__15982\
        );

    \I__3351\ : Odrv12
    port map (
            O => \N__15985\,
            I => port_address_in_1
        );

    \I__3350\ : Odrv12
    port map (
            O => \N__15982\,
            I => port_address_in_1
        );

    \I__3349\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15968\
        );

    \I__3348\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15968\
        );

    \I__3347\ : InMux
    port map (
            O => \N__15975\,
            I => \N__15968\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__15968\,
            I => \N__15965\
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__15965\,
            I => \N_218\
        );

    \I__3344\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15959\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__15959\,
            I => \N_204\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__15956\,
            I => \N__15952\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__15955\,
            I => \N__15949\
        );

    \I__3340\ : InMux
    port map (
            O => \N__15952\,
            I => \N__15946\
        );

    \I__3339\ : InMux
    port map (
            O => \N__15949\,
            I => \N__15943\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__15946\,
            I => \N__15940\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__15943\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__15940\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__3335\ : InMux
    port map (
            O => \N__15935\,
            I => \un1_M_this_data_count_q_cry_11\
        );

    \I__3334\ : SRMux
    port map (
            O => \N__15932\,
            I => \N__15929\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__15929\,
            I => \N__15926\
        );

    \I__3332\ : Span4Mux_v
    port map (
            O => \N__15926\,
            I => \N__15922\
        );

    \I__3331\ : SRMux
    port map (
            O => \N__15925\,
            I => \N__15919\
        );

    \I__3330\ : Span4Mux_h
    port map (
            O => \N__15922\,
            I => \N__15916\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__15919\,
            I => \N__15913\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__15916\,
            I => \M_this_state_q_RNI20CEZ0Z_0\
        );

    \I__3327\ : Odrv12
    port map (
            O => \N__15913\,
            I => \M_this_state_q_RNI20CEZ0Z_0\
        );

    \I__3326\ : SRMux
    port map (
            O => \N__15908\,
            I => \N__15899\
        );

    \I__3325\ : SRMux
    port map (
            O => \N__15907\,
            I => \N__15896\
        );

    \I__3324\ : SRMux
    port map (
            O => \N__15906\,
            I => \N__15893\
        );

    \I__3323\ : SRMux
    port map (
            O => \N__15905\,
            I => \N__15890\
        );

    \I__3322\ : SRMux
    port map (
            O => \N__15904\,
            I => \N__15884\
        );

    \I__3321\ : SRMux
    port map (
            O => \N__15903\,
            I => \N__15877\
        );

    \I__3320\ : SRMux
    port map (
            O => \N__15902\,
            I => \N__15872\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__15899\,
            I => \N__15869\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__15896\,
            I => \N__15866\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__15893\,
            I => \N__15861\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__15890\,
            I => \N__15861\
        );

    \I__3315\ : SRMux
    port map (
            O => \N__15889\,
            I => \N__15858\
        );

    \I__3314\ : SRMux
    port map (
            O => \N__15888\,
            I => \N__15855\
        );

    \I__3313\ : SRMux
    port map (
            O => \N__15887\,
            I => \N__15850\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__15884\,
            I => \N__15845\
        );

    \I__3311\ : SRMux
    port map (
            O => \N__15883\,
            I => \N__15842\
        );

    \I__3310\ : SRMux
    port map (
            O => \N__15882\,
            I => \N__15837\
        );

    \I__3309\ : SRMux
    port map (
            O => \N__15881\,
            I => \N__15834\
        );

    \I__3308\ : SRMux
    port map (
            O => \N__15880\,
            I => \N__15831\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__15877\,
            I => \N__15826\
        );

    \I__3306\ : SRMux
    port map (
            O => \N__15876\,
            I => \N__15823\
        );

    \I__3305\ : SRMux
    port map (
            O => \N__15875\,
            I => \N__15820\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__15872\,
            I => \N__15817\
        );

    \I__3303\ : Span4Mux_s3_v
    port map (
            O => \N__15869\,
            I => \N__15806\
        );

    \I__3302\ : Span4Mux_h
    port map (
            O => \N__15866\,
            I => \N__15806\
        );

    \I__3301\ : Span4Mux_s3_v
    port map (
            O => \N__15861\,
            I => \N__15806\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__15858\,
            I => \N__15806\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__15855\,
            I => \N__15806\
        );

    \I__3298\ : SRMux
    port map (
            O => \N__15854\,
            I => \N__15803\
        );

    \I__3297\ : SRMux
    port map (
            O => \N__15853\,
            I => \N__15800\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__15850\,
            I => \N__15794\
        );

    \I__3295\ : SRMux
    port map (
            O => \N__15849\,
            I => \N__15791\
        );

    \I__3294\ : SRMux
    port map (
            O => \N__15848\,
            I => \N__15787\
        );

    \I__3293\ : Span4Mux_h
    port map (
            O => \N__15845\,
            I => \N__15781\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__15842\,
            I => \N__15781\
        );

    \I__3291\ : SRMux
    port map (
            O => \N__15841\,
            I => \N__15778\
        );

    \I__3290\ : SRMux
    port map (
            O => \N__15840\,
            I => \N__15775\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__15837\,
            I => \N__15769\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__15834\,
            I => \N__15769\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__15831\,
            I => \N__15766\
        );

    \I__3286\ : SRMux
    port map (
            O => \N__15830\,
            I => \N__15763\
        );

    \I__3285\ : SRMux
    port map (
            O => \N__15829\,
            I => \N__15760\
        );

    \I__3284\ : Span4Mux_v
    port map (
            O => \N__15826\,
            I => \N__15753\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__15823\,
            I => \N__15753\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__15820\,
            I => \N__15750\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__15817\,
            I => \N__15741\
        );

    \I__3280\ : Span4Mux_v
    port map (
            O => \N__15806\,
            I => \N__15741\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__15803\,
            I => \N__15741\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__15800\,
            I => \N__15741\
        );

    \I__3277\ : SRMux
    port map (
            O => \N__15799\,
            I => \N__15738\
        );

    \I__3276\ : SRMux
    port map (
            O => \N__15798\,
            I => \N__15735\
        );

    \I__3275\ : IoInMux
    port map (
            O => \N__15797\,
            I => \N__15730\
        );

    \I__3274\ : Span4Mux_v
    port map (
            O => \N__15794\,
            I => \N__15727\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__15791\,
            I => \N__15724\
        );

    \I__3272\ : SRMux
    port map (
            O => \N__15790\,
            I => \N__15721\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__15787\,
            I => \N__15718\
        );

    \I__3270\ : SRMux
    port map (
            O => \N__15786\,
            I => \N__15715\
        );

    \I__3269\ : Span4Mux_v
    port map (
            O => \N__15781\,
            I => \N__15710\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__15778\,
            I => \N__15710\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__15775\,
            I => \N__15707\
        );

    \I__3266\ : SRMux
    port map (
            O => \N__15774\,
            I => \N__15704\
        );

    \I__3265\ : Span4Mux_v
    port map (
            O => \N__15769\,
            I => \N__15695\
        );

    \I__3264\ : Span4Mux_h
    port map (
            O => \N__15766\,
            I => \N__15695\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__15763\,
            I => \N__15695\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__15760\,
            I => \N__15695\
        );

    \I__3261\ : SRMux
    port map (
            O => \N__15759\,
            I => \N__15692\
        );

    \I__3260\ : SRMux
    port map (
            O => \N__15758\,
            I => \N__15689\
        );

    \I__3259\ : Span4Mux_v
    port map (
            O => \N__15753\,
            I => \N__15677\
        );

    \I__3258\ : Span4Mux_h
    port map (
            O => \N__15750\,
            I => \N__15677\
        );

    \I__3257\ : Span4Mux_v
    port map (
            O => \N__15741\,
            I => \N__15677\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__15738\,
            I => \N__15677\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__15735\,
            I => \N__15677\
        );

    \I__3254\ : SRMux
    port map (
            O => \N__15734\,
            I => \N__15674\
        );

    \I__3253\ : SRMux
    port map (
            O => \N__15733\,
            I => \N__15671\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__15730\,
            I => \N__15665\
        );

    \I__3251\ : Span4Mux_h
    port map (
            O => \N__15727\,
            I => \N__15660\
        );

    \I__3250\ : Span4Mux_v
    port map (
            O => \N__15724\,
            I => \N__15660\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__15721\,
            I => \N__15657\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__15718\,
            I => \N__15652\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__15715\,
            I => \N__15652\
        );

    \I__3246\ : Span4Mux_v
    port map (
            O => \N__15710\,
            I => \N__15645\
        );

    \I__3245\ : Span4Mux_h
    port map (
            O => \N__15707\,
            I => \N__15645\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__15704\,
            I => \N__15645\
        );

    \I__3243\ : Span4Mux_v
    port map (
            O => \N__15695\,
            I => \N__15638\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__15692\,
            I => \N__15638\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__15689\,
            I => \N__15638\
        );

    \I__3240\ : SRMux
    port map (
            O => \N__15688\,
            I => \N__15635\
        );

    \I__3239\ : Span4Mux_v
    port map (
            O => \N__15677\,
            I => \N__15628\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__15674\,
            I => \N__15628\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__15671\,
            I => \N__15628\
        );

    \I__3236\ : InMux
    port map (
            O => \N__15670\,
            I => \N__15625\
        );

    \I__3235\ : InMux
    port map (
            O => \N__15669\,
            I => \N__15620\
        );

    \I__3234\ : InMux
    port map (
            O => \N__15668\,
            I => \N__15620\
        );

    \I__3233\ : Span4Mux_s1_h
    port map (
            O => \N__15665\,
            I => \N__15617\
        );

    \I__3232\ : Sp12to4
    port map (
            O => \N__15660\,
            I => \N__15614\
        );

    \I__3231\ : Span4Mux_h
    port map (
            O => \N__15657\,
            I => \N__15611\
        );

    \I__3230\ : Span4Mux_v
    port map (
            O => \N__15652\,
            I => \N__15606\
        );

    \I__3229\ : Span4Mux_v
    port map (
            O => \N__15645\,
            I => \N__15606\
        );

    \I__3228\ : Span4Mux_v
    port map (
            O => \N__15638\,
            I => \N__15599\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__15635\,
            I => \N__15599\
        );

    \I__3226\ : Span4Mux_v
    port map (
            O => \N__15628\,
            I => \N__15599\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__15625\,
            I => \N__15594\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15620\,
            I => \N__15594\
        );

    \I__3223\ : Sp12to4
    port map (
            O => \N__15617\,
            I => \N__15591\
        );

    \I__3222\ : Span12Mux_s9_h
    port map (
            O => \N__15614\,
            I => \N__15588\
        );

    \I__3221\ : Span4Mux_v
    port map (
            O => \N__15611\,
            I => \N__15581\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__15606\,
            I => \N__15581\
        );

    \I__3219\ : Span4Mux_h
    port map (
            O => \N__15599\,
            I => \N__15581\
        );

    \I__3218\ : Span4Mux_h
    port map (
            O => \N__15594\,
            I => \N__15578\
        );

    \I__3217\ : Span12Mux_v
    port map (
            O => \N__15591\,
            I => \N__15575\
        );

    \I__3216\ : Span12Mux_v
    port map (
            O => \N__15588\,
            I => \N__15570\
        );

    \I__3215\ : Sp12to4
    port map (
            O => \N__15581\,
            I => \N__15570\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__15578\,
            I => \N__15567\
        );

    \I__3213\ : Odrv12
    port map (
            O => \N__15575\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3212\ : Odrv12
    port map (
            O => \N__15570\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__15567\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3210\ : InMux
    port map (
            O => \N__15560\,
            I => \bfn_17_25_0_\
        );

    \I__3209\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15553\
        );

    \I__3208\ : InMux
    port map (
            O => \N__15556\,
            I => \N__15550\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__15553\,
            I => \N__15547\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__15550\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__15547\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__15542\,
            I => \this_ppu.un1_M_haddress_q_c2_cascade_\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__15539\,
            I => \this_ppu.un1_M_haddress_q_c5_cascade_\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__15536\,
            I => \N__15532\
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__15535\,
            I => \N__15529\
        );

    \I__3200\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15526\
        );

    \I__3199\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15523\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__15526\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__15523\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15518\,
            I => \un1_M_this_data_count_q_cry_3\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__15515\,
            I => \N__15512\
        );

    \I__3194\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15508\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15505\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__15508\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__15505\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__3190\ : InMux
    port map (
            O => \N__15500\,
            I => \un1_M_this_data_count_q_cry_4\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__15497\,
            I => \N__15494\
        );

    \I__3188\ : InMux
    port map (
            O => \N__15494\,
            I => \N__15490\
        );

    \I__3187\ : InMux
    port map (
            O => \N__15493\,
            I => \N__15487\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__15490\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__15487\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__3184\ : InMux
    port map (
            O => \N__15482\,
            I => \un1_M_this_data_count_q_cry_5\
        );

    \I__3183\ : CascadeMux
    port map (
            O => \N__15479\,
            I => \N__15476\
        );

    \I__3182\ : InMux
    port map (
            O => \N__15476\,
            I => \N__15472\
        );

    \I__3181\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15469\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__15472\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__15469\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__3178\ : InMux
    port map (
            O => \N__15464\,
            I => \un1_M_this_data_count_q_cry_6\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__15461\,
            I => \N__15457\
        );

    \I__3176\ : InMux
    port map (
            O => \N__15460\,
            I => \N__15454\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15451\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__15454\,
            I => \N__15448\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__15451\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__3172\ : Odrv4
    port map (
            O => \N__15448\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15443\,
            I => \bfn_17_24_0_\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__15440\,
            I => \N__15436\
        );

    \I__3169\ : InMux
    port map (
            O => \N__15439\,
            I => \N__15433\
        );

    \I__3168\ : InMux
    port map (
            O => \N__15436\,
            I => \N__15430\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__15433\,
            I => \N__15427\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__15430\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__3165\ : Odrv4
    port map (
            O => \N__15427\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__3164\ : InMux
    port map (
            O => \N__15422\,
            I => \un1_M_this_data_count_q_cry_8\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__15419\,
            I => \N__15415\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__15418\,
            I => \N__15412\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15415\,
            I => \N__15409\
        );

    \I__3160\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15406\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__15409\,
            I => \N__15403\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__15406\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__3157\ : Odrv4
    port map (
            O => \N__15403\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__3156\ : InMux
    port map (
            O => \N__15398\,
            I => \un1_M_this_data_count_q_cry_9\
        );

    \I__3155\ : CascadeMux
    port map (
            O => \N__15395\,
            I => \N__15391\
        );

    \I__3154\ : InMux
    port map (
            O => \N__15394\,
            I => \N__15388\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15385\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__15388\,
            I => \N__15382\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__15385\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__15382\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3149\ : InMux
    port map (
            O => \N__15377\,
            I => \un1_M_this_data_count_q_cry_10\
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__15374\,
            I => \N__15371\
        );

    \I__3147\ : CascadeBuf
    port map (
            O => \N__15371\,
            I => \N__15368\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__15368\,
            I => \N__15365\
        );

    \I__3145\ : CascadeBuf
    port map (
            O => \N__15365\,
            I => \N__15362\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__15362\,
            I => \N__15359\
        );

    \I__3143\ : CascadeBuf
    port map (
            O => \N__15359\,
            I => \N__15356\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__15356\,
            I => \N__15353\
        );

    \I__3141\ : CascadeBuf
    port map (
            O => \N__15353\,
            I => \N__15350\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__15350\,
            I => \N__15347\
        );

    \I__3139\ : CascadeBuf
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__15344\,
            I => \N__15341\
        );

    \I__3137\ : CascadeBuf
    port map (
            O => \N__15341\,
            I => \N__15338\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__15338\,
            I => \N__15335\
        );

    \I__3135\ : CascadeBuf
    port map (
            O => \N__15335\,
            I => \N__15332\
        );

    \I__3134\ : CascadeMux
    port map (
            O => \N__15332\,
            I => \N__15329\
        );

    \I__3133\ : CascadeBuf
    port map (
            O => \N__15329\,
            I => \N__15326\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__15326\,
            I => \N__15323\
        );

    \I__3131\ : CascadeBuf
    port map (
            O => \N__15323\,
            I => \N__15320\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__15320\,
            I => \N__15317\
        );

    \I__3129\ : CascadeBuf
    port map (
            O => \N__15317\,
            I => \N__15314\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__15314\,
            I => \N__15311\
        );

    \I__3127\ : CascadeBuf
    port map (
            O => \N__15311\,
            I => \N__15308\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__15308\,
            I => \N__15305\
        );

    \I__3125\ : CascadeBuf
    port map (
            O => \N__15305\,
            I => \N__15302\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__15302\,
            I => \N__15299\
        );

    \I__3123\ : CascadeBuf
    port map (
            O => \N__15299\,
            I => \N__15296\
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__15296\,
            I => \N__15293\
        );

    \I__3121\ : CascadeBuf
    port map (
            O => \N__15293\,
            I => \N__15290\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__15290\,
            I => \N__15287\
        );

    \I__3119\ : CascadeBuf
    port map (
            O => \N__15287\,
            I => \N__15284\
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__15284\,
            I => \N__15280\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15283\,
            I => \N__15277\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15280\,
            I => \N__15274\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__15277\,
            I => \N__15271\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__15274\,
            I => \N__15267\
        );

    \I__3113\ : Span4Mux_h
    port map (
            O => \N__15271\,
            I => \N__15264\
        );

    \I__3112\ : InMux
    port map (
            O => \N__15270\,
            I => \N__15261\
        );

    \I__3111\ : Span12Mux_s11_v
    port map (
            O => \N__15267\,
            I => \N__15258\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__15264\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15261\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__3108\ : Odrv12
    port map (
            O => \N__15258\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__3107\ : InMux
    port map (
            O => \N__15251\,
            I => \N__15248\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__15248\,
            I => \M_this_sprites_address_q_3_ns_1_0\
        );

    \I__3105\ : InMux
    port map (
            O => \N__15245\,
            I => \N__15242\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__15242\,
            I => \M_this_state_q_srsts_i_a2_1_8_1\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__15239\,
            I => \M_this_state_q_srsts_i_a2_1_7_1_cascade_\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15236\,
            I => \N__15233\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__15233\,
            I => \M_this_state_q_srsts_i_a2_1_9_1\
        );

    \I__3100\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15227\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__15227\,
            I => \M_this_state_q_srsts_i_a2_1_6_1\
        );

    \I__3098\ : CascadeMux
    port map (
            O => \N__15224\,
            I => \N__15221\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15217\
        );

    \I__3096\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15214\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15217\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__15214\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__15209\,
            I => \N__15206\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15202\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15199\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__15202\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__15199\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15194\,
            I => \un1_M_this_data_count_q_cry_0\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__15191\,
            I => \N__15188\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15184\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15181\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__15184\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__15181\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3082\ : InMux
    port map (
            O => \N__15176\,
            I => \un1_M_this_data_count_q_cry_1\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__15173\,
            I => \N__15170\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15170\,
            I => \N__15166\
        );

    \I__3079\ : InMux
    port map (
            O => \N__15169\,
            I => \N__15163\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__15166\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__15163\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3076\ : InMux
    port map (
            O => \N__15158\,
            I => \un1_M_this_data_count_q_cry_2\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15155\,
            I => \N__15152\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__15152\,
            I => \this_ppu.M_haddress_d8lto6_4\
        );

    \I__3073\ : InMux
    port map (
            O => \N__15149\,
            I => \N__15146\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__15146\,
            I => \this_ppu.un1_M_line_clk_out_ns_1_0\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15143\,
            I => \N__15140\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__15140\,
            I => \N__15134\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15129\
        );

    \I__3068\ : InMux
    port map (
            O => \N__15138\,
            I => \N__15129\
        );

    \I__3067\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15126\
        );

    \I__3066\ : Span4Mux_v
    port map (
            O => \N__15134\,
            I => \N__15121\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__15129\,
            I => \N__15121\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__15126\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__15121\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__15116\,
            I => \N__15111\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__15115\,
            I => \N__15108\
        );

    \I__3060\ : CascadeMux
    port map (
            O => \N__15114\,
            I => \N__15105\
        );

    \I__3059\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15102\
        );

    \I__3058\ : InMux
    port map (
            O => \N__15108\,
            I => \N__15096\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15096\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__15102\,
            I => \N__15093\
        );

    \I__3055\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15090\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__15096\,
            I => \N__15087\
        );

    \I__3053\ : Span4Mux_h
    port map (
            O => \N__15093\,
            I => \N__15084\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__15090\,
            I => \this_ppu.line_clk.M_last_qZ0\
        );

    \I__3051\ : Odrv12
    port map (
            O => \N__15087\,
            I => \this_ppu.line_clk.M_last_qZ0\
        );

    \I__3050\ : Odrv4
    port map (
            O => \N__15084\,
            I => \this_ppu.line_clk.M_last_qZ0\
        );

    \I__3049\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15074\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__15074\,
            I => \N__15070\
        );

    \I__3047\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15067\
        );

    \I__3046\ : Span4Mux_h
    port map (
            O => \N__15070\,
            I => \N__15064\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__15067\,
            I => \N__15061\
        );

    \I__3044\ : Odrv4
    port map (
            O => \N__15064\,
            I => \this_vga_signals.M_vcounter_d8\
        );

    \I__3043\ : Odrv12
    port map (
            O => \N__15061\,
            I => \this_vga_signals.M_vcounter_d8\
        );

    \I__3042\ : SRMux
    port map (
            O => \N__15056\,
            I => \N__15052\
        );

    \I__3041\ : SRMux
    port map (
            O => \N__15055\,
            I => \N__15049\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15052\,
            I => \N__15044\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__15049\,
            I => \N__15041\
        );

    \I__3038\ : SRMux
    port map (
            O => \N__15048\,
            I => \N__15038\
        );

    \I__3037\ : InMux
    port map (
            O => \N__15047\,
            I => \N__15034\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__15044\,
            I => \N__15029\
        );

    \I__3035\ : Span4Mux_v
    port map (
            O => \N__15041\,
            I => \N__15029\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__15038\,
            I => \N__15026\
        );

    \I__3033\ : SRMux
    port map (
            O => \N__15037\,
            I => \N__15023\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__15034\,
            I => \N__15020\
        );

    \I__3031\ : Span4Mux_h
    port map (
            O => \N__15029\,
            I => \N__15016\
        );

    \I__3030\ : Span12Mux_s11_v
    port map (
            O => \N__15026\,
            I => \N__15011\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__15023\,
            I => \N__15011\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__15020\,
            I => \N__15008\
        );

    \I__3027\ : InMux
    port map (
            O => \N__15019\,
            I => \N__15005\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__15016\,
            I => \this_vga_signals.M_vcounter_q_249_0\
        );

    \I__3025\ : Odrv12
    port map (
            O => \N__15011\,
            I => \this_vga_signals.M_vcounter_q_249_0\
        );

    \I__3024\ : Odrv4
    port map (
            O => \N__15008\,
            I => \this_vga_signals.M_vcounter_q_249_0\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__15005\,
            I => \this_vga_signals.M_vcounter_q_249_0\
        );

    \I__3022\ : IoInMux
    port map (
            O => \N__14996\,
            I => \N__14993\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__14993\,
            I => \N__14990\
        );

    \I__3020\ : IoSpan4Mux
    port map (
            O => \N__14990\,
            I => \N__14987\
        );

    \I__3019\ : Span4Mux_s2_h
    port map (
            O => \N__14987\,
            I => \N__14984\
        );

    \I__3018\ : Sp12to4
    port map (
            O => \N__14984\,
            I => \N__14981\
        );

    \I__3017\ : Odrv12
    port map (
            O => \N__14981\,
            I => \this_vga_signals.M_vcounter_q_esr_RNIRO2H5Z0Z_9\
        );

    \I__3016\ : InMux
    port map (
            O => \N__14978\,
            I => \N__14975\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__14975\,
            I => \N__14972\
        );

    \I__3014\ : Span4Mux_v
    port map (
            O => \N__14972\,
            I => \N__14969\
        );

    \I__3013\ : Odrv4
    port map (
            O => \N__14969\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_0\
        );

    \I__3012\ : InMux
    port map (
            O => \N__14966\,
            I => \N__14961\
        );

    \I__3011\ : InMux
    port map (
            O => \N__14965\,
            I => \N__14956\
        );

    \I__3010\ : InMux
    port map (
            O => \N__14964\,
            I => \N__14956\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__14961\,
            I => \this_pixel_clk.M_counter_qZ0Z_0\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__14956\,
            I => \this_pixel_clk.M_counter_qZ0Z_0\
        );

    \I__3007\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14948\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__14948\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_9\
        );

    \I__3005\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14942\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__14942\,
            I => \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\
        );

    \I__3003\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14936\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__14936\,
            I => \M_this_sprites_address_q_3_ns_1_6\
        );

    \I__3001\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14930\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__14930\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_6\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__14927\,
            I => \N__14924\
        );

    \I__2998\ : CascadeBuf
    port map (
            O => \N__14924\,
            I => \N__14921\
        );

    \I__2997\ : CascadeMux
    port map (
            O => \N__14921\,
            I => \N__14918\
        );

    \I__2996\ : CascadeBuf
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__14915\,
            I => \N__14912\
        );

    \I__2994\ : CascadeBuf
    port map (
            O => \N__14912\,
            I => \N__14909\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__14909\,
            I => \N__14906\
        );

    \I__2992\ : CascadeBuf
    port map (
            O => \N__14906\,
            I => \N__14903\
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__14903\,
            I => \N__14900\
        );

    \I__2990\ : CascadeBuf
    port map (
            O => \N__14900\,
            I => \N__14897\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__14897\,
            I => \N__14894\
        );

    \I__2988\ : CascadeBuf
    port map (
            O => \N__14894\,
            I => \N__14891\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__14891\,
            I => \N__14888\
        );

    \I__2986\ : CascadeBuf
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__2985\ : CascadeMux
    port map (
            O => \N__14885\,
            I => \N__14882\
        );

    \I__2984\ : CascadeBuf
    port map (
            O => \N__14882\,
            I => \N__14879\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__14879\,
            I => \N__14876\
        );

    \I__2982\ : CascadeBuf
    port map (
            O => \N__14876\,
            I => \N__14873\
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__14873\,
            I => \N__14870\
        );

    \I__2980\ : CascadeBuf
    port map (
            O => \N__14870\,
            I => \N__14867\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__14867\,
            I => \N__14864\
        );

    \I__2978\ : CascadeBuf
    port map (
            O => \N__14864\,
            I => \N__14861\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__14861\,
            I => \N__14858\
        );

    \I__2976\ : CascadeBuf
    port map (
            O => \N__14858\,
            I => \N__14855\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__14855\,
            I => \N__14852\
        );

    \I__2974\ : CascadeBuf
    port map (
            O => \N__14852\,
            I => \N__14849\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__14849\,
            I => \N__14846\
        );

    \I__2972\ : CascadeBuf
    port map (
            O => \N__14846\,
            I => \N__14843\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__14843\,
            I => \N__14840\
        );

    \I__2970\ : CascadeBuf
    port map (
            O => \N__14840\,
            I => \N__14837\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__14837\,
            I => \N__14834\
        );

    \I__2968\ : InMux
    port map (
            O => \N__14834\,
            I => \N__14831\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__14831\,
            I => \N__14826\
        );

    \I__2966\ : InMux
    port map (
            O => \N__14830\,
            I => \N__14823\
        );

    \I__2965\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14820\
        );

    \I__2964\ : Span12Mux_s9_v
    port map (
            O => \N__14826\,
            I => \N__14817\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__14823\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__14820\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__2961\ : Odrv12
    port map (
            O => \N__14817\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__14810\,
            I => \N__14807\
        );

    \I__2959\ : CascadeBuf
    port map (
            O => \N__14807\,
            I => \N__14804\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__14804\,
            I => \N__14801\
        );

    \I__2957\ : CascadeBuf
    port map (
            O => \N__14801\,
            I => \N__14798\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__14798\,
            I => \N__14795\
        );

    \I__2955\ : CascadeBuf
    port map (
            O => \N__14795\,
            I => \N__14792\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__14792\,
            I => \N__14789\
        );

    \I__2953\ : CascadeBuf
    port map (
            O => \N__14789\,
            I => \N__14786\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__14786\,
            I => \N__14783\
        );

    \I__2951\ : CascadeBuf
    port map (
            O => \N__14783\,
            I => \N__14780\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__14780\,
            I => \N__14777\
        );

    \I__2949\ : CascadeBuf
    port map (
            O => \N__14777\,
            I => \N__14774\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__14774\,
            I => \N__14771\
        );

    \I__2947\ : CascadeBuf
    port map (
            O => \N__14771\,
            I => \N__14768\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__14768\,
            I => \N__14765\
        );

    \I__2945\ : CascadeBuf
    port map (
            O => \N__14765\,
            I => \N__14762\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__14762\,
            I => \N__14759\
        );

    \I__2943\ : CascadeBuf
    port map (
            O => \N__14759\,
            I => \N__14756\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__14756\,
            I => \N__14753\
        );

    \I__2941\ : CascadeBuf
    port map (
            O => \N__14753\,
            I => \N__14750\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__14750\,
            I => \N__14747\
        );

    \I__2939\ : CascadeBuf
    port map (
            O => \N__14747\,
            I => \N__14744\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__14744\,
            I => \N__14741\
        );

    \I__2937\ : CascadeBuf
    port map (
            O => \N__14741\,
            I => \N__14738\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__14738\,
            I => \N__14735\
        );

    \I__2935\ : CascadeBuf
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__14732\,
            I => \N__14729\
        );

    \I__2933\ : CascadeBuf
    port map (
            O => \N__14729\,
            I => \N__14726\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__14726\,
            I => \N__14723\
        );

    \I__2931\ : CascadeBuf
    port map (
            O => \N__14723\,
            I => \N__14720\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__14720\,
            I => \N__14717\
        );

    \I__2929\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14714\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__14714\,
            I => \N__14711\
        );

    \I__2927\ : Span4Mux_s2_v
    port map (
            O => \N__14711\,
            I => \N__14708\
        );

    \I__2926\ : Span4Mux_h
    port map (
            O => \N__14708\,
            I => \N__14705\
        );

    \I__2925\ : Span4Mux_h
    port map (
            O => \N__14705\,
            I => \N__14700\
        );

    \I__2924\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14697\
        );

    \I__2923\ : InMux
    port map (
            O => \N__14703\,
            I => \N__14694\
        );

    \I__2922\ : Span4Mux_v
    port map (
            O => \N__14700\,
            I => \N__14691\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__14697\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__14694\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__14691\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__14684\,
            I => \N__14681\
        );

    \I__2917\ : InMux
    port map (
            O => \N__14681\,
            I => \N__14678\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__14678\,
            I => \N__14675\
        );

    \I__2915\ : Odrv4
    port map (
            O => \N__14675\,
            I => \M_this_sprites_address_q_3_ns_1_9\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__14672\,
            I => \N__14669\
        );

    \I__2913\ : CascadeBuf
    port map (
            O => \N__14669\,
            I => \N__14666\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__14666\,
            I => \N__14663\
        );

    \I__2911\ : CascadeBuf
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__14660\,
            I => \N__14657\
        );

    \I__2909\ : CascadeBuf
    port map (
            O => \N__14657\,
            I => \N__14654\
        );

    \I__2908\ : CascadeMux
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__2907\ : CascadeBuf
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__14648\,
            I => \N__14645\
        );

    \I__2905\ : CascadeBuf
    port map (
            O => \N__14645\,
            I => \N__14642\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__14642\,
            I => \N__14639\
        );

    \I__2903\ : CascadeBuf
    port map (
            O => \N__14639\,
            I => \N__14636\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__14636\,
            I => \N__14633\
        );

    \I__2901\ : CascadeBuf
    port map (
            O => \N__14633\,
            I => \N__14630\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__14630\,
            I => \N__14627\
        );

    \I__2899\ : CascadeBuf
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__14624\,
            I => \N__14621\
        );

    \I__2897\ : CascadeBuf
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__14618\,
            I => \N__14615\
        );

    \I__2895\ : CascadeBuf
    port map (
            O => \N__14615\,
            I => \N__14612\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__14612\,
            I => \N__14609\
        );

    \I__2893\ : CascadeBuf
    port map (
            O => \N__14609\,
            I => \N__14606\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__2891\ : CascadeBuf
    port map (
            O => \N__14603\,
            I => \N__14600\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__14600\,
            I => \N__14597\
        );

    \I__2889\ : CascadeBuf
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__14594\,
            I => \N__14591\
        );

    \I__2887\ : CascadeBuf
    port map (
            O => \N__14591\,
            I => \N__14588\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__14588\,
            I => \N__14585\
        );

    \I__2885\ : CascadeBuf
    port map (
            O => \N__14585\,
            I => \N__14582\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__14582\,
            I => \N__14579\
        );

    \I__2883\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14576\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__14576\,
            I => \N__14573\
        );

    \I__2881\ : Span4Mux_h
    port map (
            O => \N__14573\,
            I => \N__14570\
        );

    \I__2880\ : Span4Mux_h
    port map (
            O => \N__14570\,
            I => \N__14566\
        );

    \I__2879\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14563\
        );

    \I__2878\ : Span4Mux_h
    port map (
            O => \N__14566\,
            I => \N__14559\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__14563\,
            I => \N__14556\
        );

    \I__2876\ : InMux
    port map (
            O => \N__14562\,
            I => \N__14553\
        );

    \I__2875\ : Span4Mux_v
    port map (
            O => \N__14559\,
            I => \N__14550\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__14556\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__14553\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__14550\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__2871\ : InMux
    port map (
            O => \N__14543\,
            I => \N__14540\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__14540\,
            I => \M_this_sprites_address_q_3_ns_1_1\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__14537\,
            I => \this_ppu.un1_M_haddress_q_c3_cascade_\
        );

    \I__2868\ : InMux
    port map (
            O => \N__14534\,
            I => \N__14528\
        );

    \I__2867\ : InMux
    port map (
            O => \N__14533\,
            I => \N__14528\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__14528\,
            I => \N__14525\
        );

    \I__2865\ : Span4Mux_v
    port map (
            O => \N__14525\,
            I => \N__14516\
        );

    \I__2864\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14505\
        );

    \I__2863\ : InMux
    port map (
            O => \N__14523\,
            I => \N__14505\
        );

    \I__2862\ : InMux
    port map (
            O => \N__14522\,
            I => \N__14505\
        );

    \I__2861\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14505\
        );

    \I__2860\ : InMux
    port map (
            O => \N__14520\,
            I => \N__14505\
        );

    \I__2859\ : IoInMux
    port map (
            O => \N__14519\,
            I => \N__14502\
        );

    \I__2858\ : Span4Mux_h
    port map (
            O => \N__14516\,
            I => \N__14498\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__14505\,
            I => \N__14495\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__14502\,
            I => \N__14492\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14489\
        );

    \I__2854\ : Sp12to4
    port map (
            O => \N__14498\,
            I => \N__14484\
        );

    \I__2853\ : Span12Mux_s8_h
    port map (
            O => \N__14495\,
            I => \N__14484\
        );

    \I__2852\ : Span12Mux_s1_v
    port map (
            O => \N__14492\,
            I => \N__14481\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__14489\,
            I => \M_this_state_q_nss_0\
        );

    \I__2850\ : Odrv12
    port map (
            O => \N__14484\,
            I => \M_this_state_q_nss_0\
        );

    \I__2849\ : Odrv12
    port map (
            O => \N__14481\,
            I => \M_this_state_q_nss_0\
        );

    \I__2848\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14468\
        );

    \I__2847\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14468\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__14468\,
            I => \this_pixel_clk.M_counter_q_i_1\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__2844\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14459\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__14459\,
            I => \N__14456\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__14456\,
            I => \N__14453\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__14453\,
            I => \M_this_state_q_srsts_i_1_2\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__14450\,
            I => \N__14447\
        );

    \I__2839\ : InMux
    port map (
            O => \N__14447\,
            I => \N__14441\
        );

    \I__2838\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14441\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__14441\,
            I => \N__14438\
        );

    \I__2836\ : Span4Mux_v
    port map (
            O => \N__14438\,
            I => \N__14435\
        );

    \I__2835\ : Sp12to4
    port map (
            O => \N__14435\,
            I => \N__14432\
        );

    \I__2834\ : Span12Mux_h
    port map (
            O => \N__14432\,
            I => \N__14428\
        );

    \I__2833\ : InMux
    port map (
            O => \N__14431\,
            I => \N__14425\
        );

    \I__2832\ : Odrv12
    port map (
            O => \N__14428\,
            I => port_rw_in
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__14425\,
            I => port_rw_in
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__14420\,
            I => \N_171_0_cascade_\
        );

    \I__2829\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14414\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__14414\,
            I => \N__14411\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__14411\,
            I => \N_176_0\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__14408\,
            I => \N__14403\
        );

    \I__2825\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14400\
        );

    \I__2824\ : InMux
    port map (
            O => \N__14406\,
            I => \N__14395\
        );

    \I__2823\ : InMux
    port map (
            O => \N__14403\,
            I => \N__14395\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__14400\,
            I => \N__14390\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__14395\,
            I => \N__14390\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__14390\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__14387\,
            I => \N__14383\
        );

    \I__2818\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14380\
        );

    \I__2817\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14377\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__14380\,
            I => \N_153_0\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__14377\,
            I => \N_153_0\
        );

    \I__2814\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14369\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__14369\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_2\
        );

    \I__2812\ : InMux
    port map (
            O => \N__14366\,
            I => \N__14361\
        );

    \I__2811\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14358\
        );

    \I__2810\ : InMux
    port map (
            O => \N__14364\,
            I => \N__14355\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__14361\,
            I => \N__14352\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__14358\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__14355\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__14352\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__2805\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14342\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__14342\,
            I => \this_vga_signals.un1_M_hcounter_d7_1_0\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__14339\,
            I => \this_vga_signals.CO0_cascade_\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14336\,
            I => \N__14331\
        );

    \I__2801\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14326\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14326\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__14331\,
            I => \N__14323\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__14326\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__14323\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14318\,
            I => \N__14315\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__14315\,
            I => \this_ppu.M_line_clk_out_0\
        );

    \I__2794\ : InMux
    port map (
            O => \N__14312\,
            I => \N__14309\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__14309\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__2792\ : InMux
    port map (
            O => \N__14306\,
            I => \N__14294\
        );

    \I__2791\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14294\
        );

    \I__2790\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14294\
        );

    \I__2789\ : InMux
    port map (
            O => \N__14303\,
            I => \N__14294\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__14294\,
            I => \N__14291\
        );

    \I__2787\ : Sp12to4
    port map (
            O => \N__14291\,
            I => \N__14288\
        );

    \I__2786\ : Span12Mux_v
    port map (
            O => \N__14288\,
            I => \N__14285\
        );

    \I__2785\ : Odrv12
    port map (
            O => \N__14285\,
            I => rst_n_c
        );

    \I__2784\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14279\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__14279\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__2782\ : InMux
    port map (
            O => \N__14276\,
            I => \N__14273\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__14273\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__2780\ : InMux
    port map (
            O => \N__14270\,
            I => \N__14247\
        );

    \I__2779\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14247\
        );

    \I__2778\ : InMux
    port map (
            O => \N__14268\,
            I => \N__14247\
        );

    \I__2777\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14247\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14240\
        );

    \I__2775\ : InMux
    port map (
            O => \N__14265\,
            I => \N__14240\
        );

    \I__2774\ : InMux
    port map (
            O => \N__14264\,
            I => \N__14240\
        );

    \I__2773\ : InMux
    port map (
            O => \N__14263\,
            I => \N__14236\
        );

    \I__2772\ : CEMux
    port map (
            O => \N__14262\,
            I => \N__14232\
        );

    \I__2771\ : InMux
    port map (
            O => \N__14261\,
            I => \N__14228\
        );

    \I__2770\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14225\
        );

    \I__2769\ : InMux
    port map (
            O => \N__14259\,
            I => \N__14220\
        );

    \I__2768\ : InMux
    port map (
            O => \N__14258\,
            I => \N__14220\
        );

    \I__2767\ : InMux
    port map (
            O => \N__14257\,
            I => \N__14215\
        );

    \I__2766\ : InMux
    port map (
            O => \N__14256\,
            I => \N__14215\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__14247\,
            I => \N__14212\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__14240\,
            I => \N__14209\
        );

    \I__2763\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14206\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__14236\,
            I => \N__14201\
        );

    \I__2761\ : InMux
    port map (
            O => \N__14235\,
            I => \N__14198\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__14232\,
            I => \N__14195\
        );

    \I__2759\ : InMux
    port map (
            O => \N__14231\,
            I => \N__14192\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__14228\,
            I => \N__14187\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__14225\,
            I => \N__14187\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__14220\,
            I => \N__14184\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__14215\,
            I => \N__14181\
        );

    \I__2754\ : Span4Mux_v
    port map (
            O => \N__14212\,
            I => \N__14178\
        );

    \I__2753\ : Span4Mux_v
    port map (
            O => \N__14209\,
            I => \N__14173\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__14206\,
            I => \N__14173\
        );

    \I__2751\ : InMux
    port map (
            O => \N__14205\,
            I => \N__14168\
        );

    \I__2750\ : InMux
    port map (
            O => \N__14204\,
            I => \N__14168\
        );

    \I__2749\ : Span12Mux_s3_h
    port map (
            O => \N__14201\,
            I => \N__14165\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__14198\,
            I => \N__14162\
        );

    \I__2747\ : Span4Mux_v
    port map (
            O => \N__14195\,
            I => \N__14159\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__14192\,
            I => \N__14154\
        );

    \I__2745\ : Span4Mux_v
    port map (
            O => \N__14187\,
            I => \N__14154\
        );

    \I__2744\ : Span4Mux_h
    port map (
            O => \N__14184\,
            I => \N__14149\
        );

    \I__2743\ : Span4Mux_h
    port map (
            O => \N__14181\,
            I => \N__14149\
        );

    \I__2742\ : Span4Mux_h
    port map (
            O => \N__14178\,
            I => \N__14144\
        );

    \I__2741\ : Span4Mux_h
    port map (
            O => \N__14173\,
            I => \N__14144\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__14168\,
            I => \N__14139\
        );

    \I__2739\ : Span12Mux_h
    port map (
            O => \N__14165\,
            I => \N__14139\
        );

    \I__2738\ : Span4Mux_v
    port map (
            O => \N__14162\,
            I => \N__14132\
        );

    \I__2737\ : Span4Mux_h
    port map (
            O => \N__14159\,
            I => \N__14132\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__14154\,
            I => \N__14132\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__14149\,
            I => \M_counter_q_RNIFKS8_1\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__14144\,
            I => \M_counter_q_RNIFKS8_1\
        );

    \I__2733\ : Odrv12
    port map (
            O => \N__14139\,
            I => \M_counter_q_RNIFKS8_1\
        );

    \I__2732\ : Odrv4
    port map (
            O => \N__14132\,
            I => \M_counter_q_RNIFKS8_1\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__14123\,
            I => \M_counter_q_RNIFKS8_1_cascade_\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__14120\,
            I => \N__14111\
        );

    \I__2729\ : InMux
    port map (
            O => \N__14119\,
            I => \N__14102\
        );

    \I__2728\ : InMux
    port map (
            O => \N__14118\,
            I => \N__14102\
        );

    \I__2727\ : InMux
    port map (
            O => \N__14117\,
            I => \N__14102\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14116\,
            I => \N__14096\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14115\,
            I => \N__14096\
        );

    \I__2724\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14093\
        );

    \I__2723\ : InMux
    port map (
            O => \N__14111\,
            I => \N__14090\
        );

    \I__2722\ : InMux
    port map (
            O => \N__14110\,
            I => \N__14085\
        );

    \I__2721\ : InMux
    port map (
            O => \N__14109\,
            I => \N__14085\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__14102\,
            I => \N__14082\
        );

    \I__2719\ : InMux
    port map (
            O => \N__14101\,
            I => \N__14079\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__14096\,
            I => \N__14076\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__14093\,
            I => \N__14071\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__14090\,
            I => \N__14071\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__14085\,
            I => \N__14068\
        );

    \I__2714\ : Span4Mux_v
    port map (
            O => \N__14082\,
            I => \N__14063\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__14079\,
            I => \N__14063\
        );

    \I__2712\ : Span4Mux_v
    port map (
            O => \N__14076\,
            I => \N__14060\
        );

    \I__2711\ : Span4Mux_v
    port map (
            O => \N__14071\,
            I => \N__14057\
        );

    \I__2710\ : Span4Mux_h
    port map (
            O => \N__14068\,
            I => \N__14054\
        );

    \I__2709\ : Span4Mux_h
    port map (
            O => \N__14063\,
            I => \N__14051\
        );

    \I__2708\ : Odrv4
    port map (
            O => \N__14060\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__14057\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__2706\ : Odrv4
    port map (
            O => \N__14054\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__2705\ : Odrv4
    port map (
            O => \N__14051\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__2704\ : InMux
    port map (
            O => \N__14042\,
            I => \un1_M_this_sprites_address_q_cry_12\
        );

    \I__2703\ : InMux
    port map (
            O => \N__14039\,
            I => \N__14036\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__14036\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_8\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__14033\,
            I => \M_this_sprites_address_q_3_ns_1_8_cascade_\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__14030\,
            I => \N__14027\
        );

    \I__2699\ : CascadeBuf
    port map (
            O => \N__14027\,
            I => \N__14024\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__14024\,
            I => \N__14021\
        );

    \I__2697\ : CascadeBuf
    port map (
            O => \N__14021\,
            I => \N__14018\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__14018\,
            I => \N__14015\
        );

    \I__2695\ : CascadeBuf
    port map (
            O => \N__14015\,
            I => \N__14012\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__14012\,
            I => \N__14009\
        );

    \I__2693\ : CascadeBuf
    port map (
            O => \N__14009\,
            I => \N__14006\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__14006\,
            I => \N__14003\
        );

    \I__2691\ : CascadeBuf
    port map (
            O => \N__14003\,
            I => \N__14000\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__14000\,
            I => \N__13997\
        );

    \I__2689\ : CascadeBuf
    port map (
            O => \N__13997\,
            I => \N__13994\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__13994\,
            I => \N__13991\
        );

    \I__2687\ : CascadeBuf
    port map (
            O => \N__13991\,
            I => \N__13988\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__13988\,
            I => \N__13985\
        );

    \I__2685\ : CascadeBuf
    port map (
            O => \N__13985\,
            I => \N__13982\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__13982\,
            I => \N__13979\
        );

    \I__2683\ : CascadeBuf
    port map (
            O => \N__13979\,
            I => \N__13976\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__13976\,
            I => \N__13973\
        );

    \I__2681\ : CascadeBuf
    port map (
            O => \N__13973\,
            I => \N__13970\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__13970\,
            I => \N__13967\
        );

    \I__2679\ : CascadeBuf
    port map (
            O => \N__13967\,
            I => \N__13964\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__2677\ : CascadeBuf
    port map (
            O => \N__13961\,
            I => \N__13958\
        );

    \I__2676\ : CascadeMux
    port map (
            O => \N__13958\,
            I => \N__13955\
        );

    \I__2675\ : CascadeBuf
    port map (
            O => \N__13955\,
            I => \N__13952\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__13952\,
            I => \N__13949\
        );

    \I__2673\ : CascadeBuf
    port map (
            O => \N__13949\,
            I => \N__13946\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__13946\,
            I => \N__13943\
        );

    \I__2671\ : CascadeBuf
    port map (
            O => \N__13943\,
            I => \N__13940\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__13940\,
            I => \N__13937\
        );

    \I__2669\ : InMux
    port map (
            O => \N__13937\,
            I => \N__13934\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__13934\,
            I => \N__13931\
        );

    \I__2667\ : Span4Mux_h
    port map (
            O => \N__13931\,
            I => \N__13928\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__13928\,
            I => \N__13925\
        );

    \I__2665\ : Span4Mux_v
    port map (
            O => \N__13925\,
            I => \N__13920\
        );

    \I__2664\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13917\
        );

    \I__2663\ : InMux
    port map (
            O => \N__13923\,
            I => \N__13914\
        );

    \I__2662\ : Span4Mux_v
    port map (
            O => \N__13920\,
            I => \N__13911\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__13917\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__13914\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__13911\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__2658\ : InMux
    port map (
            O => \N__13904\,
            I => \N__13901\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__13901\,
            I => \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_11\
        );

    \I__2656\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__13895\,
            I => \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\
        );

    \I__2654\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__13889\,
            I => \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_12\
        );

    \I__2652\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__13883\,
            I => \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\
        );

    \I__2650\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13877\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__2648\ : Odrv12
    port map (
            O => \N__13874\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_1\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__13871\,
            I => \this_vga_signals.un1_M_hcounter_d7_1_0_cascade_\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__2645\ : CascadeBuf
    port map (
            O => \N__13865\,
            I => \N__13862\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__13862\,
            I => \N__13859\
        );

    \I__2643\ : CascadeBuf
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__13856\,
            I => \N__13853\
        );

    \I__2641\ : CascadeBuf
    port map (
            O => \N__13853\,
            I => \N__13850\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__13850\,
            I => \N__13847\
        );

    \I__2639\ : CascadeBuf
    port map (
            O => \N__13847\,
            I => \N__13844\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__13844\,
            I => \N__13841\
        );

    \I__2637\ : CascadeBuf
    port map (
            O => \N__13841\,
            I => \N__13838\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__13838\,
            I => \N__13835\
        );

    \I__2635\ : CascadeBuf
    port map (
            O => \N__13835\,
            I => \N__13832\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__13832\,
            I => \N__13829\
        );

    \I__2633\ : CascadeBuf
    port map (
            O => \N__13829\,
            I => \N__13826\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__13826\,
            I => \N__13823\
        );

    \I__2631\ : CascadeBuf
    port map (
            O => \N__13823\,
            I => \N__13820\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__13820\,
            I => \N__13817\
        );

    \I__2629\ : CascadeBuf
    port map (
            O => \N__13817\,
            I => \N__13814\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__13814\,
            I => \N__13811\
        );

    \I__2627\ : CascadeBuf
    port map (
            O => \N__13811\,
            I => \N__13808\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__13808\,
            I => \N__13805\
        );

    \I__2625\ : CascadeBuf
    port map (
            O => \N__13805\,
            I => \N__13802\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__13802\,
            I => \N__13799\
        );

    \I__2623\ : CascadeBuf
    port map (
            O => \N__13799\,
            I => \N__13796\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__13796\,
            I => \N__13793\
        );

    \I__2621\ : CascadeBuf
    port map (
            O => \N__13793\,
            I => \N__13790\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__13790\,
            I => \N__13787\
        );

    \I__2619\ : CascadeBuf
    port map (
            O => \N__13787\,
            I => \N__13784\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__13784\,
            I => \N__13781\
        );

    \I__2617\ : CascadeBuf
    port map (
            O => \N__13781\,
            I => \N__13778\
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__13778\,
            I => \N__13775\
        );

    \I__2615\ : InMux
    port map (
            O => \N__13775\,
            I => \N__13772\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__13772\,
            I => \N__13767\
        );

    \I__2613\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13764\
        );

    \I__2612\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13761\
        );

    \I__2611\ : Span12Mux_h
    port map (
            O => \N__13767\,
            I => \N__13758\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__13764\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__13761\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__2608\ : Odrv12
    port map (
            O => \N__13758\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__2607\ : InMux
    port map (
            O => \N__13751\,
            I => \N__13748\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__13748\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_4\
        );

    \I__2605\ : InMux
    port map (
            O => \N__13745\,
            I => \un1_M_this_sprites_address_q_cry_3\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__13742\,
            I => \N__13739\
        );

    \I__2603\ : CascadeBuf
    port map (
            O => \N__13739\,
            I => \N__13736\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__13736\,
            I => \N__13733\
        );

    \I__2601\ : CascadeBuf
    port map (
            O => \N__13733\,
            I => \N__13730\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__13730\,
            I => \N__13727\
        );

    \I__2599\ : CascadeBuf
    port map (
            O => \N__13727\,
            I => \N__13724\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__13724\,
            I => \N__13721\
        );

    \I__2597\ : CascadeBuf
    port map (
            O => \N__13721\,
            I => \N__13718\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__13718\,
            I => \N__13715\
        );

    \I__2595\ : CascadeBuf
    port map (
            O => \N__13715\,
            I => \N__13712\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__13712\,
            I => \N__13709\
        );

    \I__2593\ : CascadeBuf
    port map (
            O => \N__13709\,
            I => \N__13706\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__13706\,
            I => \N__13703\
        );

    \I__2591\ : CascadeBuf
    port map (
            O => \N__13703\,
            I => \N__13700\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__13700\,
            I => \N__13697\
        );

    \I__2589\ : CascadeBuf
    port map (
            O => \N__13697\,
            I => \N__13694\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__13694\,
            I => \N__13691\
        );

    \I__2587\ : CascadeBuf
    port map (
            O => \N__13691\,
            I => \N__13688\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__13688\,
            I => \N__13685\
        );

    \I__2585\ : CascadeBuf
    port map (
            O => \N__13685\,
            I => \N__13682\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__13682\,
            I => \N__13679\
        );

    \I__2583\ : CascadeBuf
    port map (
            O => \N__13679\,
            I => \N__13676\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__13676\,
            I => \N__13673\
        );

    \I__2581\ : CascadeBuf
    port map (
            O => \N__13673\,
            I => \N__13670\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__13670\,
            I => \N__13667\
        );

    \I__2579\ : CascadeBuf
    port map (
            O => \N__13667\,
            I => \N__13664\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__13664\,
            I => \N__13661\
        );

    \I__2577\ : CascadeBuf
    port map (
            O => \N__13661\,
            I => \N__13658\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__13658\,
            I => \N__13655\
        );

    \I__2575\ : CascadeBuf
    port map (
            O => \N__13655\,
            I => \N__13652\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__13652\,
            I => \N__13649\
        );

    \I__2573\ : InMux
    port map (
            O => \N__13649\,
            I => \N__13646\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__13646\,
            I => \N__13643\
        );

    \I__2571\ : Span4Mux_s1_v
    port map (
            O => \N__13643\,
            I => \N__13640\
        );

    \I__2570\ : Span4Mux_h
    port map (
            O => \N__13640\,
            I => \N__13637\
        );

    \I__2569\ : Sp12to4
    port map (
            O => \N__13637\,
            I => \N__13632\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13636\,
            I => \N__13629\
        );

    \I__2567\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13626\
        );

    \I__2566\ : Span12Mux_s11_v
    port map (
            O => \N__13632\,
            I => \N__13623\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__13629\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__13626\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__2563\ : Odrv12
    port map (
            O => \N__13623\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__2562\ : InMux
    port map (
            O => \N__13616\,
            I => \N__13613\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__13613\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_5\
        );

    \I__2560\ : InMux
    port map (
            O => \N__13610\,
            I => \un1_M_this_sprites_address_q_cry_4\
        );

    \I__2559\ : InMux
    port map (
            O => \N__13607\,
            I => \un1_M_this_sprites_address_q_cry_5\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__13604\,
            I => \N__13601\
        );

    \I__2557\ : CascadeBuf
    port map (
            O => \N__13601\,
            I => \N__13598\
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__13598\,
            I => \N__13595\
        );

    \I__2555\ : CascadeBuf
    port map (
            O => \N__13595\,
            I => \N__13592\
        );

    \I__2554\ : CascadeMux
    port map (
            O => \N__13592\,
            I => \N__13589\
        );

    \I__2553\ : CascadeBuf
    port map (
            O => \N__13589\,
            I => \N__13586\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__13586\,
            I => \N__13583\
        );

    \I__2551\ : CascadeBuf
    port map (
            O => \N__13583\,
            I => \N__13580\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__13580\,
            I => \N__13577\
        );

    \I__2549\ : CascadeBuf
    port map (
            O => \N__13577\,
            I => \N__13574\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__13574\,
            I => \N__13571\
        );

    \I__2547\ : CascadeBuf
    port map (
            O => \N__13571\,
            I => \N__13568\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__13568\,
            I => \N__13565\
        );

    \I__2545\ : CascadeBuf
    port map (
            O => \N__13565\,
            I => \N__13562\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__13562\,
            I => \N__13559\
        );

    \I__2543\ : CascadeBuf
    port map (
            O => \N__13559\,
            I => \N__13556\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__13556\,
            I => \N__13553\
        );

    \I__2541\ : CascadeBuf
    port map (
            O => \N__13553\,
            I => \N__13550\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__13550\,
            I => \N__13547\
        );

    \I__2539\ : CascadeBuf
    port map (
            O => \N__13547\,
            I => \N__13544\
        );

    \I__2538\ : CascadeMux
    port map (
            O => \N__13544\,
            I => \N__13541\
        );

    \I__2537\ : CascadeBuf
    port map (
            O => \N__13541\,
            I => \N__13538\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__13538\,
            I => \N__13535\
        );

    \I__2535\ : CascadeBuf
    port map (
            O => \N__13535\,
            I => \N__13532\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__13532\,
            I => \N__13529\
        );

    \I__2533\ : CascadeBuf
    port map (
            O => \N__13529\,
            I => \N__13526\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__13526\,
            I => \N__13523\
        );

    \I__2531\ : CascadeBuf
    port map (
            O => \N__13523\,
            I => \N__13520\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__13520\,
            I => \N__13517\
        );

    \I__2529\ : CascadeBuf
    port map (
            O => \N__13517\,
            I => \N__13514\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__13514\,
            I => \N__13511\
        );

    \I__2527\ : InMux
    port map (
            O => \N__13511\,
            I => \N__13508\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13508\,
            I => \N__13505\
        );

    \I__2525\ : Sp12to4
    port map (
            O => \N__13505\,
            I => \N__13500\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13504\,
            I => \N__13497\
        );

    \I__2523\ : InMux
    port map (
            O => \N__13503\,
            I => \N__13494\
        );

    \I__2522\ : Span12Mux_s11_v
    port map (
            O => \N__13500\,
            I => \N__13491\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__13497\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__13494\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__2519\ : Odrv12
    port map (
            O => \N__13491\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13484\,
            I => \N__13481\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__13481\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_7\
        );

    \I__2516\ : InMux
    port map (
            O => \N__13478\,
            I => \un1_M_this_sprites_address_q_cry_6\
        );

    \I__2515\ : InMux
    port map (
            O => \N__13475\,
            I => \bfn_15_23_0_\
        );

    \I__2514\ : InMux
    port map (
            O => \N__13472\,
            I => \un1_M_this_sprites_address_q_cry_8\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13469\,
            I => \un1_M_this_sprites_address_q_cry_9\
        );

    \I__2512\ : InMux
    port map (
            O => \N__13466\,
            I => \un1_M_this_sprites_address_q_cry_10\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13463\,
            I => \un1_M_this_sprites_address_q_cry_11\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13460\,
            I => \N__13457\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__13457\,
            I => \M_this_ppu_vga_is_drawing_0\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__13454\,
            I => \this_ppu.M_line_clk_out_0_cascade_\
        );

    \I__2507\ : InMux
    port map (
            O => \N__13451\,
            I => \N__13448\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__13448\,
            I => \M_this_sprites_address_q_3_ns_1_5\
        );

    \I__2505\ : InMux
    port map (
            O => \N__13445\,
            I => \N__13442\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__13442\,
            I => \M_this_sprites_address_q_3_ns_1_4\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__13439\,
            I => \M_this_sprites_address_q_3_ns_1_7_cascade_\
        );

    \I__2502\ : InMux
    port map (
            O => \N__13436\,
            I => \un1_M_this_sprites_address_q_cry_0\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13433\,
            I => \un1_M_this_sprites_address_q_cry_1\
        );

    \I__2500\ : InMux
    port map (
            O => \N__13430\,
            I => \un1_M_this_sprites_address_q_cry_2\
        );

    \I__2499\ : CascadeMux
    port map (
            O => \N__13427\,
            I => \N__13420\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__13426\,
            I => \N__13414\
        );

    \I__2497\ : InMux
    port map (
            O => \N__13425\,
            I => \N__13411\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13424\,
            I => \N__13408\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13423\,
            I => \N__13405\
        );

    \I__2494\ : InMux
    port map (
            O => \N__13420\,
            I => \N__13397\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13419\,
            I => \N__13394\
        );

    \I__2492\ : InMux
    port map (
            O => \N__13418\,
            I => \N__13389\
        );

    \I__2491\ : InMux
    port map (
            O => \N__13417\,
            I => \N__13389\
        );

    \I__2490\ : InMux
    port map (
            O => \N__13414\,
            I => \N__13386\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__13411\,
            I => \N__13381\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__13408\,
            I => \N__13381\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__13405\,
            I => \N__13378\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13404\,
            I => \N__13371\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13403\,
            I => \N__13371\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13402\,
            I => \N__13371\
        );

    \I__2483\ : InMux
    port map (
            O => \N__13401\,
            I => \N__13368\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13400\,
            I => \N__13365\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__13397\,
            I => \N__13358\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__13394\,
            I => \N__13358\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__13389\,
            I => \N__13353\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__13386\,
            I => \N__13353\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__13381\,
            I => \N__13346\
        );

    \I__2476\ : Span4Mux_h
    port map (
            O => \N__13378\,
            I => \N__13346\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__13371\,
            I => \N__13346\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__13368\,
            I => \N__13343\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__13365\,
            I => \N__13340\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__13364\,
            I => \N__13336\
        );

    \I__2471\ : InMux
    port map (
            O => \N__13363\,
            I => \N__13333\
        );

    \I__2470\ : Span4Mux_v
    port map (
            O => \N__13358\,
            I => \N__13328\
        );

    \I__2469\ : Span4Mux_v
    port map (
            O => \N__13353\,
            I => \N__13328\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__13346\,
            I => \N__13325\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__13343\,
            I => \N__13320\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__13340\,
            I => \N__13320\
        );

    \I__2465\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13315\
        );

    \I__2464\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13315\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__13333\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__13328\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__13325\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__13320\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__13315\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2458\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13297\
        );

    \I__2457\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13292\
        );

    \I__2456\ : InMux
    port map (
            O => \N__13302\,
            I => \N__13292\
        );

    \I__2455\ : InMux
    port map (
            O => \N__13301\,
            I => \N__13289\
        );

    \I__2454\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13286\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__13297\,
            I => \N__13282\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__13292\,
            I => \N__13279\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__13289\,
            I => \N__13276\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__13286\,
            I => \N__13273\
        );

    \I__2449\ : InMux
    port map (
            O => \N__13285\,
            I => \N__13269\
        );

    \I__2448\ : Span4Mux_v
    port map (
            O => \N__13282\,
            I => \N__13264\
        );

    \I__2447\ : Span4Mux_h
    port map (
            O => \N__13279\,
            I => \N__13264\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__13276\,
            I => \N__13259\
        );

    \I__2445\ : Span4Mux_v
    port map (
            O => \N__13273\,
            I => \N__13259\
        );

    \I__2444\ : InMux
    port map (
            O => \N__13272\,
            I => \N__13256\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__13269\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__13264\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__13259\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__13256\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__13247\,
            I => \N__13244\
        );

    \I__2438\ : InMux
    port map (
            O => \N__13244\,
            I => \N__13241\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__13241\,
            I => \N__13238\
        );

    \I__2436\ : Span4Mux_h
    port map (
            O => \N__13238\,
            I => \N__13235\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__13235\,
            I => \this_vga_signals.g0_0\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__13232\,
            I => \N_206_cascade_\
        );

    \I__2433\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__13226\,
            I => \N_207\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13220\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__13220\,
            I => \M_this_state_q_srsts_0_a2_1_4\
        );

    \I__2429\ : IoInMux
    port map (
            O => \N__13217\,
            I => \N__13214\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__13214\,
            I => \N__13210\
        );

    \I__2427\ : InMux
    port map (
            O => \N__13213\,
            I => \N__13205\
        );

    \I__2426\ : IoSpan4Mux
    port map (
            O => \N__13210\,
            I => \N__13202\
        );

    \I__2425\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13199\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__13208\,
            I => \N__13196\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__13205\,
            I => \N__13193\
        );

    \I__2422\ : Sp12to4
    port map (
            O => \N__13202\,
            I => \N__13190\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__13199\,
            I => \N__13187\
        );

    \I__2420\ : InMux
    port map (
            O => \N__13196\,
            I => \N__13184\
        );

    \I__2419\ : Sp12to4
    port map (
            O => \N__13193\,
            I => \N__13181\
        );

    \I__2418\ : Span12Mux_h
    port map (
            O => \N__13190\,
            I => \N__13178\
        );

    \I__2417\ : Span12Mux_v
    port map (
            O => \N__13187\,
            I => \N__13175\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__13184\,
            I => \N__13170\
        );

    \I__2415\ : Span12Mux_v
    port map (
            O => \N__13181\,
            I => \N__13167\
        );

    \I__2414\ : Span12Mux_v
    port map (
            O => \N__13178\,
            I => \N__13162\
        );

    \I__2413\ : Span12Mux_h
    port map (
            O => \N__13175\,
            I => \N__13162\
        );

    \I__2412\ : InMux
    port map (
            O => \N__13174\,
            I => \N__13159\
        );

    \I__2411\ : InMux
    port map (
            O => \N__13173\,
            I => \N__13156\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__13170\,
            I => \N__13153\
        );

    \I__2409\ : Odrv12
    port map (
            O => \N__13167\,
            I => port_dmab_c
        );

    \I__2408\ : Odrv12
    port map (
            O => \N__13162\,
            I => port_dmab_c
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__13159\,
            I => port_dmab_c
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13156\,
            I => port_dmab_c
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__13153\,
            I => port_dmab_c
        );

    \I__2404\ : IoInMux
    port map (
            O => \N__13142\,
            I => \N__13138\
        );

    \I__2403\ : IoInMux
    port map (
            O => \N__13141\,
            I => \N__13135\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__13138\,
            I => \N__13130\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__13135\,
            I => \N__13130\
        );

    \I__2400\ : IoSpan4Mux
    port map (
            O => \N__13130\,
            I => \N__13126\
        );

    \I__2399\ : IoInMux
    port map (
            O => \N__13129\,
            I => \N__13121\
        );

    \I__2398\ : IoSpan4Mux
    port map (
            O => \N__13126\,
            I => \N__13117\
        );

    \I__2397\ : IoInMux
    port map (
            O => \N__13125\,
            I => \N__13114\
        );

    \I__2396\ : IoInMux
    port map (
            O => \N__13124\,
            I => \N__13111\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__13121\,
            I => \N__13106\
        );

    \I__2394\ : IoInMux
    port map (
            O => \N__13120\,
            I => \N__13103\
        );

    \I__2393\ : IoSpan4Mux
    port map (
            O => \N__13117\,
            I => \N__13092\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__13114\,
            I => \N__13092\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__13111\,
            I => \N__13092\
        );

    \I__2390\ : IoInMux
    port map (
            O => \N__13110\,
            I => \N__13089\
        );

    \I__2389\ : IoInMux
    port map (
            O => \N__13109\,
            I => \N__13086\
        );

    \I__2388\ : IoSpan4Mux
    port map (
            O => \N__13106\,
            I => \N__13081\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__13103\,
            I => \N__13081\
        );

    \I__2386\ : IoInMux
    port map (
            O => \N__13102\,
            I => \N__13078\
        );

    \I__2385\ : IoInMux
    port map (
            O => \N__13101\,
            I => \N__13075\
        );

    \I__2384\ : IoInMux
    port map (
            O => \N__13100\,
            I => \N__13072\
        );

    \I__2383\ : IoInMux
    port map (
            O => \N__13099\,
            I => \N__13069\
        );

    \I__2382\ : IoSpan4Mux
    port map (
            O => \N__13092\,
            I => \N__13061\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__13089\,
            I => \N__13061\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__13086\,
            I => \N__13061\
        );

    \I__2379\ : IoSpan4Mux
    port map (
            O => \N__13081\,
            I => \N__13056\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__13078\,
            I => \N__13056\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__13075\,
            I => \N__13053\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__13072\,
            I => \N__13049\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__13069\,
            I => \N__13046\
        );

    \I__2374\ : IoInMux
    port map (
            O => \N__13068\,
            I => \N__13043\
        );

    \I__2373\ : IoSpan4Mux
    port map (
            O => \N__13061\,
            I => \N__13036\
        );

    \I__2372\ : IoSpan4Mux
    port map (
            O => \N__13056\,
            I => \N__13036\
        );

    \I__2371\ : Span4Mux_s2_h
    port map (
            O => \N__13053\,
            I => \N__13032\
        );

    \I__2370\ : IoInMux
    port map (
            O => \N__13052\,
            I => \N__13029\
        );

    \I__2369\ : IoSpan4Mux
    port map (
            O => \N__13049\,
            I => \N__13022\
        );

    \I__2368\ : IoSpan4Mux
    port map (
            O => \N__13046\,
            I => \N__13022\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__13043\,
            I => \N__13022\
        );

    \I__2366\ : IoInMux
    port map (
            O => \N__13042\,
            I => \N__13019\
        );

    \I__2365\ : IoInMux
    port map (
            O => \N__13041\,
            I => \N__13016\
        );

    \I__2364\ : Span4Mux_s3_h
    port map (
            O => \N__13036\,
            I => \N__13013\
        );

    \I__2363\ : IoInMux
    port map (
            O => \N__13035\,
            I => \N__13010\
        );

    \I__2362\ : Span4Mux_h
    port map (
            O => \N__13032\,
            I => \N__13007\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__13029\,
            I => \N__13004\
        );

    \I__2360\ : IoSpan4Mux
    port map (
            O => \N__13022\,
            I => \N__12997\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__13019\,
            I => \N__12997\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__13016\,
            I => \N__12997\
        );

    \I__2357\ : Sp12to4
    port map (
            O => \N__13013\,
            I => \N__12992\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__13010\,
            I => \N__12992\
        );

    \I__2355\ : Span4Mux_h
    port map (
            O => \N__13007\,
            I => \N__12989\
        );

    \I__2354\ : Span12Mux_s0_v
    port map (
            O => \N__13004\,
            I => \N__12986\
        );

    \I__2353\ : IoSpan4Mux
    port map (
            O => \N__12997\,
            I => \N__12983\
        );

    \I__2352\ : Span12Mux_s11_h
    port map (
            O => \N__12992\,
            I => \N__12980\
        );

    \I__2351\ : Span4Mux_h
    port map (
            O => \N__12989\,
            I => \N__12977\
        );

    \I__2350\ : Span12Mux_h
    port map (
            O => \N__12986\,
            I => \N__12972\
        );

    \I__2349\ : Sp12to4
    port map (
            O => \N__12983\,
            I => \N__12972\
        );

    \I__2348\ : Odrv12
    port map (
            O => \N__12980\,
            I => port_dmab_c_i
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__12977\,
            I => port_dmab_c_i
        );

    \I__2346\ : Odrv12
    port map (
            O => \N__12972\,
            I => port_dmab_c_i
        );

    \I__2345\ : InMux
    port map (
            O => \N__12965\,
            I => \N__12959\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__12964\,
            I => \N__12954\
        );

    \I__2343\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12945\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__12962\,
            I => \N__12942\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__12959\,
            I => \N__12939\
        );

    \I__2340\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12936\
        );

    \I__2339\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12931\
        );

    \I__2338\ : InMux
    port map (
            O => \N__12954\,
            I => \N__12931\
        );

    \I__2337\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12926\
        );

    \I__2336\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12926\
        );

    \I__2335\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12923\
        );

    \I__2334\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12920\
        );

    \I__2333\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12917\
        );

    \I__2332\ : InMux
    port map (
            O => \N__12948\,
            I => \N__12914\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__12945\,
            I => \N__12911\
        );

    \I__2330\ : InMux
    port map (
            O => \N__12942\,
            I => \N__12908\
        );

    \I__2329\ : Span4Mux_v
    port map (
            O => \N__12939\,
            I => \N__12901\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__12936\,
            I => \N__12901\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__12931\,
            I => \N__12901\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__12926\,
            I => \N__12898\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__12923\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__12920\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__12917\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__12914\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__12911\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__12908\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__12901\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2318\ : Odrv12
    port map (
            O => \N__12898\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__12881\,
            I => \N__12878\
        );

    \I__2316\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12875\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__12875\,
            I => \N__12872\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__12872\,
            I => \N__12869\
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__12869\,
            I => \this_vga_signals.g1_0\
        );

    \I__2312\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12863\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__12863\,
            I => \N__12859\
        );

    \I__2310\ : InMux
    port map (
            O => \N__12862\,
            I => \N__12856\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__12859\,
            I => \N__12853\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__12856\,
            I => \N__12847\
        );

    \I__2307\ : Span4Mux_h
    port map (
            O => \N__12853\,
            I => \N__12847\
        );

    \I__2306\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12844\
        );

    \I__2305\ : Odrv4
    port map (
            O => \N__12847\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__12844\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__12839\,
            I => \N__12833\
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__12838\,
            I => \N__12829\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__12837\,
            I => \N__12823\
        );

    \I__2300\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12820\
        );

    \I__2299\ : InMux
    port map (
            O => \N__12833\,
            I => \N__12813\
        );

    \I__2298\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12803\
        );

    \I__2297\ : InMux
    port map (
            O => \N__12829\,
            I => \N__12794\
        );

    \I__2296\ : InMux
    port map (
            O => \N__12828\,
            I => \N__12794\
        );

    \I__2295\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12794\
        );

    \I__2294\ : InMux
    port map (
            O => \N__12826\,
            I => \N__12794\
        );

    \I__2293\ : InMux
    port map (
            O => \N__12823\,
            I => \N__12790\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__12820\,
            I => \N__12787\
        );

    \I__2291\ : InMux
    port map (
            O => \N__12819\,
            I => \N__12784\
        );

    \I__2290\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12781\
        );

    \I__2289\ : InMux
    port map (
            O => \N__12817\,
            I => \N__12778\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__12816\,
            I => \N__12770\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__12813\,
            I => \N__12766\
        );

    \I__2286\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12763\
        );

    \I__2285\ : InMux
    port map (
            O => \N__12811\,
            I => \N__12760\
        );

    \I__2284\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12749\
        );

    \I__2283\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12749\
        );

    \I__2282\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12749\
        );

    \I__2281\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12749\
        );

    \I__2280\ : InMux
    port map (
            O => \N__12806\,
            I => \N__12749\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__12803\,
            I => \N__12746\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__12794\,
            I => \N__12743\
        );

    \I__2277\ : InMux
    port map (
            O => \N__12793\,
            I => \N__12740\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__12790\,
            I => \N__12729\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__12787\,
            I => \N__12729\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__12784\,
            I => \N__12729\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__12781\,
            I => \N__12729\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__12778\,
            I => \N__12729\
        );

    \I__2271\ : InMux
    port map (
            O => \N__12777\,
            I => \N__12725\
        );

    \I__2270\ : InMux
    port map (
            O => \N__12776\,
            I => \N__12720\
        );

    \I__2269\ : InMux
    port map (
            O => \N__12775\,
            I => \N__12720\
        );

    \I__2268\ : InMux
    port map (
            O => \N__12774\,
            I => \N__12711\
        );

    \I__2267\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12711\
        );

    \I__2266\ : InMux
    port map (
            O => \N__12770\,
            I => \N__12711\
        );

    \I__2265\ : InMux
    port map (
            O => \N__12769\,
            I => \N__12711\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__12766\,
            I => \N__12701\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__12763\,
            I => \N__12701\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__12760\,
            I => \N__12701\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__12749\,
            I => \N__12701\
        );

    \I__2260\ : Span4Mux_v
    port map (
            O => \N__12746\,
            I => \N__12692\
        );

    \I__2259\ : Span4Mux_v
    port map (
            O => \N__12743\,
            I => \N__12692\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__12740\,
            I => \N__12692\
        );

    \I__2257\ : Span4Mux_v
    port map (
            O => \N__12729\,
            I => \N__12692\
        );

    \I__2256\ : InMux
    port map (
            O => \N__12728\,
            I => \N__12689\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__12725\,
            I => \N__12682\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__12720\,
            I => \N__12682\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__12711\,
            I => \N__12682\
        );

    \I__2252\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12677\
        );

    \I__2251\ : Span4Mux_v
    port map (
            O => \N__12701\,
            I => \N__12674\
        );

    \I__2250\ : Span4Mux_h
    port map (
            O => \N__12692\,
            I => \N__12671\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__12689\,
            I => \N__12666\
        );

    \I__2248\ : Span4Mux_h
    port map (
            O => \N__12682\,
            I => \N__12666\
        );

    \I__2247\ : InMux
    port map (
            O => \N__12681\,
            I => \N__12661\
        );

    \I__2246\ : InMux
    port map (
            O => \N__12680\,
            I => \N__12661\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__12677\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__12674\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__12671\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__12666\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__12661\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2240\ : InMux
    port map (
            O => \N__12650\,
            I => \N__12636\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__12649\,
            I => \N__12632\
        );

    \I__2238\ : InMux
    port map (
            O => \N__12648\,
            I => \N__12629\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12647\,
            I => \N__12626\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__12646\,
            I => \N__12620\
        );

    \I__2235\ : InMux
    port map (
            O => \N__12645\,
            I => \N__12614\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__12644\,
            I => \N__12611\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__12643\,
            I => \N__12606\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__12642\,
            I => \N__12603\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__12641\,
            I => \N__12597\
        );

    \I__2230\ : CascadeMux
    port map (
            O => \N__12640\,
            I => \N__12592\
        );

    \I__2229\ : InMux
    port map (
            O => \N__12639\,
            I => \N__12587\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__12636\,
            I => \N__12584\
        );

    \I__2227\ : InMux
    port map (
            O => \N__12635\,
            I => \N__12579\
        );

    \I__2226\ : InMux
    port map (
            O => \N__12632\,
            I => \N__12579\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__12629\,
            I => \N__12576\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__12626\,
            I => \N__12573\
        );

    \I__2223\ : InMux
    port map (
            O => \N__12625\,
            I => \N__12570\
        );

    \I__2222\ : InMux
    port map (
            O => \N__12624\,
            I => \N__12567\
        );

    \I__2221\ : InMux
    port map (
            O => \N__12623\,
            I => \N__12564\
        );

    \I__2220\ : InMux
    port map (
            O => \N__12620\,
            I => \N__12559\
        );

    \I__2219\ : InMux
    port map (
            O => \N__12619\,
            I => \N__12559\
        );

    \I__2218\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12554\
        );

    \I__2217\ : InMux
    port map (
            O => \N__12617\,
            I => \N__12554\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__12614\,
            I => \N__12551\
        );

    \I__2215\ : InMux
    port map (
            O => \N__12611\,
            I => \N__12546\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12610\,
            I => \N__12546\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__12609\,
            I => \N__12542\
        );

    \I__2212\ : InMux
    port map (
            O => \N__12606\,
            I => \N__12535\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12603\,
            I => \N__12535\
        );

    \I__2210\ : InMux
    port map (
            O => \N__12602\,
            I => \N__12535\
        );

    \I__2209\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12532\
        );

    \I__2208\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12528\
        );

    \I__2207\ : InMux
    port map (
            O => \N__12597\,
            I => \N__12525\
        );

    \I__2206\ : InMux
    port map (
            O => \N__12596\,
            I => \N__12516\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12516\
        );

    \I__2204\ : InMux
    port map (
            O => \N__12592\,
            I => \N__12516\
        );

    \I__2203\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12516\
        );

    \I__2202\ : InMux
    port map (
            O => \N__12590\,
            I => \N__12513\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__12587\,
            I => \N__12510\
        );

    \I__2200\ : Span4Mux_v
    port map (
            O => \N__12584\,
            I => \N__12505\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__12579\,
            I => \N__12505\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__12576\,
            I => \N__12498\
        );

    \I__2197\ : Span4Mux_v
    port map (
            O => \N__12573\,
            I => \N__12498\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__12570\,
            I => \N__12483\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__12567\,
            I => \N__12483\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__12564\,
            I => \N__12483\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__12559\,
            I => \N__12483\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__12554\,
            I => \N__12483\
        );

    \I__2191\ : Span4Mux_v
    port map (
            O => \N__12551\,
            I => \N__12483\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__12546\,
            I => \N__12483\
        );

    \I__2189\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12480\
        );

    \I__2188\ : InMux
    port map (
            O => \N__12542\,
            I => \N__12477\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__12535\,
            I => \N__12472\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__12532\,
            I => \N__12472\
        );

    \I__2185\ : InMux
    port map (
            O => \N__12531\,
            I => \N__12469\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__12528\,
            I => \N__12460\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__12525\,
            I => \N__12460\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__12516\,
            I => \N__12460\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__12513\,
            I => \N__12460\
        );

    \I__2180\ : Span4Mux_h
    port map (
            O => \N__12510\,
            I => \N__12455\
        );

    \I__2179\ : Span4Mux_v
    port map (
            O => \N__12505\,
            I => \N__12455\
        );

    \I__2178\ : InMux
    port map (
            O => \N__12504\,
            I => \N__12450\
        );

    \I__2177\ : InMux
    port map (
            O => \N__12503\,
            I => \N__12450\
        );

    \I__2176\ : Span4Mux_h
    port map (
            O => \N__12498\,
            I => \N__12445\
        );

    \I__2175\ : Span4Mux_v
    port map (
            O => \N__12483\,
            I => \N__12445\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__12480\,
            I => \N__12438\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__12477\,
            I => \N__12438\
        );

    \I__2172\ : Span4Mux_v
    port map (
            O => \N__12472\,
            I => \N__12438\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__12469\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2170\ : Odrv12
    port map (
            O => \N__12460\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__12455\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__12450\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__12445\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__12438\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__12425\,
            I => \N__12422\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12422\,
            I => \N__12415\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__12421\,
            I => \N__12410\
        );

    \I__2162\ : InMux
    port map (
            O => \N__12420\,
            I => \N__12405\
        );

    \I__2161\ : InMux
    port map (
            O => \N__12419\,
            I => \N__12402\
        );

    \I__2160\ : InMux
    port map (
            O => \N__12418\,
            I => \N__12396\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__12415\,
            I => \N__12393\
        );

    \I__2158\ : InMux
    port map (
            O => \N__12414\,
            I => \N__12390\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12413\,
            I => \N__12387\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12380\
        );

    \I__2155\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12380\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__12408\,
            I => \N__12376\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__12405\,
            I => \N__12373\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__12402\,
            I => \N__12370\
        );

    \I__2151\ : InMux
    port map (
            O => \N__12401\,
            I => \N__12363\
        );

    \I__2150\ : InMux
    port map (
            O => \N__12400\,
            I => \N__12363\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12399\,
            I => \N__12363\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__12396\,
            I => \N__12358\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__12393\,
            I => \N__12351\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__12390\,
            I => \N__12351\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__12387\,
            I => \N__12351\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12386\,
            I => \N__12346\
        );

    \I__2143\ : InMux
    port map (
            O => \N__12385\,
            I => \N__12346\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__12380\,
            I => \N__12343\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__12379\,
            I => \N__12335\
        );

    \I__2140\ : InMux
    port map (
            O => \N__12376\,
            I => \N__12331\
        );

    \I__2139\ : Span4Mux_v
    port map (
            O => \N__12373\,
            I => \N__12326\
        );

    \I__2138\ : Span4Mux_v
    port map (
            O => \N__12370\,
            I => \N__12326\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__12363\,
            I => \N__12323\
        );

    \I__2136\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12318\
        );

    \I__2135\ : InMux
    port map (
            O => \N__12361\,
            I => \N__12318\
        );

    \I__2134\ : Span4Mux_h
    port map (
            O => \N__12358\,
            I => \N__12309\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__12351\,
            I => \N__12309\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__12346\,
            I => \N__12309\
        );

    \I__2131\ : Span4Mux_h
    port map (
            O => \N__12343\,
            I => \N__12309\
        );

    \I__2130\ : InMux
    port map (
            O => \N__12342\,
            I => \N__12298\
        );

    \I__2129\ : InMux
    port map (
            O => \N__12341\,
            I => \N__12298\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12340\,
            I => \N__12298\
        );

    \I__2127\ : InMux
    port map (
            O => \N__12339\,
            I => \N__12298\
        );

    \I__2126\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12298\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12335\,
            I => \N__12293\
        );

    \I__2124\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12293\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__12331\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__12326\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2121\ : Odrv12
    port map (
            O => \N__12323\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__12318\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__12309\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__12298\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__12293\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2116\ : InMux
    port map (
            O => \N__12278\,
            I => \N__12274\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__12277\,
            I => \N__12271\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__12274\,
            I => \N__12268\
        );

    \I__2113\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12265\
        );

    \I__2112\ : Span4Mux_h
    port map (
            O => \N__12268\,
            I => \N__12262\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__12265\,
            I => \this_vga_signals.M_vcounter_d7lt8_0\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__12262\,
            I => \this_vga_signals.M_vcounter_d7lt8_0\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__12257\,
            I => \N__12250\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__12256\,
            I => \N__12243\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__12255\,
            I => \N__12239\
        );

    \I__2106\ : InMux
    port map (
            O => \N__12254\,
            I => \N__12236\
        );

    \I__2105\ : InMux
    port map (
            O => \N__12253\,
            I => \N__12231\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12250\,
            I => \N__12231\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__12249\,
            I => \N__12228\
        );

    \I__2102\ : InMux
    port map (
            O => \N__12248\,
            I => \N__12225\
        );

    \I__2101\ : InMux
    port map (
            O => \N__12247\,
            I => \N__12220\
        );

    \I__2100\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12220\
        );

    \I__2099\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12215\
        );

    \I__2098\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12212\
        );

    \I__2097\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12206\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__12236\,
            I => \N__12203\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__12231\,
            I => \N__12200\
        );

    \I__2094\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12197\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__12225\,
            I => \N__12192\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__12220\,
            I => \N__12192\
        );

    \I__2091\ : InMux
    port map (
            O => \N__12219\,
            I => \N__12187\
        );

    \I__2090\ : InMux
    port map (
            O => \N__12218\,
            I => \N__12187\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__12215\,
            I => \N__12180\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__12212\,
            I => \N__12177\
        );

    \I__2087\ : InMux
    port map (
            O => \N__12211\,
            I => \N__12174\
        );

    \I__2086\ : InMux
    port map (
            O => \N__12210\,
            I => \N__12169\
        );

    \I__2085\ : InMux
    port map (
            O => \N__12209\,
            I => \N__12169\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__12206\,
            I => \N__12164\
        );

    \I__2083\ : Span4Mux_v
    port map (
            O => \N__12203\,
            I => \N__12164\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__12200\,
            I => \N__12157\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__12197\,
            I => \N__12157\
        );

    \I__2080\ : Span4Mux_v
    port map (
            O => \N__12192\,
            I => \N__12157\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__12187\,
            I => \N__12154\
        );

    \I__2078\ : InMux
    port map (
            O => \N__12186\,
            I => \N__12149\
        );

    \I__2077\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12149\
        );

    \I__2076\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12144\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12183\,
            I => \N__12144\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__12180\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__12177\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__12174\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__12169\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__12164\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__12157\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__12154\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__12149\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__12144\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__12125\,
            I => \this_vga_signals.un4_lvisibility_1_cascade_\
        );

    \I__2064\ : InMux
    port map (
            O => \N__12122\,
            I => \N__12119\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__12119\,
            I => \N__12113\
        );

    \I__2062\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12107\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__12117\,
            I => \N__12104\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__12116\,
            I => \N__12101\
        );

    \I__2059\ : Span4Mux_v
    port map (
            O => \N__12113\,
            I => \N__12098\
        );

    \I__2058\ : InMux
    port map (
            O => \N__12112\,
            I => \N__12095\
        );

    \I__2057\ : InMux
    port map (
            O => \N__12111\,
            I => \N__12090\
        );

    \I__2056\ : InMux
    port map (
            O => \N__12110\,
            I => \N__12090\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__12107\,
            I => \N__12087\
        );

    \I__2054\ : InMux
    port map (
            O => \N__12104\,
            I => \N__12084\
        );

    \I__2053\ : InMux
    port map (
            O => \N__12101\,
            I => \N__12081\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__12098\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__12095\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__12090\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__12087\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__12084\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__12081\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2046\ : InMux
    port map (
            O => \N__12068\,
            I => \N__12062\
        );

    \I__2045\ : InMux
    port map (
            O => \N__12067\,
            I => \N__12062\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__12062\,
            I => \this_vga_signals.line_clk_1\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__12059\,
            I => \N__12056\
        );

    \I__2042\ : InMux
    port map (
            O => \N__12056\,
            I => \N__12053\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__12053\,
            I => \this_vga_signals.un4_lvisibility_1\
        );

    \I__2040\ : InMux
    port map (
            O => \N__12050\,
            I => \N__12043\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12040\
        );

    \I__2038\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12035\
        );

    \I__2037\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12032\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12046\,
            I => \N__12029\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__12043\,
            I => \N__12024\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__12040\,
            I => \N__12024\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12020\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__12038\,
            I => \N__12016\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__12035\,
            I => \N__12013\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__12032\,
            I => \N__12010\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__12029\,
            I => \N__12005\
        );

    \I__2028\ : Span4Mux_v
    port map (
            O => \N__12024\,
            I => \N__12005\
        );

    \I__2027\ : InMux
    port map (
            O => \N__12023\,
            I => \N__12002\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__12020\,
            I => \N__11999\
        );

    \I__2025\ : InMux
    port map (
            O => \N__12019\,
            I => \N__11994\
        );

    \I__2024\ : InMux
    port map (
            O => \N__12016\,
            I => \N__11994\
        );

    \I__2023\ : Span4Mux_h
    port map (
            O => \N__12013\,
            I => \N__11991\
        );

    \I__2022\ : Odrv12
    port map (
            O => \N__12010\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__12005\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__12002\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__11999\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__11994\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__11991\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__11978\,
            I => \N__11974\
        );

    \I__2015\ : InMux
    port map (
            O => \N__11977\,
            I => \N__11971\
        );

    \I__2014\ : InMux
    port map (
            O => \N__11974\,
            I => \N__11968\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__11971\,
            I => \N__11965\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__11968\,
            I => \N__11960\
        );

    \I__2011\ : Span4Mux_h
    port map (
            O => \N__11965\,
            I => \N__11957\
        );

    \I__2010\ : InMux
    port map (
            O => \N__11964\,
            I => \N__11954\
        );

    \I__2009\ : InMux
    port map (
            O => \N__11963\,
            I => \N__11951\
        );

    \I__2008\ : Span4Mux_h
    port map (
            O => \N__11960\,
            I => \N__11946\
        );

    \I__2007\ : Span4Mux_h
    port map (
            O => \N__11957\,
            I => \N__11946\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__11954\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__11951\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__11946\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__11939\,
            I => \N__11932\
        );

    \I__2002\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11927\
        );

    \I__2001\ : InMux
    port map (
            O => \N__11937\,
            I => \N__11924\
        );

    \I__2000\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11919\
        );

    \I__1999\ : InMux
    port map (
            O => \N__11935\,
            I => \N__11919\
        );

    \I__1998\ : InMux
    port map (
            O => \N__11932\,
            I => \N__11914\
        );

    \I__1997\ : InMux
    port map (
            O => \N__11931\,
            I => \N__11914\
        );

    \I__1996\ : InMux
    port map (
            O => \N__11930\,
            I => \N__11911\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__11927\,
            I => \N__11906\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__11924\,
            I => \N__11906\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__11919\,
            I => \N__11901\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__11914\,
            I => \N__11901\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__11911\,
            I => \N__11897\
        );

    \I__1990\ : Span4Mux_v
    port map (
            O => \N__11906\,
            I => \N__11894\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__11901\,
            I => \N__11891\
        );

    \I__1988\ : InMux
    port map (
            O => \N__11900\,
            I => \N__11888\
        );

    \I__1987\ : Span4Mux_v
    port map (
            O => \N__11897\,
            I => \N__11881\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__11894\,
            I => \N__11881\
        );

    \I__1985\ : Span4Mux_h
    port map (
            O => \N__11891\,
            I => \N__11881\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__11888\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__11881\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1982\ : InMux
    port map (
            O => \N__11876\,
            I => \N__11873\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__11873\,
            I => \N__11870\
        );

    \I__1980\ : Span4Mux_h
    port map (
            O => \N__11870\,
            I => \N__11867\
        );

    \I__1979\ : Span4Mux_h
    port map (
            O => \N__11867\,
            I => \N__11864\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__11864\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__1977\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11858\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__11858\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__1975\ : InMux
    port map (
            O => \N__11855\,
            I => \N__11846\
        );

    \I__1974\ : InMux
    port map (
            O => \N__11854\,
            I => \N__11846\
        );

    \I__1973\ : InMux
    port map (
            O => \N__11853\,
            I => \N__11846\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__11846\,
            I => \M_this_delay_clk_out_0\
        );

    \I__1971\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11834\
        );

    \I__1970\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11834\
        );

    \I__1969\ : InMux
    port map (
            O => \N__11841\,
            I => \N__11834\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__11834\,
            I => \N__11831\
        );

    \I__1967\ : Sp12to4
    port map (
            O => \N__11831\,
            I => \N__11828\
        );

    \I__1966\ : Span12Mux_v
    port map (
            O => \N__11828\,
            I => \N__11825\
        );

    \I__1965\ : Span12Mux_h
    port map (
            O => \N__11825\,
            I => \N__11822\
        );

    \I__1964\ : Odrv12
    port map (
            O => \N__11822\,
            I => port_enb_c
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__11819\,
            I => \N__11816\
        );

    \I__1962\ : InMux
    port map (
            O => \N__11816\,
            I => \N__11810\
        );

    \I__1961\ : InMux
    port map (
            O => \N__11815\,
            I => \N__11810\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__11810\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__1959\ : InMux
    port map (
            O => \N__11807\,
            I => \N__11803\
        );

    \I__1958\ : InMux
    port map (
            O => \N__11806\,
            I => \N__11800\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__11803\,
            I => \N__11797\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__11800\,
            I => \N__11794\
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__11797\,
            I => \this_vga_signals.vaddress_ac0_9_0_a0_0\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__11794\,
            I => \this_vga_signals.vaddress_ac0_9_0_a0_0\
        );

    \I__1953\ : InMux
    port map (
            O => \N__11789\,
            I => \N__11786\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__11786\,
            I => \N__11783\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__11783\,
            I => \this_vga_signals.un6_vvisibilitylt9_0\
        );

    \I__1950\ : InMux
    port map (
            O => \N__11780\,
            I => \N__11777\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__11777\,
            I => \N__11773\
        );

    \I__1948\ : InMux
    port map (
            O => \N__11776\,
            I => \N__11770\
        );

    \I__1947\ : Span4Mux_h
    port map (
            O => \N__11773\,
            I => \N__11764\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__11770\,
            I => \N__11764\
        );

    \I__1945\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11761\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__11764\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__11761\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__1942\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11753\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__11753\,
            I => \N__11749\
        );

    \I__1940\ : InMux
    port map (
            O => \N__11752\,
            I => \N__11745\
        );

    \I__1939\ : Span4Mux_h
    port map (
            O => \N__11749\,
            I => \N__11742\
        );

    \I__1938\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11739\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__11745\,
            I => \N__11736\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__11742\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__11739\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1934\ : Odrv12
    port map (
            O => \N__11736\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1933\ : InMux
    port map (
            O => \N__11729\,
            I => \N__11724\
        );

    \I__1932\ : InMux
    port map (
            O => \N__11728\,
            I => \N__11721\
        );

    \I__1931\ : InMux
    port map (
            O => \N__11727\,
            I => \N__11718\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__11724\,
            I => \N__11715\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__11721\,
            I => \N__11712\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__11718\,
            I => \N__11709\
        );

    \I__1927\ : Span4Mux_h
    port map (
            O => \N__11715\,
            I => \N__11706\
        );

    \I__1926\ : Span4Mux_h
    port map (
            O => \N__11712\,
            I => \N__11703\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__11709\,
            I => \N__11700\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__11706\,
            I => \this_vga_signals.vaddress_5_6\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__11703\,
            I => \this_vga_signals.vaddress_5_6\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__11700\,
            I => \this_vga_signals.vaddress_5_6\
        );

    \I__1921\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11690\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__11690\,
            I => \N__11685\
        );

    \I__1919\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11682\
        );

    \I__1918\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11678\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__11685\,
            I => \N__11675\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__11682\,
            I => \N__11672\
        );

    \I__1915\ : InMux
    port map (
            O => \N__11681\,
            I => \N__11669\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__11678\,
            I => \N__11666\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__11675\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1912\ : Odrv12
    port map (
            O => \N__11672\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__11669\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__11666\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__11657\,
            I => \N__11653\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11650\
        );

    \I__1907\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11647\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__11650\,
            I => \N__11644\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__11647\,
            I => \N__11641\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__11644\,
            I => \N__11638\
        );

    \I__1903\ : Span4Mux_h
    port map (
            O => \N__11641\,
            I => \N__11635\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__11638\,
            I => \this_vga_signals.vaddress_3_5\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__11635\,
            I => \this_vga_signals.vaddress_3_5\
        );

    \I__1900\ : InMux
    port map (
            O => \N__11630\,
            I => \N__11627\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__11627\,
            I => \N__11623\
        );

    \I__1898\ : InMux
    port map (
            O => \N__11626\,
            I => \N__11620\
        );

    \I__1897\ : Span4Mux_h
    port map (
            O => \N__11623\,
            I => \N__11615\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__11620\,
            I => \N__11615\
        );

    \I__1895\ : Span4Mux_v
    port map (
            O => \N__11615\,
            I => \N__11611\
        );

    \I__1894\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11608\
        );

    \I__1893\ : Span4Mux_h
    port map (
            O => \N__11611\,
            I => \N__11605\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__11608\,
            I => \N__11602\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__11605\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__11602\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__1889\ : CEMux
    port map (
            O => \N__11597\,
            I => \N__11573\
        );

    \I__1888\ : CEMux
    port map (
            O => \N__11596\,
            I => \N__11573\
        );

    \I__1887\ : CEMux
    port map (
            O => \N__11595\,
            I => \N__11573\
        );

    \I__1886\ : CEMux
    port map (
            O => \N__11594\,
            I => \N__11573\
        );

    \I__1885\ : CEMux
    port map (
            O => \N__11593\,
            I => \N__11573\
        );

    \I__1884\ : CEMux
    port map (
            O => \N__11592\,
            I => \N__11573\
        );

    \I__1883\ : CEMux
    port map (
            O => \N__11591\,
            I => \N__11573\
        );

    \I__1882\ : CEMux
    port map (
            O => \N__11590\,
            I => \N__11573\
        );

    \I__1881\ : GlobalMux
    port map (
            O => \N__11573\,
            I => \N__11570\
        );

    \I__1880\ : gio2CtrlBuf
    port map (
            O => \N__11570\,
            I => \this_vga_signals.N_340_0_g\
        );

    \I__1879\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11564\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__11564\,
            I => \N__11552\
        );

    \I__1877\ : SRMux
    port map (
            O => \N__11563\,
            I => \N__11531\
        );

    \I__1876\ : SRMux
    port map (
            O => \N__11562\,
            I => \N__11531\
        );

    \I__1875\ : SRMux
    port map (
            O => \N__11561\,
            I => \N__11531\
        );

    \I__1874\ : SRMux
    port map (
            O => \N__11560\,
            I => \N__11531\
        );

    \I__1873\ : SRMux
    port map (
            O => \N__11559\,
            I => \N__11531\
        );

    \I__1872\ : SRMux
    port map (
            O => \N__11558\,
            I => \N__11531\
        );

    \I__1871\ : SRMux
    port map (
            O => \N__11557\,
            I => \N__11531\
        );

    \I__1870\ : SRMux
    port map (
            O => \N__11556\,
            I => \N__11531\
        );

    \I__1869\ : SRMux
    port map (
            O => \N__11555\,
            I => \N__11531\
        );

    \I__1868\ : Glb2LocalMux
    port map (
            O => \N__11552\,
            I => \N__11531\
        );

    \I__1867\ : GlobalMux
    port map (
            O => \N__11531\,
            I => \N__11528\
        );

    \I__1866\ : gio2CtrlBuf
    port map (
            O => \N__11528\,
            I => \this_vga_signals.N_515_g\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__11525\,
            I => \N__11522\
        );

    \I__1864\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11516\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11521\,
            I => \N__11513\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__11520\,
            I => \N__11509\
        );

    \I__1861\ : InMux
    port map (
            O => \N__11519\,
            I => \N__11505\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__11516\,
            I => \N__11500\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__11513\,
            I => \N__11500\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11512\,
            I => \N__11497\
        );

    \I__1857\ : InMux
    port map (
            O => \N__11509\,
            I => \N__11492\
        );

    \I__1856\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11492\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__11505\,
            I => \N__11481\
        );

    \I__1854\ : Span4Mux_h
    port map (
            O => \N__11500\,
            I => \N__11481\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__11497\,
            I => \N__11476\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__11492\,
            I => \N__11476\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11469\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11490\,
            I => \N__11469\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11469\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11462\
        );

    \I__1847\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11462\
        );

    \I__1846\ : InMux
    port map (
            O => \N__11486\,
            I => \N__11462\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__11481\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1844\ : Odrv12
    port map (
            O => \N__11476\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__11469\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__11462\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1841\ : InMux
    port map (
            O => \N__11453\,
            I => \N__11445\
        );

    \I__1840\ : InMux
    port map (
            O => \N__11452\,
            I => \N__11442\
        );

    \I__1839\ : InMux
    port map (
            O => \N__11451\,
            I => \N__11433\
        );

    \I__1838\ : InMux
    port map (
            O => \N__11450\,
            I => \N__11433\
        );

    \I__1837\ : InMux
    port map (
            O => \N__11449\,
            I => \N__11433\
        );

    \I__1836\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11433\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__11445\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__11442\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__11433\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1832\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11419\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11416\
        );

    \I__1830\ : InMux
    port map (
            O => \N__11424\,
            I => \N__11409\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11423\,
            I => \N__11409\
        );

    \I__1828\ : InMux
    port map (
            O => \N__11422\,
            I => \N__11409\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__11419\,
            I => \N__11406\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__11416\,
            I => \N__11401\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__11409\,
            I => \N__11401\
        );

    \I__1824\ : Span4Mux_h
    port map (
            O => \N__11406\,
            I => \N__11398\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__11401\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__11398\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__11393\,
            I => \N__11384\
        );

    \I__1820\ : InMux
    port map (
            O => \N__11392\,
            I => \N__11381\
        );

    \I__1819\ : InMux
    port map (
            O => \N__11391\,
            I => \N__11372\
        );

    \I__1818\ : InMux
    port map (
            O => \N__11390\,
            I => \N__11372\
        );

    \I__1817\ : InMux
    port map (
            O => \N__11389\,
            I => \N__11372\
        );

    \I__1816\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11367\
        );

    \I__1815\ : InMux
    port map (
            O => \N__11387\,
            I => \N__11367\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11384\,
            I => \N__11364\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__11381\,
            I => \N__11361\
        );

    \I__1812\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11353\
        );

    \I__1811\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11350\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__11372\,
            I => \N__11343\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__11367\,
            I => \N__11343\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__11364\,
            I => \N__11343\
        );

    \I__1807\ : Span4Mux_v
    port map (
            O => \N__11361\,
            I => \N__11335\
        );

    \I__1806\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11332\
        );

    \I__1805\ : InMux
    port map (
            O => \N__11359\,
            I => \N__11323\
        );

    \I__1804\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11323\
        );

    \I__1803\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11323\
        );

    \I__1802\ : InMux
    port map (
            O => \N__11356\,
            I => \N__11323\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__11353\,
            I => \N__11320\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__11350\,
            I => \N__11315\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__11343\,
            I => \N__11315\
        );

    \I__1798\ : InMux
    port map (
            O => \N__11342\,
            I => \N__11310\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11341\,
            I => \N__11310\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11340\,
            I => \N__11303\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11339\,
            I => \N__11303\
        );

    \I__1794\ : InMux
    port map (
            O => \N__11338\,
            I => \N__11303\
        );

    \I__1793\ : Odrv4
    port map (
            O => \N__11335\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__11332\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__11323\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__11320\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__11315\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__11310\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__11303\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z2\
        );

    \I__1786\ : InMux
    port map (
            O => \N__11288\,
            I => \N__11285\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__11285\,
            I => \this_vga_signals.vaddress_4_6\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__11282\,
            I => \this_vga_signals.M_vcounter_d7lto8_1_cascade_\
        );

    \I__1783\ : InMux
    port map (
            O => \N__11279\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__1782\ : InMux
    port map (
            O => \N__11276\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__1781\ : InMux
    port map (
            O => \N__11273\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__1780\ : InMux
    port map (
            O => \N__11270\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__1779\ : InMux
    port map (
            O => \N__11267\,
            I => \N__11261\
        );

    \I__1778\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11261\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__11261\,
            I => \N__11257\
        );

    \I__1776\ : InMux
    port map (
            O => \N__11260\,
            I => \N__11254\
        );

    \I__1775\ : Span4Mux_h
    port map (
            O => \N__11257\,
            I => \N__11251\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__11254\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__11251\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11246\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11243\,
            I => \bfn_13_18_0_\
        );

    \I__1770\ : InMux
    port map (
            O => \N__11240\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11237\,
            I => \N__11234\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__11234\,
            I => \N__11229\
        );

    \I__1767\ : InMux
    port map (
            O => \N__11233\,
            I => \N__11226\
        );

    \I__1766\ : InMux
    port map (
            O => \N__11232\,
            I => \N__11223\
        );

    \I__1765\ : Odrv12
    port map (
            O => \N__11229\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__11226\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__11223\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11213\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__11213\,
            I => \this_vga_signals.vsync_1_3\
        );

    \I__1760\ : IoInMux
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__11207\,
            I => \N__11204\
        );

    \I__1758\ : Span4Mux_s2_v
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__1757\ : Sp12to4
    port map (
            O => \N__11201\,
            I => \N__11198\
        );

    \I__1756\ : Span12Mux_s11_h
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__1755\ : Odrv12
    port map (
            O => \N__11195\,
            I => this_vga_signals_vsync_1_i
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__11192\,
            I => \N__11188\
        );

    \I__1753\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11183\
        );

    \I__1752\ : InMux
    port map (
            O => \N__11188\,
            I => \N__11179\
        );

    \I__1751\ : InMux
    port map (
            O => \N__11187\,
            I => \N__11176\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__11186\,
            I => \N__11170\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__11183\,
            I => \N__11166\
        );

    \I__1748\ : InMux
    port map (
            O => \N__11182\,
            I => \N__11163\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__11179\,
            I => \N__11158\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__11176\,
            I => \N__11158\
        );

    \I__1745\ : InMux
    port map (
            O => \N__11175\,
            I => \N__11155\
        );

    \I__1744\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11152\
        );

    \I__1743\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11145\
        );

    \I__1742\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11145\
        );

    \I__1741\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11145\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__11166\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__11163\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1738\ : Odrv12
    port map (
            O => \N__11158\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__11155\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11152\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__11145\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__11132\,
            I => \N__11124\
        );

    \I__1733\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11115\
        );

    \I__1732\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11115\
        );

    \I__1731\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11112\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__11128\,
            I => \N__11108\
        );

    \I__1729\ : InMux
    port map (
            O => \N__11127\,
            I => \N__11103\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11124\,
            I => \N__11100\
        );

    \I__1727\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11095\
        );

    \I__1726\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11095\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11092\
        );

    \I__1724\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11089\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__11115\,
            I => \N__11084\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__11112\,
            I => \N__11084\
        );

    \I__1721\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11075\
        );

    \I__1720\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11075\
        );

    \I__1719\ : InMux
    port map (
            O => \N__11107\,
            I => \N__11075\
        );

    \I__1718\ : InMux
    port map (
            O => \N__11106\,
            I => \N__11075\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__11103\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__11100\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__11095\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__11092\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__11089\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__11084\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__11075\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1710\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11052\
        );

    \I__1709\ : CascadeMux
    port map (
            O => \N__11059\,
            I => \N__11049\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__11058\,
            I => \N__11044\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__11057\,
            I => \N__11041\
        );

    \I__1706\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11038\
        );

    \I__1705\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11035\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__11052\,
            I => \N__11032\
        );

    \I__1703\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11029\
        );

    \I__1702\ : InMux
    port map (
            O => \N__11048\,
            I => \N__11023\
        );

    \I__1701\ : InMux
    port map (
            O => \N__11047\,
            I => \N__11020\
        );

    \I__1700\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11015\
        );

    \I__1699\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11015\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__11038\,
            I => \N__11006\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__11035\,
            I => \N__11006\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__11032\,
            I => \N__11006\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__11029\,
            I => \N__11006\
        );

    \I__1694\ : InMux
    port map (
            O => \N__11028\,
            I => \N__10999\
        );

    \I__1693\ : InMux
    port map (
            O => \N__11027\,
            I => \N__10999\
        );

    \I__1692\ : InMux
    port map (
            O => \N__11026\,
            I => \N__10999\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__11023\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__11020\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__11015\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__11006\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__10999\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1686\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10984\
        );

    \I__1685\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10978\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__10984\,
            I => \N__10975\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__10983\,
            I => \N__10968\
        );

    \I__1682\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10965\
        );

    \I__1681\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10962\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__10978\,
            I => \N__10957\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__10975\,
            I => \N__10957\
        );

    \I__1678\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10954\
        );

    \I__1677\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10951\
        );

    \I__1676\ : InMux
    port map (
            O => \N__10972\,
            I => \N__10944\
        );

    \I__1675\ : InMux
    port map (
            O => \N__10971\,
            I => \N__10944\
        );

    \I__1674\ : InMux
    port map (
            O => \N__10968\,
            I => \N__10944\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__10965\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__10962\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__10957\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__10954\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__10951\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__10944\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__10931\,
            I => \this_vga_signals.M_hcounter_d7lto7_0_cascade_\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__10928\,
            I => \N__10924\
        );

    \I__1665\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10920\
        );

    \I__1664\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10916\
        );

    \I__1663\ : InMux
    port map (
            O => \N__10923\,
            I => \N__10913\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__10920\,
            I => \N__10910\
        );

    \I__1661\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10902\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__10916\,
            I => \N__10895\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__10913\,
            I => \N__10895\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__10910\,
            I => \N__10895\
        );

    \I__1657\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10892\
        );

    \I__1656\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10889\
        );

    \I__1655\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10882\
        );

    \I__1654\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10882\
        );

    \I__1653\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10882\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__10902\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__10895\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__10892\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__10889\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__10882\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1647\ : InMux
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__10868\,
            I => \this_vga_signals.un2_vsynclt8\
        );

    \I__1645\ : CEMux
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__10862\,
            I => \this_vga_signals.N_340_1\
        );

    \I__1643\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10856\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__10856\,
            I => \this_vga_signals.vsync_1_2\
        );

    \I__1641\ : InMux
    port map (
            O => \N__10853\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__1640\ : InMux
    port map (
            O => \N__10850\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__1639\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__10844\,
            I => \this_vga_signals.g2_1\
        );

    \I__1637\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10838\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__10838\,
            I => \N__10834\
        );

    \I__1635\ : InMux
    port map (
            O => \N__10837\,
            I => \N__10831\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__10834\,
            I => \this_vga_signals.if_N_5\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__10831\,
            I => \this_vga_signals.if_N_5\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__10826\,
            I => \N__10823\
        );

    \I__1631\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10820\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__10820\,
            I => \this_vga_signals.vaddress_4_5\
        );

    \I__1629\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10814\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__10814\,
            I => \this_vga_signals.vaddress_3_6\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__10811\,
            I => \N__10802\
        );

    \I__1626\ : InMux
    port map (
            O => \N__10810\,
            I => \N__10796\
        );

    \I__1625\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10796\
        );

    \I__1624\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10793\
        );

    \I__1623\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10784\
        );

    \I__1622\ : InMux
    port map (
            O => \N__10806\,
            I => \N__10784\
        );

    \I__1621\ : InMux
    port map (
            O => \N__10805\,
            I => \N__10780\
        );

    \I__1620\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10774\
        );

    \I__1619\ : InMux
    port map (
            O => \N__10801\,
            I => \N__10774\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__10796\,
            I => \N__10768\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__10793\,
            I => \N__10768\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__10792\,
            I => \N__10761\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__10791\,
            I => \N__10757\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__10790\,
            I => \N__10752\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__10789\,
            I => \N__10749\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__10784\,
            I => \N__10746\
        );

    \I__1611\ : InMux
    port map (
            O => \N__10783\,
            I => \N__10743\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__10780\,
            I => \N__10740\
        );

    \I__1609\ : InMux
    port map (
            O => \N__10779\,
            I => \N__10737\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__10774\,
            I => \N__10734\
        );

    \I__1607\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10731\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__10768\,
            I => \N__10728\
        );

    \I__1605\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10715\
        );

    \I__1604\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10715\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10765\,
            I => \N__10715\
        );

    \I__1602\ : InMux
    port map (
            O => \N__10764\,
            I => \N__10715\
        );

    \I__1601\ : InMux
    port map (
            O => \N__10761\,
            I => \N__10715\
        );

    \I__1600\ : InMux
    port map (
            O => \N__10760\,
            I => \N__10715\
        );

    \I__1599\ : InMux
    port map (
            O => \N__10757\,
            I => \N__10704\
        );

    \I__1598\ : InMux
    port map (
            O => \N__10756\,
            I => \N__10704\
        );

    \I__1597\ : InMux
    port map (
            O => \N__10755\,
            I => \N__10704\
        );

    \I__1596\ : InMux
    port map (
            O => \N__10752\,
            I => \N__10704\
        );

    \I__1595\ : InMux
    port map (
            O => \N__10749\,
            I => \N__10704\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__10746\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__10743\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__10740\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__10737\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__10734\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__10731\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__10728\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__10715\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__10704\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__10685\,
            I => \this_vga_signals.vaddress_0_5_cascade_\
        );

    \I__1584\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10677\
        );

    \I__1583\ : InMux
    port map (
            O => \N__10681\,
            I => \N__10674\
        );

    \I__1582\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10666\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__10677\,
            I => \N__10663\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__10674\,
            I => \N__10660\
        );

    \I__1579\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10655\
        );

    \I__1578\ : InMux
    port map (
            O => \N__10672\,
            I => \N__10655\
        );

    \I__1577\ : InMux
    port map (
            O => \N__10671\,
            I => \N__10652\
        );

    \I__1576\ : InMux
    port map (
            O => \N__10670\,
            I => \N__10649\
        );

    \I__1575\ : InMux
    port map (
            O => \N__10669\,
            I => \N__10635\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__10666\,
            I => \N__10630\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__10663\,
            I => \N__10630\
        );

    \I__1572\ : Span4Mux_h
    port map (
            O => \N__10660\,
            I => \N__10627\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__10655\,
            I => \N__10624\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__10652\,
            I => \N__10621\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__10649\,
            I => \N__10618\
        );

    \I__1568\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10607\
        );

    \I__1567\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10607\
        );

    \I__1566\ : InMux
    port map (
            O => \N__10646\,
            I => \N__10607\
        );

    \I__1565\ : InMux
    port map (
            O => \N__10645\,
            I => \N__10607\
        );

    \I__1564\ : InMux
    port map (
            O => \N__10644\,
            I => \N__10607\
        );

    \I__1563\ : InMux
    port map (
            O => \N__10643\,
            I => \N__10594\
        );

    \I__1562\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10594\
        );

    \I__1561\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10594\
        );

    \I__1560\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10594\
        );

    \I__1559\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10594\
        );

    \I__1558\ : InMux
    port map (
            O => \N__10638\,
            I => \N__10594\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__10635\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1556\ : Odrv4
    port map (
            O => \N__10630\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1555\ : Odrv4
    port map (
            O => \N__10627\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__10624\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__10621\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1552\ : Odrv12
    port map (
            O => \N__10618\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__10607\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__10594\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__10577\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0_cascade_\
        );

    \I__1548\ : InMux
    port map (
            O => \N__10574\,
            I => \N__10571\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__10571\,
            I => \this_vga_signals.g2\
        );

    \I__1546\ : InMux
    port map (
            O => \N__10568\,
            I => \N__10565\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__10565\,
            I => \this_vga_signals.g1\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10558\
        );

    \I__1543\ : InMux
    port map (
            O => \N__10561\,
            I => \N__10555\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__10558\,
            I => \this_vga_signals.vaddress_0_6\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__10555\,
            I => \this_vga_signals.vaddress_0_6\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10547\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__10547\,
            I => \this_vga_signals.g1_0_2\
        );

    \I__1538\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__10541\,
            I => \this_vga_signals.g0_31_1\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__10538\,
            I => \N__10535\
        );

    \I__1535\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10532\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__10532\,
            I => \this_vga_signals.g1_0_1\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10525\
        );

    \I__1532\ : InMux
    port map (
            O => \N__10528\,
            I => \N__10519\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__10525\,
            I => \N__10516\
        );

    \I__1530\ : InMux
    port map (
            O => \N__10524\,
            I => \N__10513\
        );

    \I__1529\ : InMux
    port map (
            O => \N__10523\,
            I => \N__10508\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10522\,
            I => \N__10508\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__10519\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_N_2L1\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__10516\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_N_2L1\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__10513\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_N_2L1\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__10508\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_N_2L1\
        );

    \I__1523\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10496\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__10496\,
            I => \this_vga_signals.N_5_1_0_0\
        );

    \I__1521\ : InMux
    port map (
            O => \N__10493\,
            I => \N__10490\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__10490\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2_0_1_0\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__10487\,
            I => \this_vga_signals.g0_22_1_cascade_\
        );

    \I__1518\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10481\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__10481\,
            I => \N__10478\
        );

    \I__1516\ : Odrv12
    port map (
            O => \N__10478\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0_0_0_0\
        );

    \I__1515\ : InMux
    port map (
            O => \N__10475\,
            I => \N__10471\
        );

    \I__1514\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10468\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__10471\,
            I => \this_vga_signals.mult1_un61_sum_c3_0\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__10468\,
            I => \this_vga_signals.mult1_un61_sum_c3_0\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__10463\,
            I => \this_vga_signals.vaddress_5_5_cascade_\
        );

    \I__1510\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10457\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_1\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__10454\,
            I => \N__10446\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__10453\,
            I => \N__10443\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10440\
        );

    \I__1505\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10435\
        );

    \I__1504\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10435\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10449\,
            I => \N__10430\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10430\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10427\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__10440\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__10435\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__10430\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__10427\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__10418\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_1_cascade_\
        );

    \I__1495\ : InMux
    port map (
            O => \N__10415\,
            I => \N__10409\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10409\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__10409\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0_0\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10406\,
            I => \N__10403\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__10403\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_0_0_0\
        );

    \I__1490\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__10397\,
            I => \N__10394\
        );

    \I__1488\ : Span4Mux_h
    port map (
            O => \N__10394\,
            I => \N__10383\
        );

    \I__1487\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10380\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10392\,
            I => \N__10375\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10391\,
            I => \N__10375\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10372\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10367\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10388\,
            I => \N__10367\
        );

    \I__1481\ : InMux
    port map (
            O => \N__10387\,
            I => \N__10362\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10386\,
            I => \N__10362\
        );

    \I__1479\ : Odrv4
    port map (
            O => \N__10383\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__10380\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__10375\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__10372\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__10367\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__10362\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10346\,
            I => \N__10343\
        );

    \I__1471\ : Span4Mux_h
    port map (
            O => \N__10343\,
            I => \N__10339\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10342\,
            I => \N__10336\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__10339\,
            I => \this_vga_signals.vaddress_2_0_6\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__10336\,
            I => \this_vga_signals.vaddress_2_0_6\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__1466\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10325\,
            I => \this_vga_signals.g0_7_0\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__10322\,
            I => \N__10315\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__10321\,
            I => \N__10312\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10320\,
            I => \N__10309\
        );

    \I__1461\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10306\
        );

    \I__1460\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10303\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10315\,
            I => \N__10300\
        );

    \I__1458\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10297\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__10309\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__10306\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__10303\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__10300\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__10297\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10286\,
            I => \N__10283\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__10280\,
            I => \this_vga_signals.mult1_un40_sum_axb1_0\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__10277\,
            I => \N__10274\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10264\
        );

    \I__1447\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10264\
        );

    \I__1446\ : InMux
    port map (
            O => \N__10272\,
            I => \N__10259\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10259\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10256\
        );

    \I__1443\ : InMux
    port map (
            O => \N__10269\,
            I => \N__10253\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10248\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__10259\,
            I => \N__10248\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__10256\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__10253\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__10248\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__10241\,
            I => \this_vga_signals.if_m8_0_a3_1_1_1_cascade_\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__10238\,
            I => \N__10235\
        );

    \I__1435\ : InMux
    port map (
            O => \N__10235\,
            I => \N__10227\
        );

    \I__1434\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10224\
        );

    \I__1433\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10221\
        );

    \I__1432\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10214\
        );

    \I__1431\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10214\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10214\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__10227\,
            I => \N__10209\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__10224\,
            I => \N__10209\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__10221\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__10214\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1425\ : Odrv4
    port map (
            O => \N__10209\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__10202\,
            I => \N__10199\
        );

    \I__1423\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10196\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__10196\,
            I => \N__10193\
        );

    \I__1421\ : Span4Mux_h
    port map (
            O => \N__10193\,
            I => \N__10190\
        );

    \I__1420\ : Odrv4
    port map (
            O => \N__10190\,
            I => \this_vga_signals.vaddress_2_6\
        );

    \I__1419\ : InMux
    port map (
            O => \N__10187\,
            I => \N__10184\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__10184\,
            I => \N__10181\
        );

    \I__1417\ : Span4Mux_h
    port map (
            O => \N__10181\,
            I => \N__10178\
        );

    \I__1416\ : Odrv4
    port map (
            O => \N__10178\,
            I => \this_vga_signals.vaddress_2_5\
        );

    \I__1415\ : InMux
    port map (
            O => \N__10175\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__1414\ : InMux
    port map (
            O => \N__10172\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__1413\ : InMux
    port map (
            O => \N__10169\,
            I => \bfn_11_23_0_\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__10166\,
            I => \this_vga_signals.un4_hsynclt8_0_cascade_\
        );

    \I__1411\ : IoInMux
    port map (
            O => \N__10163\,
            I => \N__10160\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__1409\ : IoSpan4Mux
    port map (
            O => \N__10157\,
            I => \N__10154\
        );

    \I__1408\ : Span4Mux_s1_v
    port map (
            O => \N__10154\,
            I => \N__10151\
        );

    \I__1407\ : Sp12to4
    port map (
            O => \N__10151\,
            I => \N__10148\
        );

    \I__1406\ : Span12Mux_s8_v
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__1405\ : Odrv12
    port map (
            O => \N__10145\,
            I => this_vga_signals_hsync_1_i
        );

    \I__1404\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10135\
        );

    \I__1403\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10135\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__10140\,
            I => \N__10130\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__10135\,
            I => \N__10124\
        );

    \I__1400\ : InMux
    port map (
            O => \N__10134\,
            I => \N__10117\
        );

    \I__1399\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10117\
        );

    \I__1398\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10114\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__10129\,
            I => \N__10110\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10128\,
            I => \N__10104\
        );

    \I__1395\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10104\
        );

    \I__1394\ : Span4Mux_v
    port map (
            O => \N__10124\,
            I => \N__10101\
        );

    \I__1393\ : InMux
    port map (
            O => \N__10123\,
            I => \N__10098\
        );

    \I__1392\ : InMux
    port map (
            O => \N__10122\,
            I => \N__10095\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__10117\,
            I => \N__10090\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__10114\,
            I => \N__10090\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10083\
        );

    \I__1388\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10083\
        );

    \I__1387\ : InMux
    port map (
            O => \N__10109\,
            I => \N__10083\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__10104\,
            I => \N__10076\
        );

    \I__1385\ : Span4Mux_h
    port map (
            O => \N__10101\,
            I => \N__10076\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__10098\,
            I => \N__10076\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__10095\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__10090\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__10083\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__10076\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__10064\,
            I => \this_vga_signals.un3_hsynclt8_0\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__10061\,
            I => \this_vga_signals.un6_vvisibilitylto8_0_cascade_\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__10058\,
            I => \this_vga_signals.un6_vvisibilitylt9_0_cascade_\
        );

    \I__1375\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10052\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__10052\,
            I => \N__10049\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__10049\,
            I => \N__10044\
        );

    \I__1372\ : InMux
    port map (
            O => \N__10048\,
            I => \N__10041\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__10047\,
            I => \N__10038\
        );

    \I__1370\ : Span4Mux_v
    port map (
            O => \N__10044\,
            I => \N__10035\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__10041\,
            I => \N__10032\
        );

    \I__1368\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10029\
        );

    \I__1367\ : Span4Mux_h
    port map (
            O => \N__10035\,
            I => \N__10026\
        );

    \I__1366\ : Span12Mux_s11_h
    port map (
            O => \N__10032\,
            I => \N__10023\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__10029\,
            I => \N__10020\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__10026\,
            I => \this_vga_signals.vvisibility\
        );

    \I__1363\ : Odrv12
    port map (
            O => \N__10023\,
            I => \this_vga_signals.vvisibility\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__10020\,
            I => \this_vga_signals.vvisibility\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__10013\,
            I => \N__10002\
        );

    \I__1360\ : InMux
    port map (
            O => \N__10012\,
            I => \N__9994\
        );

    \I__1359\ : InMux
    port map (
            O => \N__10011\,
            I => \N__9991\
        );

    \I__1358\ : InMux
    port map (
            O => \N__10010\,
            I => \N__9988\
        );

    \I__1357\ : InMux
    port map (
            O => \N__10009\,
            I => \N__9983\
        );

    \I__1356\ : InMux
    port map (
            O => \N__10008\,
            I => \N__9983\
        );

    \I__1355\ : InMux
    port map (
            O => \N__10007\,
            I => \N__9978\
        );

    \I__1354\ : InMux
    port map (
            O => \N__10006\,
            I => \N__9978\
        );

    \I__1353\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9973\
        );

    \I__1352\ : InMux
    port map (
            O => \N__10002\,
            I => \N__9973\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9962\
        );

    \I__1350\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9962\
        );

    \I__1349\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9962\
        );

    \I__1348\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9962\
        );

    \I__1347\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9962\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__9994\,
            I => \this_vga_signals.mult1_un68_sum_axb1_395\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__9991\,
            I => \this_vga_signals.mult1_un68_sum_axb1_395\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__9988\,
            I => \this_vga_signals.mult1_un68_sum_axb1_395\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__9983\,
            I => \this_vga_signals.mult1_un68_sum_axb1_395\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__9978\,
            I => \this_vga_signals.mult1_un68_sum_axb1_395\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__9973\,
            I => \this_vga_signals.mult1_un68_sum_axb1_395\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__9962\,
            I => \this_vga_signals.mult1_un68_sum_axb1_395\
        );

    \I__1339\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9944\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__9944\,
            I => \this_vga_signals.mult1_un68_sum_ac0_1_x0\
        );

    \I__1337\ : InMux
    port map (
            O => \N__9941\,
            I => \N__9938\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__9938\,
            I => \N__9933\
        );

    \I__1335\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9928\
        );

    \I__1334\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9928\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__9933\,
            I => \this_vga_signals.mult1_un61_sum_c3_1\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__9928\,
            I => \this_vga_signals.mult1_un61_sum_c3_1\
        );

    \I__1331\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9920\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__9920\,
            I => \this_vga_signals.g0_2_x1\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__9917\,
            I => \N__9903\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__9916\,
            I => \N__9899\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__9915\,
            I => \N__9896\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__9914\,
            I => \N__9891\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__9913\,
            I => \N__9888\
        );

    \I__1324\ : InMux
    port map (
            O => \N__9912\,
            I => \N__9883\
        );

    \I__1323\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9880\
        );

    \I__1322\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9869\
        );

    \I__1321\ : InMux
    port map (
            O => \N__9909\,
            I => \N__9869\
        );

    \I__1320\ : InMux
    port map (
            O => \N__9908\,
            I => \N__9869\
        );

    \I__1319\ : InMux
    port map (
            O => \N__9907\,
            I => \N__9869\
        );

    \I__1318\ : InMux
    port map (
            O => \N__9906\,
            I => \N__9869\
        );

    \I__1317\ : InMux
    port map (
            O => \N__9903\,
            I => \N__9864\
        );

    \I__1316\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9864\
        );

    \I__1315\ : InMux
    port map (
            O => \N__9899\,
            I => \N__9855\
        );

    \I__1314\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9855\
        );

    \I__1313\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9855\
        );

    \I__1312\ : InMux
    port map (
            O => \N__9894\,
            I => \N__9855\
        );

    \I__1311\ : InMux
    port map (
            O => \N__9891\,
            I => \N__9846\
        );

    \I__1310\ : InMux
    port map (
            O => \N__9888\,
            I => \N__9846\
        );

    \I__1309\ : InMux
    port map (
            O => \N__9887\,
            I => \N__9846\
        );

    \I__1308\ : InMux
    port map (
            O => \N__9886\,
            I => \N__9846\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__9883\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__9880\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__9869\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__9864\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__9855\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__9846\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__1301\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9830\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__9830\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1\
        );

    \I__1299\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9823\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__9826\,
            I => \N__9815\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__9823\,
            I => \N__9812\
        );

    \I__1296\ : InMux
    port map (
            O => \N__9822\,
            I => \N__9805\
        );

    \I__1295\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9805\
        );

    \I__1294\ : InMux
    port map (
            O => \N__9820\,
            I => \N__9805\
        );

    \I__1293\ : InMux
    port map (
            O => \N__9819\,
            I => \N__9800\
        );

    \I__1292\ : InMux
    port map (
            O => \N__9818\,
            I => \N__9800\
        );

    \I__1291\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9797\
        );

    \I__1290\ : Span4Mux_v
    port map (
            O => \N__9812\,
            I => \N__9791\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__9805\,
            I => \N__9791\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__9800\,
            I => \N__9786\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__9797\,
            I => \N__9786\
        );

    \I__1286\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9783\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__9791\,
            I => \N__9780\
        );

    \I__1284\ : Span12Mux_s10_h
    port map (
            O => \N__9786\,
            I => \N__9777\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__9783\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__9780\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1281\ : Odrv12
    port map (
            O => \N__9777\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1280\ : InMux
    port map (
            O => \N__9770\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__1279\ : CascadeMux
    port map (
            O => \N__9767\,
            I => \N__9764\
        );

    \I__1278\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9756\
        );

    \I__1277\ : InMux
    port map (
            O => \N__9763\,
            I => \N__9756\
        );

    \I__1276\ : InMux
    port map (
            O => \N__9762\,
            I => \N__9753\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__9761\,
            I => \N__9747\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__9756\,
            I => \N__9742\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__9753\,
            I => \N__9739\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__9752\,
            I => \N__9736\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__9751\,
            I => \N__9732\
        );

    \I__1270\ : InMux
    port map (
            O => \N__9750\,
            I => \N__9727\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9727\
        );

    \I__1268\ : InMux
    port map (
            O => \N__9746\,
            I => \N__9722\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9745\,
            I => \N__9722\
        );

    \I__1266\ : Span4Mux_v
    port map (
            O => \N__9742\,
            I => \N__9716\
        );

    \I__1265\ : Span4Mux_h
    port map (
            O => \N__9739\,
            I => \N__9716\
        );

    \I__1264\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9709\
        );

    \I__1263\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9709\
        );

    \I__1262\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9709\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__9727\,
            I => \N__9704\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__9722\,
            I => \N__9704\
        );

    \I__1259\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9700\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__9716\,
            I => \N__9697\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__9709\,
            I => \N__9692\
        );

    \I__1256\ : Span4Mux_v
    port map (
            O => \N__9704\,
            I => \N__9692\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9689\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__9700\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__9697\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__9692\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__9689\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1250\ : InMux
    port map (
            O => \N__9680\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__1249\ : InMux
    port map (
            O => \N__9677\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__1248\ : InMux
    port map (
            O => \N__9674\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__1247\ : InMux
    port map (
            O => \N__9671\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__9665\,
            I => \N__9662\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__9662\,
            I => \this_vga_signals.mult1_un54_sum_axb1_1_0_0\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__9659\,
            I => \this_vga_signals.N_5_i_5_cascade_\
        );

    \I__1242\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9653\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__9653\,
            I => \this_vga_signals.N_20_0\
        );

    \I__1240\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9647\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__9647\,
            I => \this_vga_signals.g1_1_1\
        );

    \I__1238\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__9641\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_0_0\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__9638\,
            I => \this_vga_signals.g0_2_x0_cascade_\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__9635\,
            I => \this_vga_signals.g1_0_0_0_cascade_\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9629\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__9629\,
            I => \this_vga_signals.N_5_i_5\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__9626\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9620\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__9620\,
            I => \this_vga_signals.g0_i_x2_0_2_0\
        );

    \I__1229\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9614\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__9614\,
            I => \N__9611\
        );

    \I__1227\ : Span4Mux_h
    port map (
            O => \N__9611\,
            I => \N__9608\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__9608\,
            I => \this_vga_signals.if_i4_mux_0_0_0\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__9605\,
            I => \this_vga_signals.vaddress_6_cascade_\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9597\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__9601\,
            I => \N__9593\
        );

    \I__1222\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9589\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__9597\,
            I => \N__9586\
        );

    \I__1220\ : InMux
    port map (
            O => \N__9596\,
            I => \N__9583\
        );

    \I__1219\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9578\
        );

    \I__1218\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9578\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__9589\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__9586\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__9583\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__9578\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1213\ : InMux
    port map (
            O => \N__9569\,
            I => \N__9566\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__9566\,
            I => \N__9563\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__9563\,
            I => \this_vga_signals.g1_3_0\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__9560\,
            I => \N__9554\
        );

    \I__1209\ : InMux
    port map (
            O => \N__9559\,
            I => \N__9551\
        );

    \I__1208\ : InMux
    port map (
            O => \N__9558\,
            I => \N__9544\
        );

    \I__1207\ : InMux
    port map (
            O => \N__9557\,
            I => \N__9544\
        );

    \I__1206\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9544\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__9551\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__9544\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__1203\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__9536\,
            I => \N__9533\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__9533\,
            I => \this_vga_signals.vaddress_4_0_6\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__9530\,
            I => \N__9527\
        );

    \I__1199\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9524\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__9524\,
            I => \this_vga_signals.vaddress_5_0_5\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__9521\,
            I => \this_vga_signals.g2_0_cascade_\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9518\,
            I => \N__9515\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__9515\,
            I => \this_vga_signals.mult1_un54_sum_axb1_1\
        );

    \I__1194\ : InMux
    port map (
            O => \N__9512\,
            I => \N__9509\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__9509\,
            I => \this_vga_signals.g1_0_0\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9500\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9505\,
            I => \N__9497\
        );

    \I__1190\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9492\
        );

    \I__1189\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9492\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__9500\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9497\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__9492\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__9485\,
            I => \N__9482\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9477\
        );

    \I__1183\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9474\
        );

    \I__1182\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9471\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__9477\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__9474\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__9471\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__1178\ : InMux
    port map (
            O => \N__9464\,
            I => \N__9461\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__9461\,
            I => \N__9458\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__9458\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__9455\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\
        );

    \I__1174\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__9449\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_0\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__9446\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\
        );

    \I__1171\ : IoInMux
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__1169\ : IoSpan4Mux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__1168\ : Span4Mux_s2_v
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__1167\ : Span4Mux_h
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__1166\ : Span4Mux_v
    port map (
            O => \N__9428\,
            I => \N__9425\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__9425\,
            I => this_vga_signals_hvisibility_i
        );

    \I__1164\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9418\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9415\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__9418\,
            I => \this_vga_signals.SUM_3_i_0_0_3\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__9415\,
            I => \this_vga_signals.SUM_3_i_0_0_3\
        );

    \I__1160\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__9407\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9396\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9403\,
            I => \N__9391\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9402\,
            I => \N__9391\
        );

    \I__1155\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9388\
        );

    \I__1154\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9385\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__9399\,
            I => \N__9382\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__9396\,
            I => \N__9376\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__9391\,
            I => \N__9376\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9388\,
            I => \N__9371\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__9385\,
            I => \N__9371\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9382\,
            I => \N__9368\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9365\
        );

    \I__1146\ : Span4Mux_h
    port map (
            O => \N__9376\,
            I => \N__9362\
        );

    \I__1145\ : Span4Mux_v
    port map (
            O => \N__9371\,
            I => \N__9355\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__9368\,
            I => \N__9355\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__9365\,
            I => \N__9355\
        );

    \I__1142\ : Span4Mux_v
    port map (
            O => \N__9362\,
            I => \N__9348\
        );

    \I__1141\ : Span4Mux_h
    port map (
            O => \N__9355\,
            I => \N__9348\
        );

    \I__1140\ : InMux
    port map (
            O => \N__9354\,
            I => \N__9345\
        );

    \I__1139\ : InMux
    port map (
            O => \N__9353\,
            I => \N__9342\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__9348\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__9345\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__9342\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__9335\,
            I => \this_vga_signals.g0_7_0_0_cascade_\
        );

    \I__1134\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9329\,
            I => \N__9326\
        );

    \I__1132\ : Span4Mux_v
    port map (
            O => \N__9326\,
            I => \N__9323\
        );

    \I__1131\ : Odrv4
    port map (
            O => \N__9323\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i_0_1_0\
        );

    \I__1130\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9314\
        );

    \I__1129\ : InMux
    port map (
            O => \N__9319\,
            I => \N__9314\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__9314\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\
        );

    \I__1127\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9304\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9310\,
            I => \N__9304\
        );

    \I__1125\ : InMux
    port map (
            O => \N__9309\,
            I => \N__9301\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__9304\,
            I => \this_vga_signals.SUM_2_i_1_2_3\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__9301\,
            I => \this_vga_signals.SUM_2_i_1_2_3\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__9296\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i_0_0_cascade_\
        );

    \I__1121\ : InMux
    port map (
            O => \N__9293\,
            I => \N__9286\
        );

    \I__1120\ : InMux
    port map (
            O => \N__9292\,
            I => \N__9286\
        );

    \I__1119\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9283\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__9286\,
            I => \this_vga_signals.SUM_2_i_1_0_3\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__9283\,
            I => \this_vga_signals.SUM_2_i_1_0_3\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__9278\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9275\,
            I => \N__9269\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9266\
        );

    \I__1113\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9261\
        );

    \I__1112\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9261\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__9269\,
            I => \N__9258\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__9266\,
            I => \N__9255\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__9261\,
            I => \N__9252\
        );

    \I__1108\ : Span4Mux_v
    port map (
            O => \N__9258\,
            I => \N__9247\
        );

    \I__1107\ : Span4Mux_h
    port map (
            O => \N__9255\,
            I => \N__9247\
        );

    \I__1106\ : Span4Mux_h
    port map (
            O => \N__9252\,
            I => \N__9244\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__9247\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_2\
        );

    \I__1104\ : Odrv4
    port map (
            O => \N__9244\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_2\
        );

    \I__1103\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__9236\,
            I => \N__9232\
        );

    \I__1101\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9229\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__9232\,
            I => \this_vga_signals.N_3_2_1\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__9229\,
            I => \this_vga_signals.N_3_2_1\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__9224\,
            I => \this_vga_signals.N_3_2_1_cascade_\
        );

    \I__1097\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9217\
        );

    \I__1096\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9214\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__9217\,
            I => \N__9211\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__9214\,
            I => \N__9208\
        );

    \I__1093\ : Sp12to4
    port map (
            O => \N__9211\,
            I => \N__9203\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__9208\,
            I => \N__9200\
        );

    \I__1091\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9197\
        );

    \I__1090\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9194\
        );

    \I__1089\ : Odrv12
    port map (
            O => \N__9203\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__9200\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__9197\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__9194\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9180\
        );

    \I__1084\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9175\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9183\,
            I => \N__9175\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__9180\,
            I => \this_vga_signals.mult1_un68_sum_axb2_1\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__9175\,
            I => \this_vga_signals.mult1_un68_sum_axb2_1\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__9170\,
            I => \this_vga_signals.mult1_un68_sum_axb2_1_cascade_\
        );

    \I__1079\ : InMux
    port map (
            O => \N__9167\,
            I => \N__9161\
        );

    \I__1078\ : InMux
    port map (
            O => \N__9166\,
            I => \N__9156\
        );

    \I__1077\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9156\
        );

    \I__1076\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9153\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__9161\,
            I => \N__9150\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__9156\,
            I => \N__9147\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9153\,
            I => \N__9144\
        );

    \I__1072\ : Span4Mux_v
    port map (
            O => \N__9150\,
            I => \N__9141\
        );

    \I__1071\ : Span4Mux_h
    port map (
            O => \N__9147\,
            I => \N__9138\
        );

    \I__1070\ : Odrv12
    port map (
            O => \N__9144\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__9141\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__9138\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__9128\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__9125\,
            I => \N__9122\
        );

    \I__1064\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9118\
        );

    \I__1063\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9115\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__9118\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__9115\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9107\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__1058\ : Span4Mux_v
    port map (
            O => \N__9104\,
            I => \N__9100\
        );

    \I__1057\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9097\
        );

    \I__1056\ : Span4Mux_v
    port map (
            O => \N__9100\,
            I => \N__9094\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__9097\,
            I => \N__9088\
        );

    \I__1054\ : Sp12to4
    port map (
            O => \N__9094\,
            I => \N__9083\
        );

    \I__1053\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9076\
        );

    \I__1052\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9076\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9076\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__9088\,
            I => \N__9073\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9087\,
            I => \N__9070\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9067\
        );

    \I__1047\ : Odrv12
    port map (
            O => \N__9083\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__9076\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__9073\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__9070\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9067\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__9056\,
            I => \this_vga_signals.SUM_3_i_0_0_3_cascade_\
        );

    \I__1041\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9050\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__9050\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_0\
        );

    \I__1039\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9044\,
            I => \this_vga_signals.vaddress_1_5\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__9041\,
            I => \this_vga_signals.vaddress_1_6_cascade_\
        );

    \I__1036\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__9035\,
            I => \this_vga_signals.mult1_un54_sum_axb1_1_0_1\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__9032\,
            I => \N__9022\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__9031\,
            I => \N__9016\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__9030\,
            I => \N__9013\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__9029\,
            I => \N__9009\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9002\
        );

    \I__1029\ : InMux
    port map (
            O => \N__9027\,
            I => \N__8997\
        );

    \I__1028\ : InMux
    port map (
            O => \N__9026\,
            I => \N__8997\
        );

    \I__1027\ : InMux
    port map (
            O => \N__9025\,
            I => \N__8990\
        );

    \I__1026\ : InMux
    port map (
            O => \N__9022\,
            I => \N__8990\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9021\,
            I => \N__8990\
        );

    \I__1024\ : InMux
    port map (
            O => \N__9020\,
            I => \N__8981\
        );

    \I__1023\ : InMux
    port map (
            O => \N__9019\,
            I => \N__8981\
        );

    \I__1022\ : InMux
    port map (
            O => \N__9016\,
            I => \N__8981\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9013\,
            I => \N__8981\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9012\,
            I => \N__8976\
        );

    \I__1019\ : InMux
    port map (
            O => \N__9009\,
            I => \N__8976\
        );

    \I__1018\ : InMux
    port map (
            O => \N__9008\,
            I => \N__8967\
        );

    \I__1017\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8967\
        );

    \I__1016\ : InMux
    port map (
            O => \N__9006\,
            I => \N__8967\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8967\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__9002\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__8997\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__8990\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__8981\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__8976\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__8967\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1008\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8951\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__8951\,
            I => \this_vga_signals.g0_12_x1\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__8948\,
            I => \this_vga_signals.g0_0_2_1_0_cascade_\
        );

    \I__1005\ : InMux
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__8939\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_0\
        );

    \I__1002\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8932\
        );

    \I__1001\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8929\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__8932\,
            I => \this_vga_signals.g0_0_2\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__8929\,
            I => \this_vga_signals.g0_0_2\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__997\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8917\
        );

    \I__996\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8914\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__8917\,
            I => \N__8911\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__8914\,
            I => \this_vga_signals.vaddress_6_5\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__8911\,
            I => \this_vga_signals.vaddress_6_5\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__8906\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_1_0_cascade_\
        );

    \I__991\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__8900\,
            I => \N__8897\
        );

    \I__989\ : Odrv4
    port map (
            O => \N__8897\,
            I => \this_vga_signals.g0_0_2_0\
        );

    \I__988\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__8891\,
            I => \this_vga_signals.N_236\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__8888\,
            I => \this_vga_signals.mult1_un68_sum_axb1_395_cascade_\
        );

    \I__985\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8882\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__8882\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0\
        );

    \I__983\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8876\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__8876\,
            I => \N__8869\
        );

    \I__981\ : InMux
    port map (
            O => \N__8875\,
            I => \N__8864\
        );

    \I__980\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8864\
        );

    \I__979\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8859\
        );

    \I__978\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8859\
        );

    \I__977\ : Odrv4
    port map (
            O => \N__8869\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__8864\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__8859\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__8852\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_cascade_\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__8849\,
            I => \this_vga_signals.g0_5_2_cascade_\
        );

    \I__972\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__8843\,
            I => \this_vga_signals.g1_2\
        );

    \I__970\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__8837\,
            I => \this_vga_signals.mult1_un68_sum_ac0_1_x1\
        );

    \I__968\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__8831\,
            I => \this_vga_signals.mult1_un68_sum_ac0_1\
        );

    \I__966\ : InMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__8825\,
            I => \this_vga_signals.N_3_1\
        );

    \I__964\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__8819\,
            I => \this_vga_signals.N_7\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__8816\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_cascade_\
        );

    \I__961\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__8810\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_0_0\
        );

    \I__959\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8804\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__8804\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__8801\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__8798\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4_cascade_\
        );

    \I__955\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__8792\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__8789\,
            I => \this_vga_signals.N_1_4_1_cascade_\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__8786\,
            I => \this_vga_signals.M_pcounter_q_3_0_cascade_\
        );

    \I__951\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8777\
        );

    \I__950\ : InMux
    port map (
            O => \N__8782\,
            I => \N__8777\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__8777\,
            I => \N__8774\
        );

    \I__948\ : Span4Mux_h
    port map (
            O => \N__8774\,
            I => \N__8771\
        );

    \I__947\ : Odrv4
    port map (
            O => \N__8771\,
            I => \this_vga_signals.N_2_0\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__8768\,
            I => \this_vga_signals.N_2_0_cascade_\
        );

    \I__945\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8761\
        );

    \I__944\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8758\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__8761\,
            I => \this_vga_signals.M_pcounter_q_i_3_0\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__8758\,
            I => \this_vga_signals.M_pcounter_q_i_3_0\
        );

    \I__941\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8747\
        );

    \I__940\ : InMux
    port map (
            O => \N__8752\,
            I => \N__8747\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8743\
        );

    \I__938\ : InMux
    port map (
            O => \N__8746\,
            I => \N__8740\
        );

    \I__937\ : Span4Mux_h
    port map (
            O => \N__8743\,
            I => \N__8737\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__8740\,
            I => \this_vga_signals.N_3_0\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__8737\,
            I => \this_vga_signals.N_3_0\
        );

    \I__934\ : InMux
    port map (
            O => \N__8732\,
            I => \N__8725\
        );

    \I__933\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8725\
        );

    \I__932\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8722\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__8725\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__8722\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__928\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8709\
        );

    \I__927\ : InMux
    port map (
            O => \N__8713\,
            I => \N__8704\
        );

    \I__926\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8704\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__8709\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__8704\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__8699\,
            I => \N__8694\
        );

    \I__922\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8688\
        );

    \I__921\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8688\
        );

    \I__920\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8683\
        );

    \I__919\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8683\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__8688\,
            I => \this_vga_signals.M_pcounter_q_i_3_1\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__8683\,
            I => \this_vga_signals.M_pcounter_q_i_3_1\
        );

    \I__916\ : InMux
    port map (
            O => \N__8678\,
            I => \N__8675\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__8675\,
            I => \this_vga_signals.M_pcounter_q_3_1\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__913\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__911\ : Span4Mux_h
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__910\ : Span4Mux_v
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__8657\,
            I => \M_this_vga_signals_address_6\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__907\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__905\ : Span4Mux_v
    port map (
            O => \N__8645\,
            I => \N__8640\
        );

    \I__904\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8635\
        );

    \I__903\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8635\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__8640\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__8635\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__8630\,
            I => \N__8627\
        );

    \I__899\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__897\ : Span4Mux_h
    port map (
            O => \N__8621\,
            I => \N__8618\
        );

    \I__896\ : Span4Mux_v
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__8615\,
            I => \M_this_vga_signals_address_3\
        );

    \I__894\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__892\ : Span4Mux_v
    port map (
            O => \N__8606\,
            I => \N__8603\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__8603\,
            I => \this_vga_signals.vaddress_1_0_6\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__8600\,
            I => \this_vga_signals.g1_2_0_cascade_\
        );

    \I__889\ : InMux
    port map (
            O => \N__8597\,
            I => \N__8594\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__887\ : Odrv12
    port map (
            O => \N__8591\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2_0_0\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__885\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__8582\,
            I => \N__8579\
        );

    \I__883\ : Odrv12
    port map (
            O => \N__8579\,
            I => \this_vga_signals.g1_3\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__881\ : InMux
    port map (
            O => \N__8573\,
            I => \N__8570\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__879\ : Span4Mux_h
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__8564\,
            I => \this_vga_signals.M_hcounter_q_RNI8OIBAZ0Z_3\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__8561\,
            I => \N__8557\
        );

    \I__876\ : InMux
    port map (
            O => \N__8560\,
            I => \N__8554\
        );

    \I__875\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8551\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__8554\,
            I => \N__8548\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__8551\,
            I => \N__8545\
        );

    \I__872\ : Span4Mux_v
    port map (
            O => \N__8548\,
            I => \N__8542\
        );

    \I__871\ : Span4Mux_h
    port map (
            O => \N__8545\,
            I => \N__8539\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__8542\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__869\ : Odrv4
    port map (
            O => \N__8539\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__868\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__866\ : Span4Mux_h
    port map (
            O => \N__8528\,
            I => \N__8525\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__8525\,
            I => \this_vga_signals.if_N_8_i_0\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__8522\,
            I => \this_vga_signals.g0_9_1_cascade_\
        );

    \I__863\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8516\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__8516\,
            I => \this_vga_signals.g0_12_x0\
        );

    \I__861\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__8510\,
            I => \this_vga_signals.g0_5_0\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__8507\,
            I => \this_vga_signals.N_6_0_cascade_\
        );

    \I__858\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8501\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__8501\,
            I => \this_vga_signals.N_5\
        );

    \I__856\ : InMux
    port map (
            O => \N__8498\,
            I => \N__8495\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__8495\,
            I => \N__8492\
        );

    \I__854\ : Odrv12
    port map (
            O => \N__8492\,
            I => \this_vga_signals.d_N_3_i_0_0_0\
        );

    \I__853\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8486\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__8483\,
            I => \this_vga_signals.g0_3_cascade_\
        );

    \I__850\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8476\
        );

    \I__849\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8473\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__8476\,
            I => \this_vga_signals.mult1_un68_sum_axb1\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__8473\,
            I => \this_vga_signals.mult1_un68_sum_axb1\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__8468\,
            I => \this_vga_signals.N_5_1_cascade_\
        );

    \I__845\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__8462\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__8459\,
            I => \this_vga_signals.if_i1_mux_0_cascade_\
        );

    \I__842\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8453\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__8453\,
            I => \this_vga_signals.g1_6_0\
        );

    \I__840\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8447\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__8447\,
            I => \this_vga_signals.mult1_un75_sum_c3_0_0\
        );

    \I__838\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8441\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__8441\,
            I => \this_vga_signals.if_m1_3\
        );

    \I__836\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__8435\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__8432\,
            I => \this_vga_signals.if_m1_3_cascade_\
        );

    \I__833\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8425\
        );

    \I__832\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8422\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8425\,
            I => \this_vga_signals.mult1_un68_sum_axbxc2\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8422\,
            I => \this_vga_signals.mult1_un68_sum_axbxc2\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__8417\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\
        );

    \I__828\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__8411\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_i\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__8408\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_i_cascade_\
        );

    \I__825\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8402\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__8402\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0\
        );

    \I__823\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__8396\,
            I => \this_vga_signals.if_N_2_1_0_0\
        );

    \I__821\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__8390\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__8387\,
            I => \this_vga_signals.vaddress_1_0_5_cascade_\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__8384\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_cascade_\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__8381\,
            I => \N__8378\
        );

    \I__816\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8375\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__8375\,
            I => \N__8372\
        );

    \I__814\ : Span4Mux_v
    port map (
            O => \N__8372\,
            I => \N__8369\
        );

    \I__813\ : Span4Mux_v
    port map (
            O => \N__8369\,
            I => \N__8366\
        );

    \I__812\ : Odrv4
    port map (
            O => \N__8366\,
            I => \M_this_vga_signals_address_7\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__8363\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_cascade_\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__8360\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_cascade_\
        );

    \I__809\ : CascadeMux
    port map (
            O => \N__8357\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_cascade_\
        );

    \I__808\ : InMux
    port map (
            O => \N__8354\,
            I => \N__8351\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__8351\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_0\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__8348\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_cascade_\
        );

    \I__805\ : InMux
    port map (
            O => \N__8345\,
            I => \N__8342\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8342\,
            I => \this_vga_signals.mult1_un89_sum_c3\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__802\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8333\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__8333\,
            I => \N__8330\
        );

    \I__800\ : Span4Mux_v
    port map (
            O => \N__8330\,
            I => \N__8327\
        );

    \I__799\ : Span4Mux_v
    port map (
            O => \N__8327\,
            I => \N__8324\
        );

    \I__798\ : Odrv4
    port map (
            O => \N__8324\,
            I => \M_this_vga_signals_address_0\
        );

    \I__797\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8311\
        );

    \I__796\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8311\
        );

    \I__795\ : InMux
    port map (
            O => \N__8319\,
            I => \N__8308\
        );

    \I__794\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8301\
        );

    \I__793\ : InMux
    port map (
            O => \N__8317\,
            I => \N__8301\
        );

    \I__792\ : InMux
    port map (
            O => \N__8316\,
            I => \N__8301\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__8311\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__8308\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__8301\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__788\ : InMux
    port map (
            O => \N__8294\,
            I => \N__8291\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__8291\,
            I => \this_vga_signals.d_N_11\
        );

    \I__786\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8285\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__8285\,
            I => \this_vga_signals.d_N_12\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__8282\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_cascade_\
        );

    \I__783\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8273\
        );

    \I__782\ : InMux
    port map (
            O => \N__8278\,
            I => \N__8273\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__8273\,
            I => \this_vga_signals.mult1_un75_sum_axb1\
        );

    \I__780\ : InMux
    port map (
            O => \N__8270\,
            I => \N__8265\
        );

    \I__779\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8262\
        );

    \I__778\ : CascadeMux
    port map (
            O => \N__8268\,
            I => \N__8259\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__8265\,
            I => \N__8253\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__8262\,
            I => \N__8253\
        );

    \I__775\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8248\
        );

    \I__774\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8248\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__8253\,
            I => \this_vga_signals.mult1_un68_sum_axbxc1\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8248\,
            I => \this_vga_signals.mult1_un68_sum_axbxc1\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__8243\,
            I => \N__8240\
        );

    \I__770\ : InMux
    port map (
            O => \N__8240\,
            I => \N__8237\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__8237\,
            I => \N__8234\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__8234\,
            I => \M_this_vga_signals_address_5\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__8231\,
            I => \N__8228\
        );

    \I__766\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8225\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__8225\,
            I => \M_this_vga_signals_address_4\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__8222\,
            I => \this_vga_signals.if_N_9_1_cascade_\
        );

    \I__763\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8216\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__8216\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__8213\,
            I => \this_vga_signals.if_m1_0_cascade_\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__8210\,
            I => \this_vga_signals.mult1_un82_sum_c3_cascade_\
        );

    \I__759\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8204\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__8204\,
            I => \this_vga_signals.N_2_7_0\
        );

    \I__757\ : InMux
    port map (
            O => \N__8201\,
            I => \N__8197\
        );

    \I__756\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8194\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__8197\,
            I => \this_vga_signals.mult1_un75_sum_c2_0\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__8194\,
            I => \this_vga_signals.mult1_un75_sum_c2_0\
        );

    \I__753\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__8186\,
            I => \N__8183\
        );

    \I__751\ : Span4Mux_h
    port map (
            O => \N__8183\,
            I => \N__8180\
        );

    \I__750\ : Span4Mux_v
    port map (
            O => \N__8180\,
            I => \N__8174\
        );

    \I__749\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8169\
        );

    \I__748\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8169\
        );

    \I__747\ : InMux
    port map (
            O => \N__8177\,
            I => \N__8166\
        );

    \I__746\ : Odrv4
    port map (
            O => \N__8174\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8169\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__8166\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__743\ : InMux
    port map (
            O => \N__8159\,
            I => \N__8155\
        );

    \I__742\ : InMux
    port map (
            O => \N__8158\,
            I => \N__8152\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__8155\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__8152\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0\
        );

    \I__739\ : InMux
    port map (
            O => \N__8147\,
            I => \N__8144\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__8144\,
            I => \N__8141\
        );

    \I__737\ : Odrv12
    port map (
            O => \N__8141\,
            I => \this_vga_ramdac.m19\
        );

    \I__736\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8134\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__8137\,
            I => \N__8131\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__8134\,
            I => \N__8128\
        );

    \I__733\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8125\
        );

    \I__732\ : Odrv12
    port map (
            O => \N__8128\,
            I => \this_vga_ramdac.N_1766_reto\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__8125\,
            I => \this_vga_ramdac.N_1766_reto\
        );

    \I__730\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8117\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__8117\,
            I => \this_vga_signals.M_this_vga_signals_pixel_clk_0_0\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__8114\,
            I => \N__8108\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__8113\,
            I => \N__8105\
        );

    \I__726\ : InMux
    port map (
            O => \N__8112\,
            I => \N__8092\
        );

    \I__725\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8092\
        );

    \I__724\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8092\
        );

    \I__723\ : InMux
    port map (
            O => \N__8105\,
            I => \N__8092\
        );

    \I__722\ : InMux
    port map (
            O => \N__8104\,
            I => \N__8092\
        );

    \I__721\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8089\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__8092\,
            I => \M_pcounter_q_ret_2_RNIRAOL5\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__8089\,
            I => \M_pcounter_q_ret_2_RNIRAOL5\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__8084\,
            I => \M_pcounter_q_ret_2_RNIRAOL5_cascade_\
        );

    \I__717\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__715\ : Odrv12
    port map (
            O => \N__8075\,
            I => \this_vga_ramdac.i2_mux_0\
        );

    \I__714\ : InMux
    port map (
            O => \N__8072\,
            I => \N__8069\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__8069\,
            I => \N__8066\
        );

    \I__712\ : Span4Mux_v
    port map (
            O => \N__8066\,
            I => \N__8062\
        );

    \I__711\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8059\
        );

    \I__710\ : Odrv4
    port map (
            O => \N__8062\,
            I => \this_vga_ramdac.N_1767_reto\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__8059\,
            I => \this_vga_ramdac.N_1767_reto\
        );

    \I__708\ : InMux
    port map (
            O => \N__8054\,
            I => \N__8051\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__8051\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__8048\,
            I => \N__8045\
        );

    \I__705\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8042\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__8042\,
            I => \N__8039\
        );

    \I__703\ : Odrv4
    port map (
            O => \N__8039\,
            I => \M_this_vga_signals_address_2\
        );

    \I__702\ : CascadeMux
    port map (
            O => \N__8036\,
            I => \N__8033\
        );

    \I__701\ : InMux
    port map (
            O => \N__8033\,
            I => \N__8030\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__8030\,
            I => \N__8027\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__698\ : Span4Mux_v
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__8021\,
            I => \M_this_vga_signals_address_1\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__8018\,
            I => \this_vga_signals.mult1_un75_sum_c2_0_cascade_\
        );

    \I__695\ : InMux
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__8012\,
            I => \this_vga_signals.if_m7_0_x4_0\
        );

    \I__693\ : InMux
    port map (
            O => \N__8009\,
            I => \N__8004\
        );

    \I__692\ : InMux
    port map (
            O => \N__8008\,
            I => \N__7999\
        );

    \I__691\ : InMux
    port map (
            O => \N__8007\,
            I => \N__7999\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__8004\,
            I => \N__7994\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7991\
        );

    \I__688\ : InMux
    port map (
            O => \N__7998\,
            I => \N__7988\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__7997\,
            I => \N__7983\
        );

    \I__686\ : Span4Mux_v
    port map (
            O => \N__7994\,
            I => \N__7980\
        );

    \I__685\ : Span4Mux_v
    port map (
            O => \N__7991\,
            I => \N__7977\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__7988\,
            I => \N__7974\
        );

    \I__683\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7969\
        );

    \I__682\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7969\
        );

    \I__681\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7966\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__7980\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__679\ : Odrv4
    port map (
            O => \N__7977\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__678\ : Odrv12
    port map (
            O => \N__7974\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__7969\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__7966\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__675\ : InMux
    port map (
            O => \N__7955\,
            I => \N__7952\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__7952\,
            I => \N__7949\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__7949\,
            I => \this_vga_ramdac.i2_mux\
        );

    \I__672\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7942\
        );

    \I__671\ : InMux
    port map (
            O => \N__7945\,
            I => \N__7939\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__7942\,
            I => \this_vga_ramdac.N_1764_reto\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__7939\,
            I => \this_vga_ramdac.N_1764_reto\
        );

    \I__668\ : InMux
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__7928\,
            I => \this_vga_ramdac.m16\
        );

    \I__665\ : InMux
    port map (
            O => \N__7925\,
            I => \N__7922\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__7922\,
            I => \N__7918\
        );

    \I__663\ : CascadeMux
    port map (
            O => \N__7921\,
            I => \N__7915\
        );

    \I__662\ : Span4Mux_v
    port map (
            O => \N__7918\,
            I => \N__7912\
        );

    \I__661\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7909\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__7912\,
            I => \this_vga_ramdac.N_1765_reto\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__7909\,
            I => \this_vga_ramdac.N_1765_reto\
        );

    \I__658\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7901\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__7901\,
            I => \N__7898\
        );

    \I__656\ : Odrv12
    port map (
            O => \N__7898\,
            I => port_clk_c
        );

    \I__655\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7892\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__7892\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__653\ : InMux
    port map (
            O => \N__7889\,
            I => \N__7886\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__7883\,
            I => \this_vga_ramdac.N_24_mux\
        );

    \I__650\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7876\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__7879\,
            I => \N__7873\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__7876\,
            I => \N__7870\
        );

    \I__647\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7867\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__7870\,
            I => \this_vga_ramdac.N_1762_reto\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__7867\,
            I => \this_vga_ramdac.N_1762_reto\
        );

    \I__644\ : InMux
    port map (
            O => \N__7862\,
            I => \N__7859\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__7859\,
            I => \N__7856\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__7856\,
            I => \this_vga_ramdac.m6\
        );

    \I__641\ : InMux
    port map (
            O => \N__7853\,
            I => \N__7849\
        );

    \I__640\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7846\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__7849\,
            I => \this_vga_ramdac.N_1763_reto\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__7846\,
            I => \this_vga_ramdac.N_1763_reto\
        );

    \I__637\ : IoInMux
    port map (
            O => \N__7841\,
            I => \N__7838\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__7838\,
            I => \N__7835\
        );

    \I__635\ : Span12Mux_s7_v
    port map (
            O => \N__7835\,
            I => \N__7832\
        );

    \I__634\ : Odrv12
    port map (
            O => \N__7832\,
            I => this_vga_signals_vvisibility_i
        );

    \I__633\ : IoInMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__7826\,
            I => \N__7823\
        );

    \I__631\ : IoSpan4Mux
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__630\ : Span4Mux_s3_h
    port map (
            O => \N__7820\,
            I => \N__7817\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__7817\,
            I => rgb_c_2
        );

    \I__628\ : IoInMux
    port map (
            O => \N__7814\,
            I => \N__7811\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__7811\,
            I => \N__7808\
        );

    \I__626\ : IoSpan4Mux
    port map (
            O => \N__7808\,
            I => \N__7805\
        );

    \I__625\ : Span4Mux_s2_h
    port map (
            O => \N__7805\,
            I => \N__7802\
        );

    \I__624\ : Odrv4
    port map (
            O => \N__7802\,
            I => rgb_c_1
        );

    \I__623\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7787\
        );

    \I__622\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7787\
        );

    \I__621\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7787\
        );

    \I__620\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7787\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__7787\,
            I => \N__7782\
        );

    \I__618\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7777\
        );

    \I__617\ : InMux
    port map (
            O => \N__7785\,
            I => \N__7777\
        );

    \I__616\ : Span4Mux_h
    port map (
            O => \N__7782\,
            I => \N__7774\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__7777\,
            I => \N__7771\
        );

    \I__614\ : Sp12to4
    port map (
            O => \N__7774\,
            I => \N__7766\
        );

    \I__613\ : Span12Mux_s7_h
    port map (
            O => \N__7771\,
            I => \N__7766\
        );

    \I__612\ : Odrv12
    port map (
            O => \N__7766\,
            I => \M_this_vram_read_data_0\
        );

    \I__611\ : InMux
    port map (
            O => \N__7763\,
            I => \N__7753\
        );

    \I__610\ : InMux
    port map (
            O => \N__7762\,
            I => \N__7753\
        );

    \I__609\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7744\
        );

    \I__608\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7744\
        );

    \I__607\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7744\
        );

    \I__606\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7744\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__7753\,
            I => \N__7739\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__7744\,
            I => \N__7739\
        );

    \I__603\ : Span4Mux_v
    port map (
            O => \N__7739\,
            I => \N__7736\
        );

    \I__602\ : Span4Mux_v
    port map (
            O => \N__7736\,
            I => \N__7733\
        );

    \I__601\ : Odrv4
    port map (
            O => \N__7733\,
            I => \M_this_vram_read_data_3\
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__7730\,
            I => \N__7723\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__7729\,
            I => \N__7720\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__7728\,
            I => \N__7717\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__7727\,
            I => \N__7714\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__7726\,
            I => \N__7711\
        );

    \I__595\ : InMux
    port map (
            O => \N__7723\,
            I => \N__7706\
        );

    \I__594\ : InMux
    port map (
            O => \N__7720\,
            I => \N__7706\
        );

    \I__593\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7703\
        );

    \I__592\ : InMux
    port map (
            O => \N__7714\,
            I => \N__7698\
        );

    \I__591\ : InMux
    port map (
            O => \N__7711\,
            I => \N__7698\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__7706\,
            I => \N__7691\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__7703\,
            I => \N__7691\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__7698\,
            I => \N__7691\
        );

    \I__587\ : Span4Mux_v
    port map (
            O => \N__7691\,
            I => \N__7688\
        );

    \I__586\ : Span4Mux_v
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__7685\,
            I => \M_this_vram_read_data_2\
        );

    \I__584\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7672\
        );

    \I__583\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7672\
        );

    \I__582\ : InMux
    port map (
            O => \N__7680\,
            I => \N__7667\
        );

    \I__581\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7667\
        );

    \I__580\ : InMux
    port map (
            O => \N__7678\,
            I => \N__7662\
        );

    \I__579\ : InMux
    port map (
            O => \N__7677\,
            I => \N__7662\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__7672\,
            I => \N__7655\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__7667\,
            I => \N__7655\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__7662\,
            I => \N__7655\
        );

    \I__575\ : Span12Mux_v
    port map (
            O => \N__7655\,
            I => \N__7652\
        );

    \I__574\ : Odrv12
    port map (
            O => \N__7652\,
            I => \M_this_vram_read_data_1\
        );

    \I__573\ : IoInMux
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__7646\,
            I => \this_vga_signals.N_340_0\
        );

    \I__571\ : IoInMux
    port map (
            O => \N__7643\,
            I => \N__7640\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__7640\,
            I => \N_198_i\
        );

    \I__569\ : IoInMux
    port map (
            O => \N__7637\,
            I => \N__7634\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__7634\,
            I => \N__7631\
        );

    \I__567\ : Span4Mux_s2_h
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__565\ : Span12Mux_v
    port map (
            O => \N__7625\,
            I => \N__7622\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__7622\,
            I => rgb_c_0
        );

    \I__563\ : IoInMux
    port map (
            O => \N__7619\,
            I => \N__7616\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__7616\,
            I => \N__7613\
        );

    \I__561\ : IoSpan4Mux
    port map (
            O => \N__7613\,
            I => \N__7610\
        );

    \I__560\ : Span4Mux_s2_h
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__559\ : Span4Mux_v
    port map (
            O => \N__7607\,
            I => \N__7604\
        );

    \I__558\ : Odrv4
    port map (
            O => \N__7604\,
            I => rgb_c_4
        );

    \I__557\ : IoInMux
    port map (
            O => \N__7601\,
            I => \N__7598\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__7598\,
            I => \N__7595\
        );

    \I__555\ : Span4Mux_s3_h
    port map (
            O => \N__7595\,
            I => \N__7592\
        );

    \I__554\ : Odrv4
    port map (
            O => \N__7592\,
            I => port_nmib_0_i
        );

    \I__553\ : IoInMux
    port map (
            O => \N__7589\,
            I => \N__7586\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__7586\,
            I => \N__7583\
        );

    \I__551\ : Span4Mux_s3_h
    port map (
            O => \N__7583\,
            I => \N__7580\
        );

    \I__550\ : Odrv4
    port map (
            O => \N__7580\,
            I => rgb_c_3
        );

    \I__549\ : IoInMux
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__547\ : Span4Mux_s3_h
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__546\ : Span4Mux_v
    port map (
            O => \N__7568\,
            I => \N__7565\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__7565\,
            I => rgb_c_5
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_21_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_17_0_\
        );

    \IN_MUX_bfv_21_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.sprites_addr_cry_8\,
            carryinitout => \bfn_21_18_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_sprites_address_q_cry_7\,
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_30_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_30_23_0_\
        );

    \IN_MUX_bfv_30_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_external_address_q_cry_7\,
            carryinitout => \bfn_30_24_0_\
        );

    \IN_MUX_bfv_17_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_23_0_\
        );

    \IN_MUX_bfv_17_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_data_count_q_cry_7\,
            carryinitout => \bfn_17_24_0_\
        );

    \IN_MUX_bfv_17_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO\,
            carryinitout => \bfn_17_25_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIRO2H5_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14996\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_515_g\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIADVP5_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7649\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_340_0_g\
        );

    \this_reset_cond.M_stage_q_RNI6VB7_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14519\,
            GLOBALBUFFEROUTPUT => \M_this_state_q_nss_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIADVP5_9_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14263\,
            in2 => \_gnd_net_\,
            in3 => \N__11567\,
            lcout => \this_vga_signals.N_340_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_rw_obuf_RNO_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__14431\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13209\,
            lcout => \N_198_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7880\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7998\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8138\,
            in2 => \_gnd_net_\,
            in3 => \N__8009\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIA0384_9_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13213\,
            in2 => \_gnd_net_\,
            in3 => \N__10055\,
            lcout => port_nmib_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7925\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8008\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8072\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_0_9_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10048\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => this_vga_signals_vvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7946\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7987\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7986\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7853\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100011011"
        )
    port map (
            in0 => \N__7763\,
            in1 => \N__7678\,
            in2 => \N__7730\,
            in3 => \N__7786\,
            lcout => \this_vga_ramdac.m6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100100101"
        )
    port map (
            in0 => \N__7762\,
            in1 => \N__7677\,
            in2 => \N__7729\,
            in3 => \N__7785\,
            lcout => \this_vga_ramdac.i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__7799\,
            in1 => \N__7758\,
            in2 => \_gnd_net_\,
            in3 => \N__7682\,
            lcout => \this_vga_ramdac.N_24_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110101110001"
        )
    port map (
            in0 => \N__7761\,
            in1 => \N__7680\,
            in2 => \N__7726\,
            in3 => \N__7798\,
            lcout => \this_vga_ramdac.m19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101100111"
        )
    port map (
            in0 => \N__7759\,
            in1 => \N__7679\,
            in2 => \N__7727\,
            in3 => \N__7796\,
            lcout => \this_vga_ramdac.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000110110111"
        )
    port map (
            in0 => \N__7797\,
            in1 => \N__7760\,
            in2 => \N__7728\,
            in3 => \N__7681\,
            lcout => \this_vga_ramdac.m16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_x4_0_0_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__8279\,
            in1 => \_gnd_net_\,
            in2 => \N__8268\,
            in3 => \N__8319\,
            lcout => \this_vga_signals.if_m7_0_x4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__9762\,
            in1 => \N__8258\,
            in2 => \N__9826\,
            in3 => \N__8278\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_q_ret_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__9401\,
            in1 => \N__8112\,
            in2 => \N__7997\,
            in3 => \N__14524\,
            lcout => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7895\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__14522\,
            in1 => \N__7945\,
            in2 => \N__8114\,
            in3 => \N__7955\,
            lcout => \this_vga_ramdac.N_1764_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__7934\,
            in1 => \N__8111\,
            in2 => \N__7921\,
            in3 => \N__14523\,
            lcout => \this_vga_ramdac.N_1765_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__7889\,
            in1 => \N__8104\,
            in2 => \N__7879\,
            in3 => \N__14520\,
            lcout => \this_vga_ramdac.N_1762_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__14521\,
            in1 => \N__7852\,
            in2 => \N__8113\,
            in3 => \N__7862\,
            lcout => \this_vga_ramdac.N_1763_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__8147\,
            in1 => \N__8103\,
            in2 => \N__8137\,
            in3 => \N__14533\,
            lcout => \this_vga_ramdac.N_1766_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_2_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8783\,
            in2 => \_gnd_net_\,
            in3 => \N__8753\,
            lcout => \this_vga_signals.M_this_vga_signals_pixel_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_2_RNIRAOL5_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__8120\,
            in1 => \N__8782\,
            in2 => \_gnd_net_\,
            in3 => \N__8752\,
            lcout => \M_pcounter_q_ret_2_RNIRAOL5\,
            ltout => \M_pcounter_q_ret_2_RNIRAOL5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__14534\,
            in1 => \N__8065\,
            in2 => \N__8084\,
            in3 => \N__8081\,
            lcout => \this_vga_ramdac.N_1767_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8054\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIHM2SG2_9_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9404\,
            in2 => \_gnd_net_\,
            in3 => \N__8189\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNICQMCG5_9_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__8179\,
            in1 => \N__8201\,
            in2 => \N__9399\,
            in3 => \N__8159\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011011101"
        )
    port map (
            in0 => \N__9820\,
            in1 => \N__9763\,
            in2 => \_gnd_net_\,
            in3 => \N__8316\,
            lcout => \this_vga_signals.mult1_un75_sum_c2_0\,
            ltout => \this_vga_signals.mult1_un75_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100010111"
        )
    port map (
            in0 => \N__11977\,
            in1 => \N__11936\,
            in2 => \N__8018\,
            in3 => \N__8015\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100011011"
        )
    port map (
            in0 => \N__9822\,
            in1 => \N__11938\,
            in2 => \N__8222\,
            in3 => \N__8178\,
            lcout => \this_vga_signals.mult1_un89_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000101111000"
        )
    port map (
            in0 => \N__8269\,
            in1 => \N__8317\,
            in2 => \N__8561\,
            in3 => \N__8219\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m5_i_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001001001100"
        )
    port map (
            in0 => \N__8318\,
            in1 => \N__11935\,
            in2 => \N__9767\,
            in3 => \N__9821\,
            lcout => \this_vga_signals.N_2_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m1_0_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8643\,
            in1 => \N__9166\,
            in2 => \N__9761\,
            in3 => \N__9272\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100000111110"
        )
    port map (
            in0 => \N__11931\,
            in1 => \N__9818\,
            in2 => \N__8213\,
            in3 => \N__8534\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__8270\,
            in1 => \_gnd_net_\,
            in2 => \N__8210\,
            in3 => \N__8320\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101000100"
        )
    port map (
            in0 => \N__8288\,
            in1 => \N__8294\,
            in2 => \N__8576\,
            in3 => \N__8207\,
            lcout => \this_vga_signals.mult1_un89_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8644\,
            in1 => \N__9165\,
            in2 => \_gnd_net_\,
            in3 => \N__9273\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8200\,
            in1 => \N__8177\,
            in2 => \_gnd_net_\,
            in3 => \N__8158\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIAPUMSC_9_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__9400\,
            in1 => \N__8354\,
            in2 => \N__8348\,
            in3 => \N__8345\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNICOOCQ_1_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101001110"
        )
    port map (
            in0 => \N__8321\,
            in1 => \N__9819\,
            in2 => \N__11939\,
            in3 => \N__9750\,
            lcout => \this_vga_signals.d_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI97PTA_1_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__11937\,
            in1 => \N__9827\,
            in2 => \_gnd_net_\,
            in3 => \N__8560\,
            lcout => \this_vga_signals.d_N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_c2_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011011101"
        )
    port map (
            in0 => \N__10141\,
            in1 => \N__11060\,
            in2 => \_gnd_net_\,
            in3 => \N__9220\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0\,
            ltout => \this_vga_signals.mult1_un61_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9746\,
            in1 => \N__9167\,
            in2 => \N__8282\,
            in3 => \N__9274\,
            lcout => \this_vga_signals.mult1_un75_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__9745\,
            in1 => \N__10142\,
            in2 => \_gnd_net_\,
            in3 => \N__9103\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIT1827_9_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__9403\,
            in1 => \N__9221\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIRETSA_9_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9402\,
            in2 => \_gnd_net_\,
            in3 => \N__9110\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11689\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22211\,
            ce => \N__11590\,
            sr => \N__11561\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_1_5_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12531\,
            in2 => \_gnd_net_\,
            in3 => \N__12419\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_1_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_26_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001100"
        )
    port map (
            in0 => \N__10806\,
            in1 => \N__10680\,
            in2 => \N__8387\,
            in3 => \N__8612\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__8429\,
            in1 => \N__8498\,
            in2 => \N__8588\,
            in3 => \N__9617\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNISQ5DA02_9_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__9381\,
            in1 => \N__8450\,
            in2 => \N__8384\,
            in3 => \N__8456\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_2_i_m2_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000101011010"
        )
    port map (
            in0 => \N__12248\,
            in1 => \N__10807\,
            in2 => \N__12425\,
            in3 => \N__10669\,
            lcout => \this_vga_signals.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__10010\,
            in1 => \N__9911\,
            in2 => \_gnd_net_\,
            in3 => \N__9026\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_ns_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8885\,
            in2 => \N__8363\,
            in3 => \N__8393\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0\,
            ltout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011110000"
        )
    port map (
            in0 => \N__13417\,
            in1 => \N__8444\,
            in2 => \N__8360\,
            in3 => \N__8480\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010001001101"
        )
    port map (
            in0 => \N__13302\,
            in1 => \N__13418\,
            in2 => \N__8357\,
            in3 => \N__8414\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_i1_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIOE1NOK_2_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__8813\,
            in1 => \N__9569\,
            in2 => \N__8459\,
            in3 => \N__8428\,
            lcout => \this_vga_signals.g1_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_11_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111000101100"
        )
    port map (
            in0 => \N__13303\,
            in1 => \N__10484\,
            in2 => \N__13427\,
            in3 => \N__8399\,
            lcout => \this_vga_signals.mult1_un75_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m1_3_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12836\,
            in1 => \N__9027\,
            in2 => \N__12641\,
            in3 => \N__10012\,
            lcout => \this_vga_signals.if_m1_3\,
            ltout => \this_vga_signals.if_m1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001001011"
        )
    port map (
            in0 => \N__12832\,
            in1 => \N__8438\,
            in2 => \N__8432\,
            in3 => \N__8834\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_x1_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__12775\,
            in1 => \N__9999\,
            in2 => \N__13426\,
            in3 => \N__9894\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10001\,
            in1 => \N__9020\,
            in2 => \N__9916\,
            in3 => \N__8875\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8465\,
            in2 => \N__8417\,
            in3 => \N__8489\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_i\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_37_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100000001111"
        )
    port map (
            in0 => \N__13419\,
            in1 => \N__8846\,
            in2 => \N__8408\,
            in3 => \N__8405\,
            lcout => \this_vga_signals.if_N_2_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x1_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011101101"
        )
    port map (
            in0 => \N__12590\,
            in1 => \N__12777\,
            in2 => \N__9030\,
            in3 => \N__9998\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10000\,
            in1 => \N__9019\,
            in2 => \N__9915\,
            in3 => \N__8874\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12776\,
            in1 => \N__9997\,
            in2 => \N__9031\,
            in3 => \N__9895\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__11521\,
            in1 => \_gnd_net_\,
            in2 => \N__11393\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.vaddress_6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_1_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10008\,
            in1 => \N__9021\,
            in2 => \N__13247\,
            in3 => \N__9908\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_0_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011111100001"
        )
    port map (
            in0 => \N__9909\,
            in1 => \N__12595\,
            in2 => \N__8483\,
            in3 => \N__12828\,
            lcout => \this_vga_signals.g0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12827\,
            in1 => \N__8935\,
            in2 => \N__12640\,
            in3 => \N__9025\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_m3_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001111111"
        )
    port map (
            in0 => \N__13423\,
            in1 => \N__8479\,
            in2 => \N__8468\,
            in3 => \N__8828\,
            lcout => \this_vga_signals.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011011101"
        )
    port map (
            in0 => \N__12591\,
            in1 => \N__12818\,
            in2 => \_gnd_net_\,
            in3 => \N__9907\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_12_x0_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111011111"
        )
    port map (
            in0 => \N__9906\,
            in1 => \N__12826\,
            in2 => \N__9032\,
            in3 => \N__10009\,
            lcout => \this_vga_signals.g0_12_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_2_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9028\,
            in1 => \N__9602\,
            in2 => \N__12838\,
            in3 => \N__9910\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_3_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000101101"
        )
    port map (
            in0 => \N__8879\,
            in1 => \N__12596\,
            in2 => \N__8600\,
            in3 => \N__8597\,
            lcout => \this_vga_signals.g1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI8OIBA_3_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001001"
        )
    port map (
            in0 => \N__10134\,
            in1 => \N__9184\,
            in2 => \N__9752\,
            in3 => \N__9093\,
            lcout => \this_vga_signals.M_hcounter_q_RNI8OIBAZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010011011011"
        )
    port map (
            in0 => \N__9091\,
            in1 => \N__9735\,
            in2 => \N__10140\,
            in3 => \N__9185\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001100110110"
        )
    port map (
            in0 => \N__10133\,
            in1 => \N__9183\,
            in2 => \N__9751\,
            in3 => \N__9092\,
            lcout => \this_vga_signals.if_N_8_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_9_1_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12600\,
            in2 => \N__12837\,
            in3 => \N__8936\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_12_ns_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8954\,
            in2 => \N__8522\,
            in3 => \N__8519\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_8_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110011001"
        )
    port map (
            in0 => \N__9038\,
            in1 => \N__8513\,
            in2 => \N__8507\,
            in3 => \N__8504\,
            lcout => \this_vga_signals.d_N_3_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNIF77A3_1_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8731\,
            in1 => \N__14261\,
            in2 => \_gnd_net_\,
            in3 => \N__8678\,
            lcout => \this_vga_signals.N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_1_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__14116\,
            in1 => \N__8732\,
            in2 => \N__8717\,
            in3 => \N__8698\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22230\,
            ce => \N__14262\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_0_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8697\,
            in1 => \N__8765\,
            in2 => \_gnd_net_\,
            in3 => \N__14115\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22230\,
            ce => \N__14262\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_RNI9C5I1_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14110\,
            in1 => \N__8693\,
            in2 => \_gnd_net_\,
            in3 => \N__8764\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_pcounter_q_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNII2VA2_0_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8713\,
            in2 => \N__8786\,
            in3 => \N__14260\,
            lcout => \this_vga_signals.N_2_0\,
            ltout => \this_vga_signals.N_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8768\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_pcounter_q_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8746\,
            lcout => \this_vga_signals.M_pcounter_q_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_RNI5GDH2_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__8730\,
            in1 => \N__8712\,
            in2 => \N__8699\,
            in3 => \N__14109\,
            lcout => \this_vga_signals.M_pcounter_q_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIHL0E5_9_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9354\,
            in2 => \_gnd_net_\,
            in3 => \N__9239\,
            lcout => \M_this_vga_signals_address_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIN0FTT_9_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100010000100"
        )
    port map (
            in0 => \N__9164\,
            in1 => \N__9353\,
            in2 => \N__8654\,
            in3 => \N__9275\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_6_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101010101"
        )
    port map (
            in0 => \N__12247\,
            in1 => \_gnd_net_\,
            in2 => \N__12421\,
            in3 => \N__12504\,
            lcout => \this_vga_signals.vaddress_1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_1_6_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__12503\,
            in1 => \N__12409\,
            in2 => \_gnd_net_\,
            in3 => \N__12246\,
            lcout => \this_vga_signals.vaddress_4_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10318\,
            in2 => \_gnd_net_\,
            in3 => \N__9505\,
            lcout => \this_vga_signals.vaddress_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11266\,
            lcout => \this_vga_signals.M_vcounter_q_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22204\,
            ce => \N__11591\,
            sr => \N__11562\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__12953\,
            in1 => \N__10319\,
            in2 => \N__10238\,
            in3 => \N__10269\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__9504\,
            in1 => \_gnd_net_\,
            in2 => \N__8801\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\,
            ltout => \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011011001100"
        )
    port map (
            in0 => \N__9291\,
            in1 => \N__10286\,
            in2 => \N__8798\,
            in3 => \N__9309\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11267\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22204\,
            ce => \N__11591\,
            sr => \N__11562\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9503\,
            in2 => \N__10321\,
            in3 => \N__8795\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_1_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNITEVS_6_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111101111"
        )
    port map (
            in0 => \N__10234\,
            in1 => \N__9481\,
            in2 => \N__8789\,
            in3 => \N__12952\,
            lcout => \this_vga_signals.SUM_2_i_1_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11693\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22204\,
            ce => \N__11591\,
            sr => \N__11562\
        );

    \this_vga_signals.un5_vaddress_g0_35_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011010010001"
        )
    port map (
            in0 => \N__10643\,
            in1 => \N__8920\,
            in2 => \N__10791\,
            in3 => \N__11729\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_1_1_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010110001"
        )
    port map (
            in0 => \N__11379\,
            in1 => \N__10400\,
            in2 => \N__12249\,
            in3 => \N__10642\,
            lcout => \this_vga_signals.g1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_14_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010010011001"
        )
    port map (
            in0 => \N__10187\,
            in1 => \N__10756\,
            in2 => \N__10202\,
            in3 => \N__10641\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100000100101"
        )
    port map (
            in0 => \N__10639\,
            in1 => \N__9558\,
            in2 => \N__10790\,
            in3 => \N__11424\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i\,
            ltout => \this_vga_signals.mult1_un54_sum_axb2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_23_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__12648\,
            in1 => \N__8822\,
            in2 => \N__8816\,
            in3 => \N__10452\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m2_1_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010000011001"
        )
    port map (
            in0 => \N__10638\,
            in1 => \N__9557\,
            in2 => \N__10789\,
            in3 => \N__11423\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010000"
        )
    port map (
            in0 => \N__11422\,
            in1 => \N__10755\,
            in2 => \N__9560\,
            in3 => \N__10640\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001001101"
        )
    port map (
            in0 => \N__11391\,
            in1 => \N__12769\,
            in2 => \N__10454\,
            in3 => \N__10522\,
            lcout => \this_vga_signals.mult1_un61_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_395_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010010100101"
        )
    port map (
            in0 => \N__8807\,
            in1 => \N__11389\,
            in2 => \N__9601\,
            in3 => \N__8873\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_395\,
            ltout => \this_vga_signals.mult1_un68_sum_axb1_395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x0_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12618\,
            in1 => \N__12773\,
            in2 => \N__8888\,
            in3 => \N__9005\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__9592\,
            in1 => \N__11390\,
            in2 => \N__10453\,
            in3 => \N__8872\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_1\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_2_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9596\,
            in1 => \N__12774\,
            in2 => \N__8852\,
            in3 => \N__9006\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_5_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100000100100"
        )
    port map (
            in0 => \N__9007\,
            in1 => \N__9512\,
            in2 => \N__8849\,
            in3 => \N__8903\,
            lcout => \this_vga_signals.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_ns_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8840\,
            in1 => \N__9947\,
            in2 => \_gnd_net_\,
            in3 => \N__9008\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_17_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101001010001"
        )
    port map (
            in0 => \N__10523\,
            in1 => \N__10449\,
            in2 => \N__12816\,
            in3 => \N__12617\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12619\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12400\,
            lcout => \this_vga_signals.vaddress_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_29_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10006\,
            in2 => \N__9029\,
            in3 => \N__9902\,
            lcout => \this_vga_signals.N_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101010101"
        )
    port map (
            in0 => \N__12253\,
            in1 => \_gnd_net_\,
            in2 => \N__12646\,
            in3 => \N__12401\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_9_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100011000011"
        )
    port map (
            in0 => \N__10810\,
            in1 => \N__9047\,
            in2 => \N__9041\,
            in3 => \N__9332\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_12_x1_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__10007\,
            in1 => \N__12819\,
            in2 => \N__9917\,
            in3 => \N__9012\,
            lcout => \this_vga_signals.g0_12_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_2_1_0_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010101011010"
        )
    port map (
            in0 => \N__11387\,
            in1 => \N__10809\,
            in2 => \N__12257\,
            in3 => \N__10671\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_2_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101111100100"
        )
    port map (
            in0 => \N__12399\,
            in1 => \N__11388\,
            in2 => \N__8948\,
            in3 => \N__8945\,
            lcout => \this_vga_signals.g0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100001000"
        )
    port map (
            in0 => \N__11122\,
            in1 => \N__9235\,
            in2 => \N__11057\,
            in3 => \N__9121\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_2_9_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__10909\,
            in1 => \N__11175\,
            in2 => \N__11132\,
            in3 => \N__10974\,
            lcout => \this_vga_signals.N_236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010011000011"
        )
    port map (
            in0 => \N__11727\,
            in1 => \N__10808\,
            in2 => \N__8924\,
            in3 => \N__10670\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axb2_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_0_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12645\,
            in2 => \N__8906\,
            in3 => \N__12817\,
            lcout => \this_vga_signals.g0_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_0_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__11123\,
            in1 => \N__8894\,
            in2 => \N__11058\,
            in3 => \N__9422\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_2_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9207\,
            in2 => \N__9278\,
            in3 => \N__9087\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111010000111"
        )
    port map (
            in0 => \N__10972\,
            in1 => \N__11173\,
            in2 => \N__11128\,
            in3 => \N__10907\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010101010111"
        )
    port map (
            in0 => \N__10906\,
            in1 => \N__11107\,
            in2 => \N__11186\,
            in3 => \N__10971\,
            lcout => \this_vga_signals.N_3_2_1\,
            ltout => \this_vga_signals.N_3_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100010000000"
        )
    port map (
            in0 => \N__11027\,
            in1 => \N__10109\,
            in2 => \N__9224\,
            in3 => \N__11121\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__9206\,
            in1 => \_gnd_net_\,
            in2 => \N__10129\,
            in3 => \N__11028\,
            lcout => \this_vga_signals.mult1_un68_sum_axb2_1\,
            ltout => \this_vga_signals.mult1_un68_sum_axb2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001101"
        )
    port map (
            in0 => \N__9703\,
            in1 => \N__10113\,
            in2 => \N__9170\,
            in3 => \N__9086\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__9053\,
            in1 => \N__9131\,
            in2 => \N__9125\,
            in3 => \N__9410\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111000000000"
        )
    port map (
            in0 => \N__11106\,
            in1 => \N__11169\,
            in2 => \N__10983\,
            in3 => \N__10905\,
            lcout => \this_vga_signals.SUM_3_i_0_0_3\,
            ltout => \this_vga_signals.SUM_3_i_0_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_0_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11111\,
            in2 => \N__9056\,
            in3 => \N__11026\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001101"
        )
    port map (
            in0 => \N__11191\,
            in1 => \N__10982\,
            in2 => \N__10928\,
            in3 => \_gnd_net_\,
            lcout => this_vga_signals_hvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110100011"
        )
    port map (
            in0 => \N__11129\,
            in1 => \N__10123\,
            in2 => \N__11059\,
            in3 => \N__9421\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIE00C4_9_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__10988\,
            in1 => \N__10927\,
            in2 => \N__10047\,
            in3 => \N__11187\,
            lcout => \M_this_vga_ramdac_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_7_1_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010010101"
        )
    port map (
            in0 => \N__12023\,
            in1 => \N__12413\,
            in2 => \N__12609\,
            in3 => \N__12254\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_7_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_13_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__9320\,
            in1 => \N__9293\,
            in2 => \N__9335\,
            in3 => \N__9311\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__9319\,
            in1 => \N__9292\,
            in2 => \N__10331\,
            in3 => \N__9310\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_axb1_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_25_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100101001001"
        )
    port map (
            in0 => \N__11656\,
            in1 => \N__10349\,
            in2 => \N__9296\,
            in3 => \N__10779\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIVA761_6_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011110101111"
        )
    port map (
            in0 => \N__10230\,
            in1 => \N__10273\,
            in2 => \N__12964\,
            in3 => \N__9480\,
            lcout => \this_vga_signals.SUM_2_i_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11756\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22202\,
            ce => \N__11593\,
            sr => \N__11560\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11237\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22202\,
            ce => \N__11593\,
            sr => \N__11560\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100101010"
        )
    port map (
            in0 => \N__10388\,
            in1 => \N__12957\,
            in2 => \N__10277\,
            in3 => \N__10231\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10320\,
            in1 => \N__9506\,
            in2 => \N__9485\,
            in3 => \N__9464\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000010111"
        )
    port map (
            in0 => \N__12958\,
            in1 => \N__10270\,
            in2 => \N__9455\,
            in3 => \N__10232\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011010000"
        )
    port map (
            in0 => \N__9452\,
            in1 => \N__11769\,
            in2 => \N__9446\,
            in3 => \N__10389\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11626\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22202\,
            ce => \N__11593\,
            sr => \N__11560\
        );

    \this_vga_signals.un5_vaddress_g0_24_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010100101"
        )
    port map (
            in0 => \N__10765\,
            in1 => \N__10342\,
            in2 => \N__11657\,
            in3 => \N__10646\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_34_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000101001001"
        )
    port map (
            in0 => \N__10647\,
            in1 => \N__10817\,
            in2 => \N__10826\,
            in3 => \N__10766\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__11508\,
            in1 => \N__11453\,
            in2 => \_gnd_net_\,
            in3 => \N__10391\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => \this_vga_signals.vaddress_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010100"
        )
    port map (
            in0 => \N__10837\,
            in1 => \N__11426\,
            in2 => \N__9605\,
            in3 => \N__10760\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_19_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10764\,
            in1 => \N__10392\,
            in2 => \N__11520\,
            in3 => \N__10645\,
            lcout => \this_vga_signals.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIPQ6L81_2_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10474\,
            in1 => \N__10568\,
            in2 => \N__12881\,
            in3 => \N__9600\,
            lcout => \this_vga_signals.g1_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_N_2L1_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010011001"
        )
    port map (
            in0 => \N__9559\,
            in1 => \N__11425\,
            in2 => \N__10792\,
            in3 => \N__10644\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_32_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000110"
        )
    port map (
            in0 => \N__10648\,
            in1 => \N__9539\,
            in2 => \N__9530\,
            in3 => \N__10767\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_2_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12610\,
            in2 => \_gnd_net_\,
            in3 => \N__12361\,
            lcout => \this_vga_signals.vaddress_5_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110101010"
        )
    port map (
            in0 => \N__10673\,
            in1 => \_gnd_net_\,
            in2 => \N__10811\,
            in3 => \N__10561\,
            lcout => \this_vga_signals.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_0_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110101010"
        )
    port map (
            in0 => \N__11728\,
            in1 => \N__10801\,
            in2 => \_gnd_net_\,
            in3 => \N__10672\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_4_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001101111"
        )
    port map (
            in0 => \N__12362\,
            in1 => \N__12623\,
            in2 => \N__9521\,
            in3 => \N__9518\,
            lcout => \this_vga_signals.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_15_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__9941\,
            in1 => \N__10011\,
            in2 => \_gnd_net_\,
            in3 => \N__9912\,
            lcout => \this_vga_signals.N_5_i_5\,
            ltout => \this_vga_signals.N_5_i_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x2_0_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13401\,
            in1 => \N__9668\,
            in2 => \N__9659\,
            in3 => \N__9833\,
            lcout => \this_vga_signals.g0_i_x2_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_1_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001010100"
        )
    port map (
            in0 => \N__9656\,
            in1 => \N__11392\,
            in2 => \N__11525\,
            in3 => \N__9650\,
            lcout => \this_vga_signals.g1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_31_1_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101001"
        )
    port map (
            in0 => \N__12793\,
            in1 => \N__9644\,
            in2 => \N__12644\,
            in3 => \N__10524\,
            lcout => \this_vga_signals.g0_31_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_x0_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110111010111"
        )
    port map (
            in0 => \N__13403\,
            in1 => \N__12809\,
            in2 => \N__9914\,
            in3 => \N__9937\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_2_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_ns_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__10005\,
            in1 => \_gnd_net_\,
            in2 => \N__9638\,
            in3 => \N__9923\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011010101"
        )
    port map (
            in0 => \N__10499\,
            in1 => \N__12810\,
            in2 => \N__9635\,
            in3 => \N__9632\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_0_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001100000"
        )
    port map (
            in0 => \N__13301\,
            in1 => \N__12866\,
            in2 => \N__9626\,
            in3 => \N__9623\,
            lcout => \this_vga_signals.if_i4_mux_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__12122\,
            in1 => \N__12625\,
            in2 => \N__12408\,
            in3 => \N__12965\,
            lcout => \this_vga_signals.vsync_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_x0_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__12806\,
            in1 => \N__13404\,
            in2 => \N__10013\,
            in3 => \N__9887\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_1_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_x1_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__13402\,
            in1 => \N__12808\,
            in2 => \N__9913\,
            in3 => \N__9936\,
            lcout => \this_vga_signals.g0_2_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_20_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010111011"
        )
    port map (
            in0 => \N__12807\,
            in1 => \N__12624\,
            in2 => \_gnd_net_\,
            in3 => \N__9886\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11930\,
            in2 => \N__11978\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14267\,
            in1 => \N__9796\,
            in2 => \_gnd_net_\,
            in3 => \N__9770\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__22221\,
            ce => 'H',
            sr => \N__15056\
        );

    \this_vga_signals.M_hcounter_q_3_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14264\,
            in1 => \N__9721\,
            in2 => \_gnd_net_\,
            in3 => \N__9680\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__22221\,
            ce => 'H',
            sr => \N__15056\
        );

    \this_vga_signals.M_hcounter_q_4_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14268\,
            in1 => \N__10122\,
            in2 => \_gnd_net_\,
            in3 => \N__9677\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__22221\,
            ce => 'H',
            sr => \N__15056\
        );

    \this_vga_signals.M_hcounter_q_5_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14265\,
            in1 => \N__11048\,
            in2 => \_gnd_net_\,
            in3 => \N__9674\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__22221\,
            ce => 'H',
            sr => \N__15056\
        );

    \this_vga_signals.M_hcounter_q_6_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14269\,
            in1 => \N__11127\,
            in2 => \_gnd_net_\,
            in3 => \N__9671\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__22221\,
            ce => 'H',
            sr => \N__15056\
        );

    \this_vga_signals.M_hcounter_q_7_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14266\,
            in1 => \N__11182\,
            in2 => \_gnd_net_\,
            in3 => \N__10175\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__22221\,
            ce => 'H',
            sr => \N__15056\
        );

    \this_vga_signals.M_hcounter_q_8_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14270\,
            in1 => \N__10919\,
            in2 => \_gnd_net_\,
            in3 => \N__10172\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__22221\,
            ce => 'H',
            sr => \N__15056\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10981\,
            in2 => \_gnd_net_\,
            in3 => \N__10169\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22223\,
            ce => \N__10865\,
            sr => \N__15048\
        );

    \this_vga_signals.M_hcounter_q_RNIC1AR_5_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11130\,
            in1 => \N__10127\,
            in2 => \_gnd_net_\,
            in3 => \N__11055\,
            lcout => OPEN,
            ltout => \this_vga_signals.un4_hsynclt8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIMBHF2_9_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__10987\,
            in1 => \N__10067\,
            in2 => \N__10166\,
            in3 => \N__10923\,
            lcout => this_vga_signals_hsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIIED41_7_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__10128\,
            in1 => \N__11056\,
            in2 => \N__11192\,
            in3 => \N__11131\,
            lcout => \this_vga_signals.un3_hsynclt8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIROQM_8_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12019\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12118\,
            lcout => OPEN,
            ltout => \this_vga_signals.un6_vvisibilitylto8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__12219\,
            in1 => \N__12545\,
            in2 => \N__10061\,
            in3 => \N__12414\,
            lcout => \this_vga_signals.un6_vvisibilitylt9_0\,
            ltout => \this_vga_signals.un6_vvisibilitylt9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_9_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__11806\,
            in1 => \N__11776\,
            in2 => \N__10058\,
            in3 => \N__12949\,
            lcout => \this_vga_signals.vvisibility\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11260\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22189\,
            ce => \N__11592\,
            sr => \N__11556\
        );

    \this_vga_signals.un5_vaddress_g0_7_0_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000111000011"
        )
    port map (
            in0 => \N__11519\,
            in1 => \N__12218\,
            in2 => \N__12038\,
            in3 => \N__11380\,
            lcout => \this_vga_signals.g0_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000010011"
        )
    port map (
            in0 => \N__11448\,
            in1 => \N__10386\,
            in2 => \N__10322\,
            in3 => \N__10271\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11681\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22194\,
            ce => \N__11594\,
            sr => \N__11558\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11748\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22194\,
            ce => \N__11594\,
            sr => \N__11558\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110110110111"
        )
    port map (
            in0 => \N__10272\,
            in1 => \N__10233\,
            in2 => \N__12962\,
            in3 => \N__10390\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m8_0_a3_1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__11449\,
            in1 => \_gnd_net_\,
            in2 => \N__10241\,
            in3 => \N__11489\,
            lcout => \this_vga_signals.if_N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11232\,
            lcout => \this_vga_signals.M_vcounter_q_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22194\,
            ce => \N__11594\,
            sr => \N__11558\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_0_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__11451\,
            in1 => \N__10387\,
            in2 => \_gnd_net_\,
            in3 => \N__11491\,
            lcout => \this_vga_signals.vaddress_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_0_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11490\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11450\,
            lcout => \this_vga_signals.vaddress_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_22_1_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111000110"
        )
    port map (
            in0 => \N__10415\,
            in1 => \N__12812\,
            in2 => \N__12643\,
            in3 => \N__10493\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_22_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_22_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10460\,
            in1 => \N__10406\,
            in2 => \N__10487\,
            in3 => \N__10475\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000101011"
        )
    port map (
            in0 => \N__12811\,
            in1 => \N__10451\,
            in2 => \N__12642\,
            in3 => \N__10528\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_0_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11340\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12386\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_5_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_38_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001010000101"
        )
    port map (
            in0 => \N__10681\,
            in1 => \N__11288\,
            in2 => \N__10463\,
            in3 => \N__10783\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i_1\,
            ltout => \this_vga_signals.mult1_un54_sum_axb2_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_36_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010101010"
        )
    port map (
            in0 => \N__10450\,
            in1 => \N__12602\,
            in2 => \N__10418\,
            in3 => \N__10414\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIC07L_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__11512\,
            in1 => \N__11338\,
            in2 => \_gnd_net_\,
            in3 => \N__10393\,
            lcout => \this_vga_signals.vaddress_2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_1_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111011100111"
        )
    port map (
            in0 => \N__11339\,
            in1 => \N__12385\,
            in2 => \N__12255\,
            in3 => \N__10773\,
            lcout => \this_vga_signals.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100101011"
        )
    port map (
            in0 => \N__12728\,
            in1 => \N__10847\,
            in2 => \N__12649\,
            in3 => \N__10841\,
            lcout => \this_vga_signals.g1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12338\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11359\,
            lcout => \this_vga_signals.vaddress_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_0_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__11358\,
            in1 => \N__12339\,
            in2 => \_gnd_net_\,
            in3 => \N__12209\,
            lcout => \this_vga_signals.vaddress_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_1_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12341\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11357\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010100101"
        )
    port map (
            in0 => \N__10562\,
            in1 => \N__10805\,
            in2 => \N__10685\,
            in3 => \N__10682\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011011001111"
        )
    port map (
            in0 => \N__12342\,
            in1 => \N__12635\,
            in2 => \N__10577\,
            in3 => \N__10574\,
            lcout => \this_vga_signals.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__11356\,
            in1 => \N__12340\,
            in2 => \_gnd_net_\,
            in3 => \N__12210\,
            lcout => \this_vga_signals.vaddress_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11630\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22212\,
            ce => \N__11597\,
            sr => \N__11563\
        );

    \this_vga_signals.un5_vaddress_g0_31_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101001"
        )
    port map (
            in0 => \N__10550\,
            in1 => \N__10544\,
            in2 => \N__10538\,
            in3 => \N__10529\,
            lcout => \this_vga_signals.N_5_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__10859\,
            in1 => \N__11216\,
            in2 => \N__12256\,
            in3 => \N__10871\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11174\,
            in2 => \_gnd_net_\,
            in3 => \N__11120\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hcounter_d7lto7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI704B1_9_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__11047\,
            in1 => \N__10973\,
            in2 => \N__10931\,
            in3 => \N__10908\,
            lcout => \this_vga_signals.M_hcounter_d7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010101"
        )
    port map (
            in0 => \N__12650\,
            in1 => \N__13424\,
            in2 => \N__12839\,
            in3 => \N__13304\,
            lcout => \this_vga_signals.un2_vsynclt8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14239\,
            in2 => \_gnd_net_\,
            in3 => \N__15047\,
            lcout => \this_vga_signals.N_340_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13425\,
            in2 => \_gnd_net_\,
            in3 => \N__12047\,
            lcout => \this_vga_signals.vsync_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14256\,
            in1 => \N__12862\,
            in2 => \N__14120\,
            in3 => \N__14114\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__22183\,
            ce => 'H',
            sr => \N__11555\
        );

    \this_vga_signals.M_vcounter_q_1_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14258\,
            in1 => \N__13285\,
            in2 => \_gnd_net_\,
            in3 => \N__10853\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__22183\,
            ce => 'H',
            sr => \N__11555\
        );

    \this_vga_signals.M_vcounter_q_2_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14257\,
            in1 => \N__13363\,
            in2 => \_gnd_net_\,
            in3 => \N__10850\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__22183\,
            ce => 'H',
            sr => \N__11555\
        );

    \this_vga_signals.M_vcounter_q_3_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14259\,
            in1 => \N__12710\,
            in2 => \_gnd_net_\,
            in3 => \N__11279\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__22183\,
            ce => 'H',
            sr => \N__11555\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12639\,
            in2 => \_gnd_net_\,
            in3 => \N__11276\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12418\,
            in2 => \_gnd_net_\,
            in3 => \N__11273\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12242\,
            in2 => \_gnd_net_\,
            in3 => \N__11270\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12046\,
            in2 => \_gnd_net_\,
            in3 => \N__11246\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12112\,
            in2 => \_gnd_net_\,
            in3 => \N__11243\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12951\,
            in2 => \_gnd_net_\,
            in3 => \N__11240\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22190\,
            ce => \N__11595\,
            sr => \N__11557\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_8_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12039\,
            in1 => \N__12948\,
            in2 => \N__12117\,
            in3 => \N__12184\,
            lcout => \this_vga_signals.vaddress_ac0_9_0_a0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11233\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22195\,
            ce => \N__11596\,
            sr => \N__11559\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11752\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22195\,
            ce => \N__11596\,
            sr => \N__11559\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__12183\,
            in1 => \N__11342\,
            in2 => \_gnd_net_\,
            in3 => \N__11488\,
            lcout => \this_vga_signals.vaddress_5_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11688\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22195\,
            ce => \N__11596\,
            sr => \N__11559\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_0_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11341\,
            in2 => \_gnd_net_\,
            in3 => \N__11487\,
            lcout => \this_vga_signals.vaddress_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11614\,
            lcout => \this_vga_signals.M_vcounter_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22195\,
            ce => \N__11596\,
            sr => \N__11559\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11486\,
            in2 => \_gnd_net_\,
            in3 => \N__11452\,
            lcout => \this_vga_signals.vaddress_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_1_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101010101"
        )
    port map (
            in0 => \N__12186\,
            in1 => \_gnd_net_\,
            in2 => \N__12379\,
            in3 => \N__11360\,
            lcout => \this_vga_signals.vaddress_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_0_8_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12048\,
            in1 => \N__12334\,
            in2 => \N__12116\,
            in3 => \N__12185\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_d7lto8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__12278\,
            in1 => \N__12601\,
            in2 => \N__11282\,
            in3 => \N__12963\,
            lcout => \this_vga_signals.M_vcounter_d8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11964\,
            in1 => \N__11900\,
            in2 => \_gnd_net_\,
            in3 => \N__14231\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22205\,
            ce => 'H',
            sr => \N__15037\
        );

    \this_delay_clk.M_pipe_q_4_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11861\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.out_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__11854\,
            in1 => \_gnd_net_\,
            in2 => \N__11819\,
            in3 => \N__11841\,
            lcout => \M_this_start_address_delay_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11876\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBJQQ_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__11843\,
            in1 => \N__11815\,
            in2 => \_gnd_net_\,
            in3 => \N__11853\,
            lcout => \M_this_start_data_delay_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11855\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11842\,
            lcout => \this_start_data_delay_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIQ80L_2_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20922\,
            in1 => \N__16213\,
            in2 => \_gnd_net_\,
            in3 => \N__20388\,
            lcout => port_dmab_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIBILS3_6_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__11807\,
            in1 => \N__11789\,
            in2 => \N__13208\,
            in3 => \N__11780\,
            lcout => \M_this_ppu_vga_is_drawing_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14336\,
            in1 => \N__14366\,
            in2 => \_gnd_net_\,
            in3 => \N__12950\,
            lcout => \this_vga_signals.line_clk_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIV19S_2_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12681\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13339\,
            lcout => \this_vga_signals.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__13272\,
            in1 => \N__12852\,
            in2 => \N__13364\,
            in3 => \N__12680\,
            lcout => \this_vga_signals.M_vcounter_d7lt8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110111"
        )
    port map (
            in0 => \N__12647\,
            in1 => \N__12420\,
            in2 => \N__12277\,
            in3 => \N__12211\,
            lcout => \this_vga_signals.un4_lvisibility_1\,
            ltout => \this_vga_signals.un4_lvisibility_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICHRV3_8_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010001010"
        )
    port map (
            in0 => \N__12067\,
            in1 => \N__12110\,
            in2 => \N__12125\,
            in3 => \N__12049\,
            lcout => \M_this_vga_signals_line_clk_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010010001100"
        )
    port map (
            in0 => \N__12111\,
            in1 => \N__12068\,
            in2 => \N__12059\,
            in3 => \N__12050\,
            lcout => \this_ppu.line_clk.M_last_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_0_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11963\,
            in2 => \_gnd_net_\,
            in3 => \N__14235\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22196\,
            ce => 'H',
            sr => \N__15055\
        );

    \M_this_sprites_address_q_RNO_0_5_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100110011"
        )
    port map (
            in0 => \N__16418\,
            in1 => \N__13635\,
            in2 => \N__21472\,
            in3 => \N__20255\,
            lcout => \M_this_sprites_address_q_3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_3_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13400\,
            in2 => \_gnd_net_\,
            in3 => \N__13300\,
            lcout => \this_vga_signals.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_4_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100110011"
        )
    port map (
            in0 => \N__16417\,
            in1 => \N__13770\,
            in2 => \N__20120\,
            in3 => \N__20254\,
            lcout => \M_this_sprites_address_q_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_2_4_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__21992\,
            in1 => \N__13173\,
            in2 => \N__22447\,
            in3 => \N__20256\,
            lcout => OPEN,
            ltout => \N_206_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__13223\,
            in1 => \N__13229\,
            in2 => \N__13232\,
            in3 => \N__14417\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22206\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_3_4_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21993\,
            in1 => \N__16277\,
            in2 => \_gnd_net_\,
            in3 => \N__16217\,
            lcout => \N_207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_0_4_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__14407\,
            in1 => \N__20377\,
            in2 => \N__20975\,
            in3 => \N__21991\,
            lcout => \M_this_state_q_srsts_0_a2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIQ80L_0_2_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__13174\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => port_dmab_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_0_2_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__16214\,
            in1 => \N__20389\,
            in2 => \N__16249\,
            in3 => \N__21995\,
            lcout => \M_this_state_q_srsts_i_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_3_ns_1_11_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__16411\,
            in1 => \N__21016\,
            in2 => \N__20119\,
            in3 => \N__20290\,
            lcout => \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNI5CEE4_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15101\,
            in2 => \_gnd_net_\,
            in3 => \N__15137\,
            lcout => \this_ppu.M_line_clk_out_0\,
            ltout => \this_ppu.M_line_clk_out_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIDFVT8_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__19368\,
            in1 => \N__13460\,
            in2 => \N__13454\,
            in3 => \N__21990\,
            lcout => \this_ppu.N_258_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_5_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__17512\,
            in1 => \N__13451\,
            in2 => \N__22420\,
            in3 => \N__13616\,
            lcout => \M_this_sprites_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22197\,
            ce => 'H',
            sr => \N__21941\
        );

    \M_this_sprites_address_q_4_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__17511\,
            in1 => \N__13445\,
            in2 => \N__22419\,
            in3 => \N__13751\,
            lcout => \M_this_sprites_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22197\,
            ce => 'H',
            sr => \N__21941\
        );

    \M_this_sprites_address_q_RNO_0_7_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__16415\,
            in1 => \N__13503\,
            in2 => \N__20163\,
            in3 => \N__20335\,
            lcout => OPEN,
            ltout => \M_this_sprites_address_q_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_7_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001110100001100"
        )
    port map (
            in0 => \N__22365\,
            in1 => \N__17513\,
            in2 => \N__13439\,
            in3 => \N__13484\,
            lcout => \M_this_sprites_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22197\,
            ce => 'H',
            sr => \N__21941\
        );

    \M_this_sprites_address_q_RNO_1_0_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15283\,
            in2 => \N__14387\,
            in3 => \N__14386\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_1_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14569\,
            in2 => \_gnd_net_\,
            in3 => \N__13436\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_0\,
            carryout => \un1_M_this_sprites_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_2_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16716\,
            in2 => \_gnd_net_\,
            in3 => \N__13433\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_1\,
            carryout => \un1_M_this_sprites_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_3_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17323\,
            in2 => \_gnd_net_\,
            in3 => \N__13430\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_2\,
            carryout => \un1_M_this_sprites_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_4_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13771\,
            in2 => \_gnd_net_\,
            in3 => \N__13745\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_3\,
            carryout => \un1_M_this_sprites_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_5_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13636\,
            in2 => \_gnd_net_\,
            in3 => \N__13610\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_4\,
            carryout => \un1_M_this_sprites_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_6_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14830\,
            in2 => \_gnd_net_\,
            in3 => \N__13607\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_5\,
            carryout => \un1_M_this_sprites_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_7_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13504\,
            in2 => \_gnd_net_\,
            in3 => \N__13478\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_6\,
            carryout => \un1_M_this_sprites_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_8_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13924\,
            in2 => \_gnd_net_\,
            in3 => \N__13475\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_9_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14704\,
            in2 => \_gnd_net_\,
            in3 => \N__13472\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_8\,
            carryout => \un1_M_this_sprites_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_10_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16444\,
            in2 => \_gnd_net_\,
            in3 => \N__13469\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_9\,
            carryout => \un1_M_this_sprites_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21015\,
            in2 => \_gnd_net_\,
            in3 => \N__13466\,
            lcout => \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_10\,
            carryout => \un1_M_this_sprites_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21281\,
            in2 => \_gnd_net_\,
            in3 => \N__13463\,
            lcout => \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_11\,
            carryout => \un1_M_this_sprites_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21092\,
            in2 => \_gnd_net_\,
            in3 => \N__14042\,
            lcout => \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_3_ns_1_12_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001111111"
        )
    port map (
            in0 => \N__20325\,
            in1 => \N__16413\,
            in2 => \N__21473\,
            in3 => \N__21282\,
            lcout => \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_8_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__16414\,
            in1 => \N__13923\,
            in2 => \N__21542\,
            in3 => \N__20331\,
            lcout => OPEN,
            ltout => \M_this_sprites_address_q_3_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_8_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101001001110"
        )
    port map (
            in0 => \N__17509\,
            in1 => \N__14039\,
            in2 => \N__14033\,
            in3 => \N__22422\,
            lcout => \M_this_sprites_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22214\,
            ce => 'H',
            sr => \N__21940\
        );

    \M_this_sprites_address_q_11_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__17507\,
            in1 => \N__13904\,
            in2 => \N__22448\,
            in3 => \N__13898\,
            lcout => \M_this_sprites_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22214\,
            ce => 'H',
            sr => \N__21940\
        );

    \M_this_sprites_address_q_12_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__17508\,
            in1 => \N__13892\,
            in2 => \N__22449\,
            in3 => \N__13886\,
            lcout => \M_this_sprites_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22214\,
            ce => 'H',
            sr => \N__21940\
        );

    \M_this_sprites_address_q_1_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__17510\,
            in1 => \N__14543\,
            in2 => \N__22450\,
            in3 => \N__13880\,
            lcout => \M_this_sprites_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22217\,
            ce => 'H',
            sr => \N__21937\
        );

    \this_vga_signals.M_lcounter_q_RNIGRI95_1_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__14334\,
            in1 => \N__15077\,
            in2 => \_gnd_net_\,
            in3 => \N__14118\,
            lcout => \this_vga_signals.un1_M_hcounter_d7_1_0\,
            ltout => \this_vga_signals.un1_M_hcounter_d7_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_0_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011011001100"
        )
    port map (
            in0 => \N__14119\,
            in1 => \N__14365\,
            in2 => \N__13871\,
            in3 => \N__14205\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_1_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14364\,
            in2 => \_gnd_net_\,
            in3 => \N__14117\,
            lcout => OPEN,
            ltout => \this_vga_signals.CO0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_1_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011101000000"
        )
    port map (
            in0 => \N__14345\,
            in1 => \N__14204\,
            in2 => \N__14339\,
            in3 => \N__14335\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_0_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010011000000000"
        )
    port map (
            in0 => \N__17943\,
            in1 => \N__14318\,
            in2 => \N__19385\,
            in3 => \N__16863\,
            lcout => \M_this_ppu_vram_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14304\,
            in2 => \_gnd_net_\,
            in3 => \N__14312\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14303\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__14306\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14276\,
            lcout => \M_this_state_q_nss_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14305\,
            in2 => \_gnd_net_\,
            in3 => \N__14282\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_RNIFKS8_1_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__14473\,
            in1 => \N__14964\,
            in2 => \_gnd_net_\,
            in3 => \N__21987\,
            lcout => \M_counter_q_RNIFKS8_1\,
            ltout => \M_counter_q_RNIFKS8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIMK0K1_9_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14123\,
            in3 => \N__14101\,
            lcout => \this_vga_signals.M_vcounter_q_249_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_0_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14501\,
            lcout => \M_this_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22188\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_1_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__14474\,
            in1 => \N__14965\,
            in2 => \_gnd_net_\,
            in3 => \N__21988\,
            lcout => \this_pixel_clk.M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22188\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_2_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001110000"
        )
    port map (
            in0 => \N__16216\,
            in1 => \N__16276\,
            in2 => \N__14465\,
            in3 => \N__20289\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_6_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011011111"
        )
    port map (
            in0 => \N__20288\,
            in1 => \N__16386\,
            in2 => \N__19796\,
            in3 => \N__14829\,
            lcout => \M_this_sprites_address_q_3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_rw_iobuf_RNIILOC1_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__14406\,
            in1 => \N__16248\,
            in2 => \N__14450\,
            in3 => \N__21989\,
            lcout => \N_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_4_4_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__14446\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16247\,
            lcout => OPEN,
            ltout => \N_171_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_1_4_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__21764\,
            in1 => \N__16019\,
            in2 => \N__14420\,
            in3 => \N__16045\,
            lcout => \N_176_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI95RM1_4_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__16215\,
            in1 => \N__19169\,
            in2 => \N__14408\,
            in3 => \N__20287\,
            lcout => \N_153_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_2_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__17494\,
            in1 => \N__22427\,
            in2 => \N__16694\,
            in3 => \N__14372\,
            lcout => \M_this_sprites_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22201\,
            ce => 'H',
            sr => \N__21939\
        );

    \M_this_sprites_address_q_9_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__17495\,
            in1 => \N__22428\,
            in2 => \N__14684\,
            in3 => \N__14951\,
            lcout => \M_this_sprites_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22201\,
            ce => 'H',
            sr => \N__21939\
        );

    \M_this_sprites_address_q_13_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__17482\,
            in1 => \N__16826\,
            in2 => \N__22452\,
            in3 => \N__14945\,
            lcout => \M_this_sprites_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22201\,
            ce => 'H',
            sr => \N__21939\
        );

    \M_this_sprites_address_q_6_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011101000100"
        )
    port map (
            in0 => \N__14939\,
            in1 => \N__17483\,
            in2 => \N__22453\,
            in3 => \N__14933\,
            lcout => \M_this_sprites_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22201\,
            ce => 'H',
            sr => \N__21939\
        );

    \M_this_state_q_RNI20CE_0_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__22375\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21996\,
            lcout => \M_this_state_q_RNI20CEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_9_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__16410\,
            in1 => \N__14703\,
            in2 => \N__19843\,
            in3 => \N__20327\,
            lcout => \M_this_sprites_address_q_3_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_1_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011011111"
        )
    port map (
            in0 => \N__20326\,
            in1 => \N__16412\,
            in2 => \N__21538\,
            in3 => \N__14562\,
            lcout => \M_this_sprites_address_q_3_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI9PQ_4_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__18585\,
            in1 => \N__17100\,
            in2 => \N__18430\,
            in3 => \N__15155\,
            lcout => \this_ppu.un1_M_line_clk_out_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNO_0_4_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18901\,
            in1 => \N__17026\,
            in2 => \N__17107\,
            in3 => \N__16120\,
            lcout => OPEN,
            ltout => \this_ppu.un1_M_haddress_q_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_4_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101000000000"
        )
    port map (
            in0 => \N__18433\,
            in1 => \N__18586\,
            in2 => \N__14537\,
            in3 => \N__16174\,
            lcout => \M_this_ppu_vram_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNITAF_6_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18265\,
            in1 => \N__17021\,
            in2 => \N__18115\,
            in3 => \N__18900\,
            lcout => \this_ppu.M_haddress_d8lto6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNI5NOQ4_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__19367\,
            in1 => \N__15149\,
            in2 => \N__15116\,
            in3 => \N__15143\,
            lcout => \this_ppu.M_last_q_RNI5NOQ4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_1_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__17796\,
            in1 => \N__16850\,
            in2 => \_gnd_net_\,
            in3 => \N__16072\,
            lcout => \this_ppu.M_vaddress_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIMT2V4_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__17939\,
            in1 => \N__19372\,
            in2 => \N__15114\,
            in3 => \N__15138\,
            lcout => \this_ppu.un1_M_vaddress_q_c1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNI2T915_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__19373\,
            in1 => \N__15139\,
            in2 => \N__15115\,
            in3 => \N__21994\,
            lcout => \this_ppu.N_250_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIRO2H5_9_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15073\,
            in2 => \_gnd_net_\,
            in3 => \N__15019\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNIRO2H5Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_0_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__17506\,
            in1 => \N__15251\,
            in2 => \N__22421\,
            in3 => \N__14978\,
            lcout => \M_this_sprites_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22198\,
            ce => 'H',
            sr => \N__21942\
        );

    \this_pixel_clk.M_counter_q_0_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14966\,
            lcout => \this_pixel_clk.M_counter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22198\,
            ce => 'H',
            sr => \N__21942\
        );

    \M_this_data_count_q_RNIBTAK_10_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15187\,
            in1 => \N__15169\,
            in2 => \N__15419\,
            in3 => \N__15205\,
            lcout => \M_this_state_q_srsts_i_a2_1_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_0_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011101010101"
        )
    port map (
            in0 => \N__15270\,
            in1 => \N__16396\,
            in2 => \N__20174\,
            in3 => \N__20281\,
            lcout => \M_this_sprites_address_q_3_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIAVRI_11_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15394\,
            in1 => \N__15439\,
            in2 => \N__15956\,
            in3 => \N__15460\,
            lcout => OPEN,
            ltout => \M_this_state_q_srsts_i_a2_1_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIDFF62_10_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15236\,
            in1 => \N__15245\,
            in2 => \N__15239\,
            in3 => \N__15230\,
            lcout => \N_233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIAQQL_4_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15493\,
            in1 => \N__15511\,
            in2 => \N__15535\,
            in3 => \N__15475\,
            lcout => \M_this_state_q_srsts_i_a2_1_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIEOD9_13_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15220\,
            in2 => \_gnd_net_\,
            in3 => \N__15557\,
            lcout => \M_this_state_q_srsts_i_a2_1_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_0_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20923\,
            in2 => \N__15224\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_23_0_\,
            carryout => \un1_M_this_data_count_q_cry_0\,
            clk => \N__22207\,
            ce => 'H',
            sr => \N__15932\
        );

    \M_this_data_count_q_1_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20927\,
            in2 => \N__15209\,
            in3 => \N__15194\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_0\,
            carryout => \un1_M_this_data_count_q_cry_1\,
            clk => \N__22207\,
            ce => 'H',
            sr => \N__15932\
        );

    \M_this_data_count_q_2_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20924\,
            in2 => \N__15191\,
            in3 => \N__15176\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_1\,
            carryout => \un1_M_this_data_count_q_cry_2\,
            clk => \N__22207\,
            ce => 'H',
            sr => \N__15932\
        );

    \M_this_data_count_q_3_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20928\,
            in2 => \N__15173\,
            in3 => \N__15158\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_2\,
            carryout => \un1_M_this_data_count_q_cry_3\,
            clk => \N__22207\,
            ce => 'H',
            sr => \N__15932\
        );

    \M_this_data_count_q_4_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20925\,
            in2 => \N__15536\,
            in3 => \N__15518\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_3\,
            carryout => \un1_M_this_data_count_q_cry_4\,
            clk => \N__22207\,
            ce => 'H',
            sr => \N__15932\
        );

    \M_this_data_count_q_5_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20929\,
            in2 => \N__15515\,
            in3 => \N__15500\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_4\,
            carryout => \un1_M_this_data_count_q_cry_5\,
            clk => \N__22207\,
            ce => 'H',
            sr => \N__15932\
        );

    \M_this_data_count_q_6_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20926\,
            in2 => \N__15497\,
            in3 => \N__15482\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_5\,
            carryout => \un1_M_this_data_count_q_cry_6\,
            clk => \N__22207\,
            ce => 'H',
            sr => \N__15932\
        );

    \M_this_data_count_q_7_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20930\,
            in2 => \N__15479\,
            in3 => \N__15464\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_6\,
            carryout => \un1_M_this_data_count_q_cry_7\,
            clk => \N__22207\,
            ce => 'H',
            sr => \N__15932\
        );

    \M_this_data_count_q_8_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20958\,
            in2 => \N__15461\,
            in3 => \N__15443\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_24_0_\,
            carryout => \un1_M_this_data_count_q_cry_8\,
            clk => \N__22215\,
            ce => 'H',
            sr => \N__15925\
        );

    \M_this_data_count_q_9_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20961\,
            in2 => \N__15440\,
            in3 => \N__15422\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_8\,
            carryout => \un1_M_this_data_count_q_cry_9\,
            clk => \N__22215\,
            ce => 'H',
            sr => \N__15925\
        );

    \M_this_data_count_q_10_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20959\,
            in2 => \N__15418\,
            in3 => \N__15398\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_9\,
            carryout => \un1_M_this_data_count_q_cry_10\,
            clk => \N__22215\,
            ce => 'H',
            sr => \N__15925\
        );

    \M_this_data_count_q_11_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20962\,
            in2 => \N__15395\,
            in3 => \N__15377\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_10\,
            carryout => \un1_M_this_data_count_q_cry_11\,
            clk => \N__22215\,
            ce => 'H',
            sr => \N__15925\
        );

    \M_this_data_count_q_12_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20960\,
            in2 => \N__15955\,
            in3 => \N__15935\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_11\,
            carryout => \un1_M_this_data_count_q_cry_12\,
            clk => \N__22215\,
            ce => 'H',
            sr => \N__15925\
        );

    \un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15668\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_12\,
            carryout => \un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15670\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO\,
            carryout => \un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15669\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO\,
            carryout => \un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__22435\,
            in1 => \N__15556\,
            in2 => \N__20973\,
            in3 => \N__15560\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22218\,
            ce => 'H',
            sr => \N__21938\
        );

    \this_ppu.M_haddress_q_RNIU60R4_1_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17085\,
            in1 => \N__18903\,
            in2 => \_gnd_net_\,
            in3 => \N__16119\,
            lcout => \this_ppu.un1_M_haddress_q_c2\,
            ltout => \this_ppu.un1_M_haddress_q_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIBMBR4_4_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18432\,
            in1 => \N__18590\,
            in2 => \N__15542\,
            in3 => \N__17025\,
            lcout => \this_ppu.un1_M_haddress_q_c5\,
            ltout => \this_ppu.un1_M_haddress_q_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_6_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__16161\,
            in1 => \N__18114\,
            in2 => \N__15539\,
            in3 => \N__18270\,
            lcout => \M_this_ppu_vram_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_2_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__17027\,
            in1 => \N__16158\,
            in2 => \_gnd_net_\,
            in3 => \N__16081\,
            lcout => \M_this_ppu_vram_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_5_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16159\,
            in1 => \N__18269\,
            in2 => \_gnd_net_\,
            in3 => \N__16088\,
            lcout => \M_this_ppu_vram_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_3_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100010001000"
        )
    port map (
            in0 => \N__18591\,
            in1 => \N__16160\,
            in2 => \N__17035\,
            in3 => \N__16082\,
            lcout => \M_this_ppu_vram_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_4_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100011000000"
        )
    port map (
            in0 => \N__19127\,
            in1 => \N__16865\,
            in2 => \N__18989\,
            in3 => \N__16103\,
            lcout => \this_ppu.M_vaddress_qZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_2_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100011000000"
        )
    port map (
            in0 => \N__17797\,
            in1 => \N__16864\,
            in2 => \N__17654\,
            in3 => \N__16073\,
            lcout => \this_ppu.M_vaddress_qZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNID0D95_2_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17646\,
            in1 => \N__17792\,
            in2 => \_gnd_net_\,
            in3 => \N__16071\,
            lcout => \this_ppu.un1_M_vaddress_q_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_5_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__20286\,
            in1 => \N__15962\,
            in2 => \N__16404\,
            in3 => \N__22000\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_0_7_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__16055\,
            in1 => \N__16018\,
            in2 => \N__21767\,
            in3 => \N__15977\,
            lcout => \N_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_0_6_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16054\,
            in1 => \N__16017\,
            in2 => \N__21766\,
            in3 => \N__15976\,
            lcout => \N_202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_0_5_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16053\,
            in1 => \N__16016\,
            in2 => \N__21765\,
            in3 => \N__15975\,
            lcout => \N_204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_6_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__21999\,
            in1 => \N__16292\,
            in2 => \N__20336\,
            in3 => \N__16286\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIVD0L_6_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__16375\,
            in1 => \N__16285\,
            in2 => \_gnd_net_\,
            in3 => \N__22395\,
            lcout => \M_this_sprites_address_q_3_sm0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNO_0_1_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__16275\,
            in1 => \N__16256\,
            in2 => \_gnd_net_\,
            in3 => \N__16204\,
            lcout => OPEN,
            ltout => \M_this_state_q_srsts_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_1_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__22396\,
            in1 => \N__20952\,
            in2 => \N__16220\,
            in3 => \N__21998\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_1_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000011000000"
        )
    port map (
            in0 => \N__18896\,
            in1 => \N__17086\,
            in2 => \N__16175\,
            in3 => \N__16133\,
            lcout => \M_this_ppu_vram_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_0_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__16132\,
            in1 => \N__16170\,
            in2 => \_gnd_net_\,
            in3 => \N__18895\,
            lcout => \M_this_ppu_vram_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16131\,
            in2 => \_gnd_net_\,
            in3 => \N__21997\,
            lcout => \M_this_ppu_vram_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_6_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010100000"
        )
    port map (
            in0 => \N__16868\,
            in1 => \N__18962\,
            in2 => \N__18941\,
            in3 => \N__16874\,
            lcout => \this_ppu.M_vaddress_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_3_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__19124\,
            in1 => \N__16866\,
            in2 => \_gnd_net_\,
            in3 => \N__16102\,
            lcout => \this_ppu.M_vaddress_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNI87NJ5_4_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18981\,
            in1 => \N__19126\,
            in2 => \_gnd_net_\,
            in3 => \N__16101\,
            lcout => \this_ppu.un1_M_vaddress_q_c5\,
            ltout => \this_ppu.un1_M_vaddress_q_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_5_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16867\,
            in1 => \_gnd_net_\,
            in2 => \N__16829\,
            in3 => \N__18961\,
            lcout => \this_ppu.M_vaddress_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_3_ns_1_13_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110101010101"
        )
    port map (
            in0 => \N__21106\,
            in1 => \N__16371\,
            in2 => \N__19795\,
            in3 => \N__20322\,
            lcout => \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_2_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100110011"
        )
    port map (
            in0 => \N__16385\,
            in1 => \N__16726\,
            in2 => \N__19844\,
            in3 => \N__20321\,
            lcout => \M_this_sprites_address_q_3_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI84774_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__19378\,
            in1 => \N__18617\,
            in2 => \N__19278\,
            in3 => \N__17216\,
            lcout => \M_this_ppu_vram_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIPF7_1_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17081\,
            in2 => \_gnd_net_\,
            in3 => \N__18894\,
            lcout => \M_this_ppu_sprites_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_10_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110101010101"
        )
    port map (
            in0 => \N__16437\,
            in1 => \N__16400\,
            in2 => \N__19985\,
            in3 => \N__20282\,
            lcout => \M_this_sprites_address_q_3_ns_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_10_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__17504\,
            in1 => \N__16556\,
            in2 => \N__22451\,
            in3 => \N__16550\,
            lcout => \M_this_sprites_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22222\,
            ce => 'H',
            sr => \N__21943\
        );

    \M_this_sprites_address_q_RNO_0_3_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001111"
        )
    port map (
            in0 => \N__16416\,
            in1 => \N__19971\,
            in2 => \N__17313\,
            in3 => \N__20323\,
            lcout => OPEN,
            ltout => \M_this_sprites_address_q_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_3_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__17505\,
            in1 => \N__22423\,
            in2 => \N__17432\,
            in3 => \N__17429\,
            lcout => \M_this_sprites_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22222\,
            ce => 'H',
            sr => \N__21943\
        );

    \M_this_state_q_3_LC_20_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20390\,
            in2 => \_gnd_net_\,
            in3 => \N__20324\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22222\,
            ce => 'H',
            sr => \N__21943\
        );

    \this_sprites_ram.mem_mem_1_1_RNIJBQ01_0_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__20495\,
            in1 => \N__17285\,
            in2 => \N__20672\,
            in3 => \N__17267\,
            lcout => \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIDT2Q1_0_LC_21_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__17255\,
            in1 => \N__20530\,
            in2 => \N__17240\,
            in3 => \N__17222\,
            lcout => \this_sprites_ram_mem_N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI04774_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__19374\,
            in1 => \N__18683\,
            in2 => \N__19268\,
            in3 => \N__17156\,
            lcout => \M_this_ppu_vram_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNI5LUP1_0_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__17192\,
            in1 => \N__20546\,
            in2 => \N__17177\,
            in3 => \N__17120\,
            lcout => \this_sprites_ram_mem_N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIF7O01_0_LC_21_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__20496\,
            in1 => \N__17150\,
            in2 => \N__20657\,
            in3 => \N__17138\,
            lcout => \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_cry_1_c_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18902\,
            in2 => \N__17099\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_21_17_0_\,
            carryout => \this_ppu.sprites_addr_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_cry_1_c_RNIB25D_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17031\,
            in2 => \_gnd_net_\,
            in3 => \N__18605\,
            lcout => \M_this_ppu_sprites_addr_2\,
            ltout => OPEN,
            carryin => \this_ppu.sprites_addr_cry_1\,
            carryout => \this_ppu.sprites_addr_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_cry_2_c_RNID56D_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18595\,
            in2 => \_gnd_net_\,
            in3 => \N__18446\,
            lcout => \M_this_ppu_sprites_addr_3\,
            ltout => OPEN,
            carryin => \this_ppu.sprites_addr_cry_2\,
            carryout => \this_ppu.sprites_addr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_cry_3_c_RNIF87D_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18431\,
            in2 => \_gnd_net_\,
            in3 => \N__18284\,
            lcout => \M_this_ppu_sprites_addr_4\,
            ltout => OPEN,
            carryin => \this_ppu.sprites_addr_cry_3\,
            carryout => \this_ppu.sprites_addr_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_cry_4_c_RNIHB8D_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18274\,
            in2 => \_gnd_net_\,
            in3 => \N__18131\,
            lcout => \M_this_ppu_sprites_addr_5\,
            ltout => OPEN,
            carryin => \this_ppu.sprites_addr_cry_4\,
            carryout => \this_ppu.sprites_addr_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_cry_5_c_RNIJE9D_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18113\,
            in2 => \_gnd_net_\,
            in3 => \N__17969\,
            lcout => \M_this_ppu_sprites_addr_6\,
            ltout => OPEN,
            carryin => \this_ppu.sprites_addr_cry_5\,
            carryout => \this_ppu.sprites_addr_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_cry_6_c_RNISIBI_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17959\,
            in2 => \_gnd_net_\,
            in3 => \N__17804\,
            lcout => \M_this_ppu_sprites_addr_7\,
            ltout => OPEN,
            carryin => \this_ppu.sprites_addr_cry_6\,
            carryout => \this_ppu.sprites_addr_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_cry_7_c_RNIULCI_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17801\,
            in2 => \_gnd_net_\,
            in3 => \N__17657\,
            lcout => \M_this_ppu_sprites_addr_8\,
            ltout => OPEN,
            carryin => \this_ppu.sprites_addr_cry_7\,
            carryout => \this_ppu.sprites_addr_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_cry_8_c_RNI0PDI_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17653\,
            in2 => \_gnd_net_\,
            in3 => \N__17516\,
            lcout => \M_this_ppu_sprites_addr_9\,
            ltout => OPEN,
            carryin => \bfn_21_18_0_\,
            carryout => \this_ppu.sprites_addr_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_cry_9_c_RNI2SEI_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19125\,
            in2 => \_gnd_net_\,
            in3 => \N__18992\,
            lcout => \M_this_ppu_sprites_addr_10\,
            ltout => OPEN,
            carryin => \this_ppu.sprites_addr_cry_9\,
            carryout => \this_ppu.sprites_addr_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_11_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18988\,
            in2 => \_gnd_net_\,
            in3 => \N__18965\,
            lcout => this_sprites_ram_mem_radreg_11,
            ltout => OPEN,
            carryin => \this_ppu.sprites_addr_cry_10\,
            carryout => \this_ppu.sprites_addr_cry_11\,
            clk => \N__22203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_12_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18960\,
            in2 => \_gnd_net_\,
            in3 => \N__18944\,
            lcout => \this_sprites_ram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \this_ppu.sprites_addr_cry_11\,
            carryout => \this_ppu.sprites_addr_cry_12\,
            clk => \N__22203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_13_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18937\,
            in2 => \_gnd_net_\,
            in3 => \N__18923\,
            lcout => \this_sprites_ram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNICN3_0_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18910\,
            lcout => \M_this_ppu_vram_addr_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNIHBQ01_0_LC_22_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__20535\,
            in1 => \N__18743\,
            in2 => \N__20683\,
            in3 => \N__18731\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNI9T2Q1_0_LC_22_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__18716\,
            in1 => \N__18695\,
            in2 => \N__18686\,
            in3 => \N__20536\,
            lcout => \this_sprites_ram_mem_N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_wclke_3_LC_22_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21338\,
            in1 => \N__21076\,
            in2 => \N__21183\,
            in3 => \N__21257\,
            lcout => \this_sprites_ram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNI9LUP1_0_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__18647\,
            in1 => \N__20534\,
            in2 => \N__18635\,
            in3 => \N__19190\,
            lcout => \this_sprites_ram_mem_N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__20258\,
            in1 => \N__19184\,
            in2 => \N__19421\,
            in3 => \N__22001\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIB2RF1_3_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__20953\,
            in1 => \N__19165\,
            in2 => \_gnd_net_\,
            in3 => \N__20257\,
            lcout => \M_this_sprites_ram_write_en_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI84774_0_LC_23_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__19391\,
            in1 => \N__19619\,
            in2 => \N__19289\,
            in3 => \N__20447\,
            lcout => \M_this_ppu_vram_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI04774_0_LC_23_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__19387\,
            in1 => \N__19493\,
            in2 => \N__19285\,
            in3 => \N__19556\,
            lcout => \M_this_ppu_vram_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIH7O01_0_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__20531\,
            in1 => \N__19217\,
            in2 => \N__20674\,
            in3 => \N__19205\,
            lcout => \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIDVQ81_7_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__19183\,
            in1 => \N__20954\,
            in2 => \_gnd_net_\,
            in3 => \N__20262\,
            lcout => \un1_M_this_state_q_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI1B0E_7_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19182\,
            in2 => \_gnd_net_\,
            in3 => \N__20373\,
            lcout => \N_170_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_7_0_wclke_3_LC_23_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21300\,
            in1 => \N__21029\,
            in2 => \N__21156\,
            in3 => \N__21234\,
            lcout => \this_sprites_ram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIH7O01_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__20547\,
            in1 => \N__19676\,
            in2 => \N__20673\,
            in3 => \N__19661\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNI9LUP1_LC_24_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__19649\,
            in1 => \N__19631\,
            in2 => \N__19622\,
            in3 => \N__20548\,
            lcout => \this_sprites_ram_mem_N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNIHBQ01_LC_24_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__20549\,
            in1 => \N__19613\,
            in2 => \N__20684\,
            in3 => \N__19598\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNI9T2Q1_LC_24_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__19586\,
            in1 => \N__19577\,
            in2 => \N__19559\,
            in3 => \N__20551\,
            lcout => \this_sprites_ram_mem_N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIF7O01_LC_24_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__19550\,
            in1 => \N__20682\,
            in2 => \N__19535\,
            in3 => \N__20550\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNI5LUP1_LC_24_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__20552\,
            in1 => \N__19517\,
            in2 => \N__19502\,
            in3 => \N__19499\,
            lcout => \this_sprites_ram_mem_N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__21326\,
            in1 => \N__21072\,
            in2 => \N__21185\,
            in3 => \N__21259\,
            lcout => \this_sprites_ram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21260\,
            in1 => \N__21182\,
            in2 => \N__21077\,
            in3 => \N__21327\,
            lcout => \this_sprites_ram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21325\,
            in1 => \N__21071\,
            in2 => \N__21184\,
            in3 => \N__21258\,
            lcout => \this_sprites_ram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNIJBQ01_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__20532\,
            in1 => \N__20696\,
            in2 => \N__20678\,
            in3 => \N__20588\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIDT2Q1_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__20576\,
            in1 => \N__20561\,
            in2 => \N__20555\,
            in3 => \N__20533\,
            lcout => \this_sprites_ram_mem_N_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21324\,
            in1 => \N__21060\,
            in2 => \N__21175\,
            in3 => \N__21249\,
            lcout => \this_sprites_ram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21331\,
            in1 => \N__21050\,
            in2 => \N__21161\,
            in3 => \N__21247\,
            lcout => \this_sprites_ram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI9MQ11_2_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20387\,
            in2 => \_gnd_net_\,
            in3 => \N__20291\,
            lcout => \M_this_sprites_ram_write_data_0_sqmuxa\,
            ltout => \M_this_sprites_ram_write_data_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_ibuf_RNIGSD53_0_LC_24_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__20173\,
            in1 => \N__20118\,
            in2 => \N__20075\,
            in3 => \N__21488\,
            lcout => \M_this_sprites_ram_write_data_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_ibuf_RNIM2E53_7_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__19978\,
            in1 => \N__21489\,
            in2 => \N__19940\,
            in3 => \N__21423\,
            lcout => \M_this_sprites_ram_write_data_0_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_ibuf_RNIK0E53_2_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__19827\,
            in1 => \N__21491\,
            in2 => \N__19788\,
            in3 => \N__21425\,
            lcout => \M_this_sprites_ram_write_data_0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_ibuf_RNIIUD53_1_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__21531\,
            in1 => \N__21490\,
            in2 => \N__21465\,
            in3 => \N__21424\,
            lcout => \M_this_sprites_ram_write_data_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__21320\,
            in1 => \N__21248\,
            in2 => \N__21160\,
            in3 => \N__21030\,
            lcout => \this_sprites_ram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_0_LC_30_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22482\,
            in1 => \N__20824\,
            in2 => \N__20974\,
            in3 => \N__20969\,
            lcout => \M_this_external_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_30_23_0_\,
            carryout => \un1_M_this_external_address_q_cry_0\,
            clk => \N__22239\,
            ce => 'H',
            sr => \N__21945\
        );

    \M_this_external_address_q_1_LC_30_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22488\,
            in1 => \N__20803\,
            in2 => \_gnd_net_\,
            in3 => \N__20792\,
            lcout => \M_this_external_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_0\,
            carryout => \un1_M_this_external_address_q_cry_1\,
            clk => \N__22239\,
            ce => 'H',
            sr => \N__21945\
        );

    \M_this_external_address_q_2_LC_30_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22483\,
            in1 => \N__20773\,
            in2 => \_gnd_net_\,
            in3 => \N__20762\,
            lcout => \M_this_external_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_1\,
            carryout => \un1_M_this_external_address_q_cry_2\,
            clk => \N__22239\,
            ce => 'H',
            sr => \N__21945\
        );

    \M_this_external_address_q_3_LC_30_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22489\,
            in1 => \N__20749\,
            in2 => \_gnd_net_\,
            in3 => \N__20738\,
            lcout => \M_this_external_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_2\,
            carryout => \un1_M_this_external_address_q_cry_3\,
            clk => \N__22239\,
            ce => 'H',
            sr => \N__21945\
        );

    \M_this_external_address_q_4_LC_30_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22484\,
            in1 => \N__20731\,
            in2 => \_gnd_net_\,
            in3 => \N__20720\,
            lcout => \M_this_external_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_3\,
            carryout => \un1_M_this_external_address_q_cry_4\,
            clk => \N__22239\,
            ce => 'H',
            sr => \N__21945\
        );

    \M_this_external_address_q_5_LC_30_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22486\,
            in1 => \N__20710\,
            in2 => \_gnd_net_\,
            in3 => \N__20699\,
            lcout => \M_this_external_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_4\,
            carryout => \un1_M_this_external_address_q_cry_5\,
            clk => \N__22239\,
            ce => 'H',
            sr => \N__21945\
        );

    \M_this_external_address_q_6_LC_30_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22485\,
            in1 => \N__21727\,
            in2 => \_gnd_net_\,
            in3 => \N__21716\,
            lcout => \M_this_external_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_5\,
            carryout => \un1_M_this_external_address_q_cry_6\,
            clk => \N__22239\,
            ce => 'H',
            sr => \N__21945\
        );

    \M_this_external_address_q_7_LC_30_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22487\,
            in1 => \N__21700\,
            in2 => \_gnd_net_\,
            in3 => \N__21689\,
            lcout => \M_this_external_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_6\,
            carryout => \un1_M_this_external_address_q_cry_7\,
            clk => \N__22239\,
            ce => 'H',
            sr => \N__21945\
        );

    \M_this_external_address_q_8_LC_30_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22507\,
            in1 => \N__21667\,
            in2 => \_gnd_net_\,
            in3 => \N__21656\,
            lcout => \M_this_external_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_30_24_0_\,
            carryout => \un1_M_this_external_address_q_cry_8\,
            clk => \N__22242\,
            ce => 'H',
            sr => \N__21944\
        );

    \M_this_external_address_q_9_LC_30_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22492\,
            in1 => \N__21646\,
            in2 => \_gnd_net_\,
            in3 => \N__21635\,
            lcout => \M_this_external_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_8\,
            carryout => \un1_M_this_external_address_q_cry_9\,
            clk => \N__22242\,
            ce => 'H',
            sr => \N__21944\
        );

    \M_this_external_address_q_10_LC_30_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22504\,
            in1 => \N__21616\,
            in2 => \_gnd_net_\,
            in3 => \N__21605\,
            lcout => \M_this_external_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_9\,
            carryout => \un1_M_this_external_address_q_cry_10\,
            clk => \N__22242\,
            ce => 'H',
            sr => \N__21944\
        );

    \M_this_external_address_q_11_LC_30_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22490\,
            in1 => \N__21598\,
            in2 => \_gnd_net_\,
            in3 => \N__21587\,
            lcout => \M_this_external_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_10\,
            carryout => \un1_M_this_external_address_q_cry_11\,
            clk => \N__22242\,
            ce => 'H',
            sr => \N__21944\
        );

    \M_this_external_address_q_12_LC_30_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22505\,
            in1 => \N__21580\,
            in2 => \_gnd_net_\,
            in3 => \N__21569\,
            lcout => \M_this_external_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_11\,
            carryout => \un1_M_this_external_address_q_cry_12\,
            clk => \N__22242\,
            ce => 'H',
            sr => \N__21944\
        );

    \M_this_external_address_q_13_LC_30_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__22491\,
            in1 => \N__21556\,
            in2 => \_gnd_net_\,
            in3 => \N__21545\,
            lcout => \M_this_external_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_12\,
            carryout => \un1_M_this_external_address_q_cry_13\,
            clk => \N__22242\,
            ce => 'H',
            sr => \N__21944\
        );

    \M_this_external_address_q_14_LC_30_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22506\,
            in1 => \N__22522\,
            in2 => \_gnd_net_\,
            in3 => \N__22511\,
            lcout => \M_this_external_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_13\,
            carryout => \un1_M_this_external_address_q_cry_14\,
            clk => \N__22242\,
            ce => 'H',
            sr => \N__21944\
        );

    \M_this_external_address_q_15_LC_30_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111101110"
        )
    port map (
            in0 => \N__22255\,
            in1 => \N__22508\,
            in2 => \_gnd_net_\,
            in3 => \N__22271\,
            lcout => \M_this_external_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22242\,
            ce => 'H',
            sr => \N__21944\
        );

    \port_address_iobuf_RNI6NG6_2_LC_32_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21857\,
            in1 => \N__21845\,
            in2 => \N__21839\,
            in3 => \N__21830\,
            lcout => OPEN,
            ltout => \M_this_state_d36_2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_address_iobuf_RNIV8P9_6_LC_32_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__21806\,
            in1 => \_gnd_net_\,
            in2 => \N__21782\,
            in3 => \N__21779\,
            lcout => \M_this_state_d37_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
