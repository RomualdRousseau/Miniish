// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 22 2022 16:14:27

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    input [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__22940;
    wire N__22939;
    wire N__22938;
    wire N__22929;
    wire N__22928;
    wire N__22927;
    wire N__22920;
    wire N__22919;
    wire N__22918;
    wire N__22911;
    wire N__22910;
    wire N__22909;
    wire N__22902;
    wire N__22901;
    wire N__22900;
    wire N__22893;
    wire N__22892;
    wire N__22891;
    wire N__22884;
    wire N__22883;
    wire N__22882;
    wire N__22875;
    wire N__22874;
    wire N__22873;
    wire N__22866;
    wire N__22865;
    wire N__22864;
    wire N__22857;
    wire N__22856;
    wire N__22855;
    wire N__22848;
    wire N__22847;
    wire N__22846;
    wire N__22839;
    wire N__22838;
    wire N__22837;
    wire N__22830;
    wire N__22829;
    wire N__22828;
    wire N__22821;
    wire N__22820;
    wire N__22819;
    wire N__22812;
    wire N__22811;
    wire N__22810;
    wire N__22803;
    wire N__22802;
    wire N__22801;
    wire N__22794;
    wire N__22793;
    wire N__22792;
    wire N__22785;
    wire N__22784;
    wire N__22783;
    wire N__22776;
    wire N__22775;
    wire N__22774;
    wire N__22767;
    wire N__22766;
    wire N__22765;
    wire N__22758;
    wire N__22757;
    wire N__22756;
    wire N__22749;
    wire N__22748;
    wire N__22747;
    wire N__22740;
    wire N__22739;
    wire N__22738;
    wire N__22731;
    wire N__22730;
    wire N__22729;
    wire N__22722;
    wire N__22721;
    wire N__22720;
    wire N__22713;
    wire N__22712;
    wire N__22711;
    wire N__22704;
    wire N__22703;
    wire N__22702;
    wire N__22695;
    wire N__22694;
    wire N__22693;
    wire N__22686;
    wire N__22685;
    wire N__22684;
    wire N__22677;
    wire N__22676;
    wire N__22675;
    wire N__22668;
    wire N__22667;
    wire N__22666;
    wire N__22659;
    wire N__22658;
    wire N__22657;
    wire N__22650;
    wire N__22649;
    wire N__22648;
    wire N__22641;
    wire N__22640;
    wire N__22639;
    wire N__22632;
    wire N__22631;
    wire N__22630;
    wire N__22623;
    wire N__22622;
    wire N__22621;
    wire N__22614;
    wire N__22613;
    wire N__22612;
    wire N__22605;
    wire N__22604;
    wire N__22603;
    wire N__22596;
    wire N__22595;
    wire N__22594;
    wire N__22587;
    wire N__22586;
    wire N__22585;
    wire N__22578;
    wire N__22577;
    wire N__22576;
    wire N__22569;
    wire N__22568;
    wire N__22567;
    wire N__22560;
    wire N__22559;
    wire N__22558;
    wire N__22551;
    wire N__22550;
    wire N__22549;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22511;
    wire N__22508;
    wire N__22507;
    wire N__22506;
    wire N__22505;
    wire N__22504;
    wire N__22493;
    wire N__22492;
    wire N__22491;
    wire N__22490;
    wire N__22489;
    wire N__22488;
    wire N__22487;
    wire N__22486;
    wire N__22485;
    wire N__22484;
    wire N__22483;
    wire N__22482;
    wire N__22479;
    wire N__22472;
    wire N__22463;
    wire N__22454;
    wire N__22453;
    wire N__22452;
    wire N__22451;
    wire N__22450;
    wire N__22449;
    wire N__22448;
    wire N__22447;
    wire N__22444;
    wire N__22439;
    wire N__22436;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22428;
    wire N__22427;
    wire N__22424;
    wire N__22423;
    wire N__22422;
    wire N__22421;
    wire N__22420;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22400;
    wire N__22397;
    wire N__22396;
    wire N__22395;
    wire N__22392;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22365;
    wire N__22362;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22343;
    wire N__22338;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22316;
    wire N__22309;
    wire N__22306;
    wire N__22301;
    wire N__22296;
    wire N__22291;
    wire N__22278;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22244;
    wire N__22243;
    wire N__22242;
    wire N__22241;
    wire N__22240;
    wire N__22239;
    wire N__22238;
    wire N__22237;
    wire N__22236;
    wire N__22235;
    wire N__22234;
    wire N__22233;
    wire N__22232;
    wire N__22231;
    wire N__22230;
    wire N__22229;
    wire N__22228;
    wire N__22227;
    wire N__22226;
    wire N__22225;
    wire N__22224;
    wire N__22223;
    wire N__22222;
    wire N__22221;
    wire N__22220;
    wire N__22219;
    wire N__22218;
    wire N__22217;
    wire N__22216;
    wire N__22215;
    wire N__22214;
    wire N__22213;
    wire N__22212;
    wire N__22211;
    wire N__22210;
    wire N__22209;
    wire N__22208;
    wire N__22207;
    wire N__22206;
    wire N__22205;
    wire N__22204;
    wire N__22203;
    wire N__22202;
    wire N__22201;
    wire N__22200;
    wire N__22199;
    wire N__22198;
    wire N__22197;
    wire N__22196;
    wire N__22195;
    wire N__22194;
    wire N__22193;
    wire N__22192;
    wire N__22191;
    wire N__22190;
    wire N__22189;
    wire N__22188;
    wire N__22187;
    wire N__22186;
    wire N__22185;
    wire N__22184;
    wire N__22183;
    wire N__22182;
    wire N__22181;
    wire N__22180;
    wire N__22179;
    wire N__22178;
    wire N__22177;
    wire N__22176;
    wire N__22175;
    wire N__22174;
    wire N__22173;
    wire N__22172;
    wire N__22171;
    wire N__22170;
    wire N__22169;
    wire N__22168;
    wire N__22167;
    wire N__22166;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__22000;
    wire N__21999;
    wire N__21998;
    wire N__21997;
    wire N__21996;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21988;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21946;
    wire N__21945;
    wire N__21944;
    wire N__21943;
    wire N__21942;
    wire N__21941;
    wire N__21940;
    wire N__21939;
    wire N__21938;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21766;
    wire N__21765;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21745;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21491;
    wire N__21490;
    wire N__21489;
    wire N__21488;
    wire N__21483;
    wire N__21478;
    wire N__21473;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21425;
    wire N__21424;
    wire N__21423;
    wire N__21418;
    wire N__21415;
    wire N__21410;
    wire N__21407;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21399;
    wire N__21394;
    wire N__21391;
    wire N__21390;
    wire N__21389;
    wire N__21384;
    wire N__21381;
    wire N__21380;
    wire N__21377;
    wire N__21376;
    wire N__21371;
    wire N__21368;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21356;
    wire N__21353;
    wire N__21348;
    wire N__21343;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21328;
    wire N__21327;
    wire N__21326;
    wire N__21325;
    wire N__21324;
    wire N__21321;
    wire N__21320;
    wire N__21317;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21301;
    wire N__21300;
    wire N__21297;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21282;
    wire N__21281;
    wire N__21270;
    wire N__21265;
    wire N__21260;
    wire N__21259;
    wire N__21258;
    wire N__21257;
    wire N__21250;
    wire N__21249;
    wire N__21248;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21185;
    wire N__21184;
    wire N__21183;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21175;
    wire N__21172;
    wire N__21165;
    wire N__21162;
    wire N__21161;
    wire N__21160;
    wire N__21157;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21106;
    wire N__21101;
    wire N__21096;
    wire N__21093;
    wire N__21092;
    wire N__21085;
    wire N__21082;
    wire N__21077;
    wire N__21076;
    wire N__21073;
    wire N__21072;
    wire N__21071;
    wire N__21068;
    wire N__21061;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21050;
    wire N__21047;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21031;
    wire N__21030;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21016;
    wire N__21015;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20993;
    wire N__20990;
    wire N__20989;
    wire N__20986;
    wire N__20983;
    wire N__20978;
    wire N__20975;
    wire N__20974;
    wire N__20973;
    wire N__20970;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20962;
    wire N__20961;
    wire N__20960;
    wire N__20959;
    wire N__20958;
    wire N__20955;
    wire N__20954;
    wire N__20953;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20938;
    wire N__20931;
    wire N__20930;
    wire N__20929;
    wire N__20928;
    wire N__20927;
    wire N__20926;
    wire N__20925;
    wire N__20924;
    wire N__20923;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20897;
    wire N__20888;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20868;
    wire N__20861;
    wire N__20854;
    wire N__20851;
    wire N__20846;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20683;
    wire N__20682;
    wire N__20679;
    wire N__20678;
    wire N__20675;
    wire N__20674;
    wire N__20673;
    wire N__20672;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20625;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20597;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20551;
    wire N__20550;
    wire N__20549;
    wire N__20548;
    wire N__20547;
    wire N__20546;
    wire N__20537;
    wire N__20536;
    wire N__20535;
    wire N__20534;
    wire N__20533;
    wire N__20532;
    wire N__20531;
    wire N__20530;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20514;
    wire N__20511;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20496;
    wire N__20495;
    wire N__20488;
    wire N__20481;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20459;
    wire N__20456;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20414;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20390;
    wire N__20389;
    wire N__20388;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20377;
    wire N__20374;
    wire N__20373;
    wire N__20370;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20343;
    wire N__20336;
    wire N__20335;
    wire N__20332;
    wire N__20331;
    wire N__20328;
    wire N__20327;
    wire N__20326;
    wire N__20325;
    wire N__20324;
    wire N__20323;
    wire N__20322;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20291;
    wire N__20290;
    wire N__20289;
    wire N__20288;
    wire N__20287;
    wire N__20286;
    wire N__20283;
    wire N__20282;
    wire N__20281;
    wire N__20270;
    wire N__20263;
    wire N__20262;
    wire N__20259;
    wire N__20258;
    wire N__20257;
    wire N__20256;
    wire N__20255;
    wire N__20254;
    wire N__20251;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20216;
    wire N__20213;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20185;
    wire N__20174;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20120;
    wire N__20119;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20051;
    wire N__20050;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20038;
    wire N__20035;
    wire N__20034;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20012;
    wire N__20009;
    wire N__20004;
    wire N__20003;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19911;
    wire N__19906;
    wire N__19903;
    wire N__19902;
    wire N__19901;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19889;
    wire N__19888;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19866;
    wire N__19863;
    wire N__19862;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19844;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19810;
    wire N__19807;
    wire N__19804;
    wire N__19799;
    wire N__19796;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19756;
    wire N__19753;
    wire N__19748;
    wire N__19745;
    wire N__19744;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19736;
    wire N__19733;
    wire N__19732;
    wire N__19727;
    wire N__19724;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19712;
    wire N__19709;
    wire N__19708;
    wire N__19703;
    wire N__19698;
    wire N__19695;
    wire N__19694;
    wire N__19691;
    wire N__19686;
    wire N__19683;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19463;
    wire N__19460;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19387;
    wire N__19386;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19378;
    wire N__19375;
    wire N__19374;
    wire N__19373;
    wire N__19372;
    wire N__19369;
    wire N__19368;
    wire N__19367;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19322;
    wire N__19319;
    wire N__19314;
    wire N__19311;
    wire N__19306;
    wire N__19303;
    wire N__19298;
    wire N__19289;
    wire N__19286;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19183;
    wire N__19182;
    wire N__19179;
    wire N__19174;
    wire N__19169;
    wire N__19166;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19151;
    wire N__19148;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19126;
    wire N__19125;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19105;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18965;
    wire N__18962;
    wire N__18961;
    wire N__18960;
    wire N__18955;
    wire N__18952;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18903;
    wire N__18902;
    wire N__18901;
    wire N__18900;
    wire N__18897;
    wire N__18896;
    wire N__18895;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18880;
    wire N__18877;
    wire N__18872;
    wire N__18869;
    wire N__18862;
    wire N__18859;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18595;
    wire N__18592;
    wire N__18591;
    wire N__18590;
    wire N__18587;
    wire N__18586;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18568;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18433;
    wire N__18432;
    wire N__18431;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18405;
    wire N__18402;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18274;
    wire N__18271;
    wire N__18270;
    wire N__18269;
    wire N__18266;
    wire N__18265;
    wire N__18262;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18115;
    wire N__18114;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18090;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17959;
    wire N__17956;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17944;
    wire N__17943;
    wire N__17940;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17797;
    wire N__17796;
    wire N__17793;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17646;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17512;
    wire N__17511;
    wire N__17510;
    wire N__17509;
    wire N__17508;
    wire N__17507;
    wire N__17506;
    wire N__17505;
    wire N__17504;
    wire N__17499;
    wire N__17496;
    wire N__17495;
    wire N__17494;
    wire N__17491;
    wire N__17484;
    wire N__17483;
    wire N__17482;
    wire N__17479;
    wire N__17474;
    wire N__17469;
    wire N__17464;
    wire N__17459;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17439;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17336;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17323;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17304;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17290;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17100;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17086;
    wire N__17085;
    wire N__17082;
    wire N__17081;
    wire N__17076;
    wire N__17073;
    wire N__17070;
    wire N__17067;
    wire N__17064;
    wire N__17061;
    wire N__17056;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17035;
    wire N__17032;
    wire N__17031;
    wire N__17028;
    wire N__17027;
    wire N__17026;
    wire N__17025;
    wire N__17022;
    wire N__17021;
    wire N__17018;
    wire N__17013;
    wire N__17010;
    wire N__17007;
    wire N__17004;
    wire N__17001;
    wire N__16998;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16867;
    wire N__16866;
    wire N__16865;
    wire N__16864;
    wire N__16863;
    wire N__16856;
    wire N__16851;
    wire N__16850;
    wire N__16847;
    wire N__16842;
    wire N__16839;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16716;
    wire N__16713;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16701;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16437;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16425;
    wire N__16418;
    wire N__16417;
    wire N__16416;
    wire N__16415;
    wire N__16414;
    wire N__16413;
    wire N__16412;
    wire N__16411;
    wire N__16410;
    wire N__16405;
    wire N__16404;
    wire N__16401;
    wire N__16400;
    wire N__16397;
    wire N__16396;
    wire N__16393;
    wire N__16390;
    wire N__16387;
    wire N__16386;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16375;
    wire N__16372;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16324;
    wire N__16313;
    wire N__16310;
    wire N__16305;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16285;
    wire N__16280;
    wire N__16277;
    wire N__16276;
    wire N__16275;
    wire N__16272;
    wire N__16269;
    wire N__16266;
    wire N__16263;
    wire N__16256;
    wire N__16253;
    wire N__16250;
    wire N__16249;
    wire N__16248;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16236;
    wire N__16233;
    wire N__16230;
    wire N__16227;
    wire N__16220;
    wire N__16217;
    wire N__16216;
    wire N__16215;
    wire N__16214;
    wire N__16213;
    wire N__16210;
    wire N__16205;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16193;
    wire N__16190;
    wire N__16185;
    wire N__16182;
    wire N__16175;
    wire N__16174;
    wire N__16171;
    wire N__16170;
    wire N__16167;
    wire N__16162;
    wire N__16161;
    wire N__16160;
    wire N__16159;
    wire N__16158;
    wire N__16153;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16133;
    wire N__16132;
    wire N__16131;
    wire N__16124;
    wire N__16121;
    wire N__16120;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16103;
    wire N__16102;
    wire N__16101;
    wire N__16098;
    wire N__16093;
    wire N__16088;
    wire N__16085;
    wire N__16082;
    wire N__16081;
    wire N__16076;
    wire N__16073;
    wire N__16072;
    wire N__16071;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16055;
    wire N__16054;
    wire N__16053;
    wire N__16046;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16019;
    wire N__16018;
    wire N__16017;
    wire N__16016;
    wire N__16013;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15985;
    wire N__15982;
    wire N__15977;
    wire N__15976;
    wire N__15975;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15925;
    wire N__15922;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15908;
    wire N__15907;
    wire N__15906;
    wire N__15905;
    wire N__15904;
    wire N__15903;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15889;
    wire N__15888;
    wire N__15887;
    wire N__15884;
    wire N__15883;
    wire N__15882;
    wire N__15881;
    wire N__15880;
    wire N__15877;
    wire N__15876;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15861;
    wire N__15858;
    wire N__15855;
    wire N__15854;
    wire N__15853;
    wire N__15850;
    wire N__15849;
    wire N__15848;
    wire N__15845;
    wire N__15842;
    wire N__15841;
    wire N__15840;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15830;
    wire N__15829;
    wire N__15826;
    wire N__15823;
    wire N__15820;
    wire N__15817;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15799;
    wire N__15798;
    wire N__15797;
    wire N__15794;
    wire N__15791;
    wire N__15790;
    wire N__15787;
    wire N__15786;
    wire N__15781;
    wire N__15778;
    wire N__15775;
    wire N__15774;
    wire N__15769;
    wire N__15766;
    wire N__15763;
    wire N__15760;
    wire N__15759;
    wire N__15758;
    wire N__15753;
    wire N__15750;
    wire N__15741;
    wire N__15738;
    wire N__15735;
    wire N__15734;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15688;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15670;
    wire N__15669;
    wire N__15668;
    wire N__15665;
    wire N__15660;
    wire N__15657;
    wire N__15652;
    wire N__15645;
    wire N__15638;
    wire N__15635;
    wire N__15628;
    wire N__15625;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15611;
    wire N__15606;
    wire N__15599;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15570;
    wire N__15567;
    wire N__15560;
    wire N__15557;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15542;
    wire N__15539;
    wire N__15536;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15493;
    wire N__15490;
    wire N__15487;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15464;
    wire N__15461;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15443;
    wire N__15440;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15422;
    wire N__15419;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15398;
    wire N__15395;
    wire N__15394;
    wire N__15391;
    wire N__15388;
    wire N__15385;
    wire N__15382;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15283;
    wire N__15280;
    wire N__15277;
    wire N__15274;
    wire N__15271;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15209;
    wire N__15206;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15187;
    wire N__15184;
    wire N__15181;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15139;
    wire N__15138;
    wire N__15137;
    wire N__15134;
    wire N__15129;
    wire N__15126;
    wire N__15121;
    wire N__15116;
    wire N__15115;
    wire N__15114;
    wire N__15111;
    wire N__15108;
    wire N__15105;
    wire N__15102;
    wire N__15101;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15087;
    wire N__15084;
    wire N__15077;
    wire N__15074;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15056;
    wire N__15055;
    wire N__15052;
    wire N__15049;
    wire N__15048;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15037;
    wire N__15034;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15019;
    wire N__15016;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14965;
    wire N__14964;
    wire N__14961;
    wire N__14956;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14830;
    wire N__14829;
    wire N__14826;
    wire N__14823;
    wire N__14820;
    wire N__14817;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14704;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14691;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14562;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14534;
    wire N__14533;
    wire N__14528;
    wire N__14525;
    wire N__14524;
    wire N__14523;
    wire N__14522;
    wire N__14521;
    wire N__14520;
    wire N__14519;
    wire N__14516;
    wire N__14505;
    wire N__14502;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14489;
    wire N__14484;
    wire N__14481;
    wire N__14474;
    wire N__14473;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14446;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14431;
    wire N__14428;
    wire N__14425;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14407;
    wire N__14406;
    wire N__14403;
    wire N__14400;
    wire N__14395;
    wire N__14390;
    wire N__14387;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14372;
    wire N__14369;
    wire N__14366;
    wire N__14365;
    wire N__14364;
    wire N__14361;
    wire N__14358;
    wire N__14355;
    wire N__14352;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14335;
    wire N__14334;
    wire N__14331;
    wire N__14326;
    wire N__14323;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14306;
    wire N__14305;
    wire N__14304;
    wire N__14303;
    wire N__14294;
    wire N__14291;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14269;
    wire N__14268;
    wire N__14267;
    wire N__14266;
    wire N__14265;
    wire N__14264;
    wire N__14263;
    wire N__14262;
    wire N__14261;
    wire N__14260;
    wire N__14259;
    wire N__14258;
    wire N__14257;
    wire N__14256;
    wire N__14247;
    wire N__14240;
    wire N__14239;
    wire N__14236;
    wire N__14235;
    wire N__14232;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14220;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14205;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14187;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14173;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14154;
    wire N__14149;
    wire N__14144;
    wire N__14139;
    wire N__14132;
    wire N__14123;
    wire N__14120;
    wire N__14119;
    wire N__14118;
    wire N__14117;
    wire N__14116;
    wire N__14115;
    wire N__14114;
    wire N__14111;
    wire N__14110;
    wire N__14109;
    wire N__14102;
    wire N__14101;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14071;
    wire N__14068;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14051;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13925;
    wire N__13924;
    wire N__13923;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13911;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13802;
    wire N__13799;
    wire N__13796;
    wire N__13793;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13781;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13771;
    wire N__13770;
    wire N__13767;
    wire N__13764;
    wire N__13761;
    wire N__13758;
    wire N__13751;
    wire N__13748;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13727;
    wire N__13724;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13676;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13636;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13504;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13494;
    wire N__13491;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13426;
    wire N__13425;
    wire N__13424;
    wire N__13423;
    wire N__13420;
    wire N__13419;
    wire N__13418;
    wire N__13417;
    wire N__13414;
    wire N__13411;
    wire N__13408;
    wire N__13405;
    wire N__13404;
    wire N__13403;
    wire N__13402;
    wire N__13401;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13389;
    wire N__13386;
    wire N__13381;
    wire N__13378;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13364;
    wire N__13363;
    wire N__13358;
    wire N__13353;
    wire N__13346;
    wire N__13343;
    wire N__13340;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13328;
    wire N__13325;
    wire N__13320;
    wire N__13315;
    wire N__13304;
    wire N__13303;
    wire N__13302;
    wire N__13301;
    wire N__13300;
    wire N__13297;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13285;
    wire N__13282;
    wire N__13279;
    wire N__13276;
    wire N__13273;
    wire N__13272;
    wire N__13269;
    wire N__13264;
    wire N__13259;
    wire N__13256;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13213;
    wire N__13210;
    wire N__13209;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13174;
    wire N__13173;
    wire N__13170;
    wire N__13167;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13142;
    wire N__13141;
    wire N__13138;
    wire N__13135;
    wire N__13130;
    wire N__13129;
    wire N__13126;
    wire N__13125;
    wire N__13124;
    wire N__13121;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13110;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13102;
    wire N__13101;
    wire N__13100;
    wire N__13099;
    wire N__13092;
    wire N__13089;
    wire N__13086;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13069;
    wire N__13068;
    wire N__13061;
    wire N__13056;
    wire N__13053;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13042;
    wire N__13041;
    wire N__13036;
    wire N__13035;
    wire N__13032;
    wire N__13029;
    wire N__13022;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13010;
    wire N__13007;
    wire N__13004;
    wire N__12997;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12972;
    wire N__12965;
    wire N__12964;
    wire N__12963;
    wire N__12962;
    wire N__12959;
    wire N__12958;
    wire N__12957;
    wire N__12954;
    wire N__12953;
    wire N__12952;
    wire N__12951;
    wire N__12950;
    wire N__12949;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12939;
    wire N__12936;
    wire N__12931;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12901;
    wire N__12898;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12862;
    wire N__12859;
    wire N__12856;
    wire N__12853;
    wire N__12852;
    wire N__12847;
    wire N__12844;
    wire N__12839;
    wire N__12838;
    wire N__12837;
    wire N__12836;
    wire N__12833;
    wire N__12832;
    wire N__12829;
    wire N__12828;
    wire N__12827;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12816;
    wire N__12813;
    wire N__12812;
    wire N__12811;
    wire N__12810;
    wire N__12809;
    wire N__12808;
    wire N__12807;
    wire N__12806;
    wire N__12803;
    wire N__12794;
    wire N__12793;
    wire N__12790;
    wire N__12787;
    wire N__12784;
    wire N__12781;
    wire N__12778;
    wire N__12777;
    wire N__12776;
    wire N__12775;
    wire N__12774;
    wire N__12773;
    wire N__12770;
    wire N__12769;
    wire N__12766;
    wire N__12763;
    wire N__12760;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12729;
    wire N__12728;
    wire N__12725;
    wire N__12720;
    wire N__12711;
    wire N__12710;
    wire N__12701;
    wire N__12692;
    wire N__12689;
    wire N__12682;
    wire N__12681;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12666;
    wire N__12661;
    wire N__12650;
    wire N__12649;
    wire N__12648;
    wire N__12647;
    wire N__12646;
    wire N__12645;
    wire N__12644;
    wire N__12643;
    wire N__12642;
    wire N__12641;
    wire N__12640;
    wire N__12639;
    wire N__12636;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12625;
    wire N__12624;
    wire N__12623;
    wire N__12620;
    wire N__12619;
    wire N__12618;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12610;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12602;
    wire N__12601;
    wire N__12600;
    wire N__12597;
    wire N__12596;
    wire N__12595;
    wire N__12592;
    wire N__12591;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12559;
    wire N__12554;
    wire N__12551;
    wire N__12546;
    wire N__12545;
    wire N__12542;
    wire N__12535;
    wire N__12532;
    wire N__12531;
    wire N__12528;
    wire N__12525;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12505;
    wire N__12504;
    wire N__12503;
    wire N__12498;
    wire N__12483;
    wire N__12480;
    wire N__12477;
    wire N__12472;
    wire N__12469;
    wire N__12460;
    wire N__12455;
    wire N__12450;
    wire N__12445;
    wire N__12438;
    wire N__12425;
    wire N__12422;
    wire N__12421;
    wire N__12420;
    wire N__12419;
    wire N__12418;
    wire N__12415;
    wire N__12414;
    wire N__12413;
    wire N__12410;
    wire N__12409;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12401;
    wire N__12400;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12387;
    wire N__12386;
    wire N__12385;
    wire N__12380;
    wire N__12379;
    wire N__12376;
    wire N__12373;
    wire N__12370;
    wire N__12363;
    wire N__12362;
    wire N__12361;
    wire N__12358;
    wire N__12351;
    wire N__12346;
    wire N__12343;
    wire N__12342;
    wire N__12341;
    wire N__12340;
    wire N__12339;
    wire N__12338;
    wire N__12335;
    wire N__12334;
    wire N__12331;
    wire N__12326;
    wire N__12323;
    wire N__12318;
    wire N__12309;
    wire N__12298;
    wire N__12293;
    wire N__12278;
    wire N__12277;
    wire N__12274;
    wire N__12271;
    wire N__12268;
    wire N__12265;
    wire N__12262;
    wire N__12257;
    wire N__12256;
    wire N__12255;
    wire N__12254;
    wire N__12253;
    wire N__12250;
    wire N__12249;
    wire N__12248;
    wire N__12247;
    wire N__12246;
    wire N__12243;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12220;
    wire N__12219;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12211;
    wire N__12210;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12192;
    wire N__12187;
    wire N__12186;
    wire N__12185;
    wire N__12184;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12169;
    wire N__12164;
    wire N__12157;
    wire N__12154;
    wire N__12149;
    wire N__12144;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12118;
    wire N__12117;
    wire N__12116;
    wire N__12113;
    wire N__12112;
    wire N__12111;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12090;
    wire N__12087;
    wire N__12084;
    wire N__12081;
    wire N__12068;
    wire N__12067;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12049;
    wire N__12048;
    wire N__12047;
    wire N__12046;
    wire N__12043;
    wire N__12040;
    wire N__12039;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12029;
    wire N__12024;
    wire N__12023;
    wire N__12020;
    wire N__12019;
    wire N__12016;
    wire N__12013;
    wire N__12010;
    wire N__12005;
    wire N__12002;
    wire N__11999;
    wire N__11994;
    wire N__11991;
    wire N__11978;
    wire N__11977;
    wire N__11974;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11964;
    wire N__11963;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11946;
    wire N__11939;
    wire N__11938;
    wire N__11937;
    wire N__11936;
    wire N__11935;
    wire N__11932;
    wire N__11931;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11919;
    wire N__11914;
    wire N__11911;
    wire N__11906;
    wire N__11901;
    wire N__11900;
    wire N__11897;
    wire N__11894;
    wire N__11891;
    wire N__11888;
    wire N__11881;
    wire N__11876;
    wire N__11873;
    wire N__11870;
    wire N__11867;
    wire N__11864;
    wire N__11861;
    wire N__11858;
    wire N__11855;
    wire N__11854;
    wire N__11853;
    wire N__11846;
    wire N__11843;
    wire N__11842;
    wire N__11841;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11815;
    wire N__11810;
    wire N__11807;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11797;
    wire N__11794;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11776;
    wire N__11773;
    wire N__11770;
    wire N__11769;
    wire N__11764;
    wire N__11761;
    wire N__11756;
    wire N__11753;
    wire N__11752;
    wire N__11749;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11729;
    wire N__11728;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11693;
    wire N__11690;
    wire N__11689;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11681;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11657;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11630;
    wire N__11627;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11615;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11597;
    wire N__11596;
    wire N__11595;
    wire N__11594;
    wire N__11593;
    wire N__11592;
    wire N__11591;
    wire N__11590;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11563;
    wire N__11562;
    wire N__11561;
    wire N__11560;
    wire N__11559;
    wire N__11558;
    wire N__11557;
    wire N__11556;
    wire N__11555;
    wire N__11552;
    wire N__11531;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11521;
    wire N__11520;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11512;
    wire N__11509;
    wire N__11508;
    wire N__11505;
    wire N__11500;
    wire N__11497;
    wire N__11492;
    wire N__11491;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11487;
    wire N__11486;
    wire N__11481;
    wire N__11476;
    wire N__11469;
    wire N__11462;
    wire N__11453;
    wire N__11452;
    wire N__11451;
    wire N__11450;
    wire N__11449;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11433;
    wire N__11426;
    wire N__11425;
    wire N__11424;
    wire N__11423;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11409;
    wire N__11406;
    wire N__11401;
    wire N__11398;
    wire N__11393;
    wire N__11392;
    wire N__11391;
    wire N__11390;
    wire N__11389;
    wire N__11388;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11380;
    wire N__11379;
    wire N__11372;
    wire N__11367;
    wire N__11364;
    wire N__11361;
    wire N__11360;
    wire N__11359;
    wire N__11358;
    wire N__11357;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11343;
    wire N__11342;
    wire N__11341;
    wire N__11340;
    wire N__11339;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11323;
    wire N__11320;
    wire N__11315;
    wire N__11310;
    wire N__11303;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11266;
    wire N__11261;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11237;
    wire N__11234;
    wire N__11233;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11191;
    wire N__11188;
    wire N__11187;
    wire N__11186;
    wire N__11183;
    wire N__11182;
    wire N__11179;
    wire N__11176;
    wire N__11175;
    wire N__11174;
    wire N__11173;
    wire N__11170;
    wire N__11169;
    wire N__11166;
    wire N__11163;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11145;
    wire N__11132;
    wire N__11131;
    wire N__11130;
    wire N__11129;
    wire N__11128;
    wire N__11127;
    wire N__11124;
    wire N__11123;
    wire N__11122;
    wire N__11121;
    wire N__11120;
    wire N__11115;
    wire N__11112;
    wire N__11111;
    wire N__11108;
    wire N__11107;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11084;
    wire N__11075;
    wire N__11060;
    wire N__11059;
    wire N__11058;
    wire N__11057;
    wire N__11056;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11048;
    wire N__11047;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11015;
    wire N__11006;
    wire N__10999;
    wire N__10988;
    wire N__10987;
    wire N__10984;
    wire N__10983;
    wire N__10982;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10974;
    wire N__10973;
    wire N__10972;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10957;
    wire N__10954;
    wire N__10951;
    wire N__10944;
    wire N__10931;
    wire N__10928;
    wire N__10927;
    wire N__10924;
    wire N__10923;
    wire N__10920;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10909;
    wire N__10908;
    wire N__10907;
    wire N__10906;
    wire N__10905;
    wire N__10902;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10882;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10837;
    wire N__10834;
    wire N__10831;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10810;
    wire N__10809;
    wire N__10808;
    wire N__10807;
    wire N__10806;
    wire N__10805;
    wire N__10802;
    wire N__10801;
    wire N__10796;
    wire N__10793;
    wire N__10792;
    wire N__10791;
    wire N__10790;
    wire N__10789;
    wire N__10784;
    wire N__10783;
    wire N__10780;
    wire N__10779;
    wire N__10774;
    wire N__10773;
    wire N__10768;
    wire N__10767;
    wire N__10766;
    wire N__10765;
    wire N__10764;
    wire N__10761;
    wire N__10760;
    wire N__10757;
    wire N__10756;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10715;
    wire N__10704;
    wire N__10685;
    wire N__10682;
    wire N__10681;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10673;
    wire N__10672;
    wire N__10671;
    wire N__10670;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10648;
    wire N__10647;
    wire N__10646;
    wire N__10645;
    wire N__10644;
    wire N__10643;
    wire N__10642;
    wire N__10641;
    wire N__10640;
    wire N__10639;
    wire N__10638;
    wire N__10635;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10607;
    wire N__10594;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10568;
    wire N__10565;
    wire N__10562;
    wire N__10561;
    wire N__10558;
    wire N__10555;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10528;
    wire N__10525;
    wire N__10524;
    wire N__10523;
    wire N__10522;
    wire N__10519;
    wire N__10516;
    wire N__10513;
    wire N__10508;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10474;
    wire N__10471;
    wire N__10468;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10453;
    wire N__10452;
    wire N__10451;
    wire N__10450;
    wire N__10449;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10435;
    wire N__10430;
    wire N__10427;
    wire N__10418;
    wire N__10415;
    wire N__10414;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10393;
    wire N__10392;
    wire N__10391;
    wire N__10390;
    wire N__10389;
    wire N__10388;
    wire N__10387;
    wire N__10386;
    wire N__10383;
    wire N__10380;
    wire N__10375;
    wire N__10372;
    wire N__10367;
    wire N__10362;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10342;
    wire N__10339;
    wire N__10336;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10321;
    wire N__10320;
    wire N__10319;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10273;
    wire N__10272;
    wire N__10271;
    wire N__10270;
    wire N__10269;
    wire N__10264;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10248;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10234;
    wire N__10233;
    wire N__10232;
    wire N__10231;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10221;
    wire N__10214;
    wire N__10209;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10141;
    wire N__10140;
    wire N__10135;
    wire N__10134;
    wire N__10133;
    wire N__10130;
    wire N__10129;
    wire N__10128;
    wire N__10127;
    wire N__10124;
    wire N__10123;
    wire N__10122;
    wire N__10117;
    wire N__10114;
    wire N__10113;
    wire N__10110;
    wire N__10109;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10090;
    wire N__10083;
    wire N__10076;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10048;
    wire N__10047;
    wire N__10044;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10029;
    wire N__10026;
    wire N__10023;
    wire N__10020;
    wire N__10013;
    wire N__10012;
    wire N__10011;
    wire N__10010;
    wire N__10009;
    wire N__10008;
    wire N__10007;
    wire N__10006;
    wire N__10005;
    wire N__10002;
    wire N__10001;
    wire N__10000;
    wire N__9999;
    wire N__9998;
    wire N__9997;
    wire N__9994;
    wire N__9991;
    wire N__9988;
    wire N__9983;
    wire N__9978;
    wire N__9973;
    wire N__9962;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9937;
    wire N__9936;
    wire N__9933;
    wire N__9928;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9916;
    wire N__9915;
    wire N__9914;
    wire N__9913;
    wire N__9912;
    wire N__9911;
    wire N__9910;
    wire N__9909;
    wire N__9908;
    wire N__9907;
    wire N__9906;
    wire N__9903;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9895;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9887;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9869;
    wire N__9864;
    wire N__9855;
    wire N__9846;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9826;
    wire N__9823;
    wire N__9822;
    wire N__9821;
    wire N__9820;
    wire N__9819;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9805;
    wire N__9800;
    wire N__9797;
    wire N__9796;
    wire N__9791;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9763;
    wire N__9762;
    wire N__9761;
    wire N__9756;
    wire N__9753;
    wire N__9752;
    wire N__9751;
    wire N__9750;
    wire N__9747;
    wire N__9746;
    wire N__9745;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9735;
    wire N__9732;
    wire N__9727;
    wire N__9722;
    wire N__9721;
    wire N__9716;
    wire N__9709;
    wire N__9704;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9692;
    wire N__9689;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9601;
    wire N__9600;
    wire N__9597;
    wire N__9596;
    wire N__9593;
    wire N__9592;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9578;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9559;
    wire N__9558;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9544;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9505;
    wire N__9504;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9492;
    wire N__9485;
    wire N__9482;
    wire N__9481;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9403;
    wire N__9402;
    wire N__9401;
    wire N__9400;
    wire N__9399;
    wire N__9396;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9381;
    wire N__9376;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9355;
    wire N__9354;
    wire N__9353;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9319;
    wire N__9314;
    wire N__9311;
    wire N__9310;
    wire N__9309;
    wire N__9304;
    wire N__9301;
    wire N__9296;
    wire N__9293;
    wire N__9292;
    wire N__9291;
    wire N__9286;
    wire N__9283;
    wire N__9278;
    wire N__9275;
    wire N__9274;
    wire N__9273;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9261;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9247;
    wire N__9244;
    wire N__9239;
    wire N__9236;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9224;
    wire N__9221;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9207;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9185;
    wire N__9184;
    wire N__9183;
    wire N__9180;
    wire N__9175;
    wire N__9170;
    wire N__9167;
    wire N__9166;
    wire N__9165;
    wire N__9164;
    wire N__9161;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9138;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9093;
    wire N__9092;
    wire N__9091;
    wire N__9088;
    wire N__9087;
    wire N__9086;
    wire N__9083;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9031;
    wire N__9030;
    wire N__9029;
    wire N__9028;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9012;
    wire N__9009;
    wire N__9008;
    wire N__9007;
    wire N__9006;
    wire N__9005;
    wire N__9002;
    wire N__8997;
    wire N__8990;
    wire N__8981;
    wire N__8976;
    wire N__8967;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8924;
    wire N__8921;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8875;
    wire N__8874;
    wire N__8873;
    wire N__8872;
    wire N__8869;
    wire N__8864;
    wire N__8859;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8782;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8753;
    wire N__8752;
    wire N__8747;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8732;
    wire N__8731;
    wire N__8730;
    wire N__8725;
    wire N__8722;
    wire N__8717;
    wire N__8714;
    wire N__8713;
    wire N__8712;
    wire N__8709;
    wire N__8704;
    wire N__8699;
    wire N__8698;
    wire N__8697;
    wire N__8694;
    wire N__8693;
    wire N__8688;
    wire N__8683;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8644;
    wire N__8643;
    wire N__8640;
    wire N__8635;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8560;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8479;
    wire N__8476;
    wire N__8473;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8320;
    wire N__8319;
    wire N__8318;
    wire N__8317;
    wire N__8316;
    wire N__8311;
    wire N__8308;
    wire N__8301;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8279;
    wire N__8278;
    wire N__8273;
    wire N__8270;
    wire N__8269;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8258;
    wire N__8253;
    wire N__8248;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8179;
    wire N__8178;
    wire N__8177;
    wire N__8174;
    wire N__8169;
    wire N__8166;
    wire N__8159;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8113;
    wire N__8112;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8104;
    wire N__8103;
    wire N__8092;
    wire N__8089;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8008;
    wire N__8007;
    wire N__8004;
    wire N__7999;
    wire N__7998;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7987;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7969;
    wire N__7966;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7945;
    wire N__7942;
    wire N__7939;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7921;
    wire N__7918;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7867;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7853;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7798;
    wire N__7797;
    wire N__7796;
    wire N__7787;
    wire N__7786;
    wire N__7785;
    wire N__7782;
    wire N__7777;
    wire N__7774;
    wire N__7771;
    wire N__7766;
    wire N__7763;
    wire N__7762;
    wire N__7761;
    wire N__7760;
    wire N__7759;
    wire N__7758;
    wire N__7753;
    wire N__7744;
    wire N__7739;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7729;
    wire N__7728;
    wire N__7727;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7706;
    wire N__7703;
    wire N__7698;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7681;
    wire N__7680;
    wire N__7679;
    wire N__7678;
    wire N__7677;
    wire N__7672;
    wire N__7667;
    wire N__7662;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire VCCG0;
    wire \this_vga_signals.N_340_0 ;
    wire N_198_i;
    wire rgb_c_0;
    wire rgb_c_4;
    wire port_nmib_0_i;
    wire rgb_c_3;
    wire rgb_c_5;
    wire this_vga_signals_vvisibility_i;
    wire rgb_c_2;
    wire rgb_c_1;
    wire M_this_vram_read_data_0;
    wire M_this_vram_read_data_3;
    wire M_this_vram_read_data_2;
    wire M_this_vram_read_data_1;
    wire \this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ;
    wire \this_vga_ramdac.i2_mux ;
    wire \this_vga_ramdac.N_1764_reto ;
    wire \this_vga_ramdac.m16 ;
    wire \this_vga_ramdac.N_1765_reto ;
    wire port_clk_c;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire \this_vga_ramdac.N_24_mux ;
    wire \this_vga_ramdac.N_1762_reto ;
    wire \this_vga_ramdac.m6 ;
    wire \this_vga_ramdac.N_1763_reto ;
    wire \this_vga_ramdac.m19 ;
    wire \this_vga_ramdac.N_1766_reto ;
    wire \this_vga_signals.M_this_vga_signals_pixel_clk_0_0 ;
    wire M_pcounter_q_ret_2_RNIRAOL5;
    wire M_pcounter_q_ret_2_RNIRAOL5_cascade_;
    wire \this_vga_ramdac.i2_mux_0 ;
    wire \this_vga_ramdac.N_1767_reto ;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire M_this_vga_signals_address_2;
    wire M_this_vga_signals_address_1;
    wire \this_vga_signals.mult1_un75_sum_c2_0_cascade_ ;
    wire \this_vga_signals.if_m7_0_x4_0 ;
    wire \this_vga_signals.if_N_9_1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1 ;
    wire \this_vga_signals.if_m1_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_c3_cascade_ ;
    wire \this_vga_signals.N_2_7_0 ;
    wire \this_vga_signals.mult1_un75_sum_c2_0 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_c3 ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.mult1_un68_sum_axbxc3 ;
    wire \this_vga_signals.d_N_11 ;
    wire \this_vga_signals.d_N_12 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc1 ;
    wire M_this_vga_signals_address_5;
    wire M_this_vga_signals_address_4;
    wire \this_vga_signals.vaddress_1_0_5_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_cascade_ ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_cascade_ ;
    wire \this_vga_signals.if_i1_mux_0_cascade_ ;
    wire \this_vga_signals.g1_6_0 ;
    wire \this_vga_signals.mult1_un75_sum_c3_0_0 ;
    wire \this_vga_signals.if_m1_3 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3 ;
    wire \this_vga_signals.if_m1_3_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc2 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_i ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_i_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0 ;
    wire \this_vga_signals.if_N_2_1_0_0 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ;
    wire \this_vga_signals.g0_3_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb1 ;
    wire \this_vga_signals.N_5_1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0 ;
    wire \this_vga_signals.g1_2_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_2_0_0 ;
    wire \this_vga_signals.g1_3 ;
    wire \this_vga_signals.M_hcounter_q_RNI8OIBAZ0Z_3 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_0 ;
    wire \this_vga_signals.if_N_8_i_0 ;
    wire \this_vga_signals.g0_9_1_cascade_ ;
    wire \this_vga_signals.g0_12_x0 ;
    wire \this_vga_signals.g0_5_0 ;
    wire \this_vga_signals.N_6_0_cascade_ ;
    wire \this_vga_signals.N_5 ;
    wire \this_vga_signals.d_N_3_i_0_0_0 ;
    wire \this_vga_signals.M_pcounter_q_3_0_cascade_ ;
    wire \this_vga_signals.N_2_0 ;
    wire \this_vga_signals.N_2_0_cascade_ ;
    wire \this_vga_signals.M_pcounter_q_i_3_0 ;
    wire \this_vga_signals.N_3_0 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_pcounter_q_i_3_1 ;
    wire \this_vga_signals.M_pcounter_q_3_1 ;
    wire M_this_vga_signals_address_6;
    wire \this_vga_signals.mult1_un61_sum_c2_0 ;
    wire M_this_vga_signals_address_3;
    wire \this_vga_signals.vaddress_1_0_6 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.N_1_4_1_cascade_ ;
    wire \this_vga_signals.N_7 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_1_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_2 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_395_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0 ;
    wire \this_vga_signals.mult1_un54_sum_axb1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_1_cascade_ ;
    wire \this_vga_signals.g0_5_2_cascade_ ;
    wire \this_vga_signals.g1_2 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_1_x1 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_1 ;
    wire \this_vga_signals.N_3_1 ;
    wire \this_vga_signals.vaddress_1_5 ;
    wire \this_vga_signals.vaddress_1_6_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb1_1_0_1 ;
    wire \this_vga_signals.mult1_un61_sum_c3 ;
    wire \this_vga_signals.g0_12_x1 ;
    wire \this_vga_signals.g0_0_2_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_0 ;
    wire \this_vga_signals.g0_0_2 ;
    wire \this_vga_signals.vaddress_6_5 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_1_0_cascade_ ;
    wire \this_vga_signals.g0_0_2_0 ;
    wire \this_vga_signals.N_236 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_3_2 ;
    wire \this_vga_signals.N_3_2_1 ;
    wire \this_vga_signals.N_3_2_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire \this_vga_signals.mult1_un68_sum_axb2_1 ;
    wire \this_vga_signals.mult1_un68_sum_axb2_1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2 ;
    wire \this_vga_signals.SUM_3_i_0_0_3_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_0 ;
    wire this_vga_signals_hvisibility_i;
    wire \this_vga_signals.SUM_3_i_0_0_3 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ;
    wire M_this_vga_ramdac_en_0;
    wire \this_vga_signals.g0_7_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i_0_1_0 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ;
    wire \this_vga_signals.SUM_2_i_1_2_3 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i_0_0_cascade_ ;
    wire \this_vga_signals.SUM_2_i_1_0_3 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_0 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ;
    wire \this_vga_signals.vaddress_6_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i ;
    wire \this_vga_signals.g1_3_0 ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.vaddress_4_0_6 ;
    wire \this_vga_signals.vaddress_5_0_5 ;
    wire \this_vga_signals.g2_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb1_1 ;
    wire \this_vga_signals.g1_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_1_0_0 ;
    wire \this_vga_signals.N_5_i_5_cascade_ ;
    wire \this_vga_signals.N_20_0 ;
    wire \this_vga_signals.g1_1_1 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_0_0 ;
    wire \this_vga_signals.g0_2_x0_cascade_ ;
    wire \this_vga_signals.g1_0_0_0_cascade_ ;
    wire \this_vga_signals.N_5_i_5 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_ ;
    wire \this_vga_signals.g0_i_x2_0_2_0 ;
    wire \this_vga_signals.if_i4_mux_0_0_0 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_395 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_1_x0 ;
    wire \this_vga_signals.mult1_un61_sum_c3_1 ;
    wire \this_vga_signals.g0_2_x1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1 ;
    wire bfn_11_22_0_;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_11_23_0_;
    wire \this_vga_signals.un4_hsynclt8_0_cascade_ ;
    wire this_vga_signals_hsync_1_i;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.un3_hsynclt8_0 ;
    wire \this_vga_signals.un6_vvisibilitylto8_0_cascade_ ;
    wire \this_vga_signals.un6_vvisibilitylt9_0_cascade_ ;
    wire \this_vga_signals.vvisibility ;
    wire \this_vga_signals.g0_7_0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_0 ;
    wire \this_vga_signals.M_vcounter_q_7_repZ0Z1 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_8_repZ0Z1 ;
    wire \this_vga_signals.vaddress_2_6 ;
    wire \this_vga_signals.vaddress_2_5 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_2_0_1_0 ;
    wire \this_vga_signals.g0_22_1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb1_0_0_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0 ;
    wire \this_vga_signals.vaddress_5_5_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb1_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_1_0_0_0 ;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.vaddress_2_0_6 ;
    wire \this_vga_signals.g2_1 ;
    wire \this_vga_signals.if_N_5 ;
    wire \this_vga_signals.vaddress_4_5 ;
    wire \this_vga_signals.vaddress_3_6 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0 ;
    wire \this_vga_signals.vaddress_0_5_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i ;
    wire \this_vga_signals.mult1_un54_sum_axb1_0_cascade_ ;
    wire \this_vga_signals.g2 ;
    wire \this_vga_signals.g1 ;
    wire \this_vga_signals.vaddress_0_6 ;
    wire \this_vga_signals.g1_0_2 ;
    wire \this_vga_signals.g0_31_1 ;
    wire \this_vga_signals.g1_0_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_N_2L1 ;
    wire \this_vga_signals.N_5_1_0_0 ;
    wire \this_vga_signals.vsync_1_3 ;
    wire this_vga_signals_vsync_1_i;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.M_hcounter_d7lto7_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.un2_vsynclt8 ;
    wire \this_vga_signals.N_340_1 ;
    wire \this_vga_signals.vsync_1_2 ;
    wire bfn_13_17_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire bfn_13_18_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.vaddress_5_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.vaddress_3_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire \this_vga_signals.N_340_0_g ;
    wire \this_vga_signals.N_515_g ;
    wire \this_vga_signals.M_vcounter_q_5_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z1 ;
    wire \this_vga_signals.vaddress_5 ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z2 ;
    wire \this_vga_signals.vaddress_4_6 ;
    wire \this_vga_signals.M_vcounter_d7lto8_1_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire M_this_delay_clk_out_0;
    wire port_enb_c;
    wire this_start_data_delay_M_last_q;
    wire \this_vga_signals.vaddress_ac0_9_0_a0_0 ;
    wire \this_vga_signals.un6_vvisibilitylt9_0 ;
    wire \this_vga_signals.vaddress_c2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire \this_vga_signals.g1_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_d7lt8_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.un4_lvisibility_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire \this_vga_signals.line_clk_1 ;
    wire \this_vga_signals.un4_lvisibility_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.g0_0 ;
    wire N_206_cascade_;
    wire N_207;
    wire M_this_state_q_srsts_0_a2_1_4;
    wire port_dmab_c;
    wire port_dmab_c_i;
    wire M_this_ppu_vga_is_drawing_0;
    wire \this_ppu.M_line_clk_out_0_cascade_ ;
    wire M_this_sprites_address_q_3_ns_1_5;
    wire M_this_sprites_address_q_3_ns_1_4;
    wire M_this_sprites_address_q_3_ns_1_7_cascade_;
    wire bfn_15_22_0_;
    wire un1_M_this_sprites_address_q_cry_0;
    wire un1_M_this_sprites_address_q_cry_1;
    wire un1_M_this_sprites_address_q_cry_2;
    wire M_this_sprites_address_qZ0Z_4;
    wire M_this_sprites_address_q_RNO_1Z0Z_4;
    wire un1_M_this_sprites_address_q_cry_3;
    wire M_this_sprites_address_qZ0Z_5;
    wire M_this_sprites_address_q_RNO_1Z0Z_5;
    wire un1_M_this_sprites_address_q_cry_4;
    wire un1_M_this_sprites_address_q_cry_5;
    wire M_this_sprites_address_qZ0Z_7;
    wire M_this_sprites_address_q_RNO_1Z0Z_7;
    wire un1_M_this_sprites_address_q_cry_6;
    wire un1_M_this_sprites_address_q_cry_7;
    wire bfn_15_23_0_;
    wire un1_M_this_sprites_address_q_cry_8;
    wire un1_M_this_sprites_address_q_cry_9;
    wire un1_M_this_sprites_address_q_cry_10;
    wire un1_M_this_sprites_address_q_cry_11;
    wire un1_M_this_sprites_address_q_cry_12;
    wire M_this_sprites_address_q_RNO_1Z0Z_8;
    wire M_this_sprites_address_q_3_ns_1_8_cascade_;
    wire M_this_sprites_address_qZ0Z_8;
    wire \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_11 ;
    wire un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0;
    wire \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_12 ;
    wire un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0;
    wire M_this_sprites_address_q_RNO_1Z0Z_1;
    wire \this_vga_signals.un1_M_hcounter_d7_1_0_cascade_ ;
    wire \this_vga_signals.M_lcounter_qZ0Z_0 ;
    wire \this_vga_signals.un1_M_hcounter_d7_1_0 ;
    wire \this_vga_signals.CO0_cascade_ ;
    wire \this_vga_signals.M_lcounter_qZ0Z_1 ;
    wire \this_ppu.M_line_clk_out_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire M_counter_q_RNIFKS8_1;
    wire M_counter_q_RNIFKS8_1_cascade_;
    wire \this_vga_signals.M_hcounter_d7_0 ;
    wire M_this_state_q_nss_0;
    wire \this_pixel_clk.M_counter_q_i_1 ;
    wire M_this_state_q_srsts_i_1_2;
    wire port_rw_in;
    wire N_171_0_cascade_;
    wire N_176_0;
    wire M_this_state_qZ0Z_4;
    wire N_153_0;
    wire M_this_sprites_address_q_RNO_1Z0Z_2;
    wire M_this_sprites_address_q_RNO_1Z0Z_9;
    wire un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0;
    wire M_this_sprites_address_q_3_ns_1_6;
    wire M_this_sprites_address_q_RNO_1Z0Z_6;
    wire M_this_sprites_address_qZ0Z_6;
    wire M_this_sprites_address_qZ0Z_9;
    wire M_this_sprites_address_q_3_ns_1_9;
    wire M_this_sprites_address_qZ0Z_1;
    wire M_this_sprites_address_q_3_ns_1_1;
    wire \this_ppu.un1_M_haddress_q_c3_cascade_ ;
    wire \this_ppu.M_haddress_d8lto6_4 ;
    wire \this_ppu.un1_M_line_clk_out_ns_1_0 ;
    wire M_this_vga_signals_line_clk_0;
    wire \this_ppu.line_clk.M_last_qZ0 ;
    wire \this_vga_signals.M_vcounter_d8 ;
    wire \this_vga_signals.M_vcounter_q_249_0 ;
    wire \this_vga_signals.M_vcounter_q_esr_RNIRO2H5Z0Z_9 ;
    wire M_this_sprites_address_q_RNO_1Z0Z_0;
    wire \this_pixel_clk.M_counter_qZ0Z_0 ;
    wire M_this_sprites_address_qZ0Z_0;
    wire M_this_sprites_address_q_3_ns_1_0;
    wire M_this_state_q_srsts_i_a2_1_8_1;
    wire M_this_state_q_srsts_i_a2_1_7_1_cascade_;
    wire M_this_state_q_srsts_i_a2_1_9_1;
    wire M_this_state_q_srsts_i_a2_1_6_1;
    wire M_this_data_count_qZ0Z_0;
    wire bfn_17_23_0_;
    wire M_this_data_count_qZ0Z_1;
    wire un1_M_this_data_count_q_cry_0;
    wire M_this_data_count_qZ0Z_2;
    wire un1_M_this_data_count_q_cry_1;
    wire M_this_data_count_qZ0Z_3;
    wire un1_M_this_data_count_q_cry_2;
    wire M_this_data_count_qZ0Z_4;
    wire un1_M_this_data_count_q_cry_3;
    wire M_this_data_count_qZ0Z_5;
    wire un1_M_this_data_count_q_cry_4;
    wire M_this_data_count_qZ0Z_6;
    wire un1_M_this_data_count_q_cry_5;
    wire M_this_data_count_qZ0Z_7;
    wire un1_M_this_data_count_q_cry_6;
    wire un1_M_this_data_count_q_cry_7;
    wire M_this_data_count_qZ0Z_8;
    wire bfn_17_24_0_;
    wire M_this_data_count_qZ0Z_9;
    wire un1_M_this_data_count_q_cry_8;
    wire M_this_data_count_qZ0Z_10;
    wire un1_M_this_data_count_q_cry_9;
    wire M_this_data_count_qZ0Z_11;
    wire un1_M_this_data_count_q_cry_10;
    wire M_this_data_count_qZ0Z_12;
    wire un1_M_this_data_count_q_cry_11;
    wire M_this_state_q_RNI20CEZ0Z_0;
    wire un1_M_this_data_count_q_cry_12;
    wire un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO;
    wire un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO;
    wire bfn_17_25_0_;
    wire M_this_data_count_qZ0Z_13;
    wire \this_ppu.un1_M_haddress_q_c2_cascade_ ;
    wire \this_ppu.un1_M_haddress_q_c5_cascade_ ;
    wire \this_ppu.un1_M_haddress_q_c5 ;
    wire \this_ppu.un1_M_haddress_q_c2 ;
    wire \this_ppu.un1_M_vaddress_q_c1 ;
    wire port_address_in_0;
    wire port_address_in_1;
    wire N_218;
    wire N_204;
    wire N_202;
    wire M_this_state_qZ0Z_6;
    wire N_233;
    wire M_this_start_address_delay_out_0;
    wire M_this_state_q_srsts_i_1_1_cascade_;
    wire M_this_state_qZ0Z_1;
    wire \this_ppu.N_250_1 ;
    wire \this_ppu.M_last_q_RNI5NOQ4 ;
    wire \this_ppu.un1_M_vaddress_q_c3 ;
    wire \this_ppu.un1_M_vaddress_q_c5 ;
    wire \this_ppu.N_258_1 ;
    wire \this_ppu.un1_M_vaddress_q_c5_cascade_ ;
    wire \this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_13 ;
    wire M_this_sprites_address_qZ0Z_2;
    wire M_this_sprites_address_q_3_ns_1_2;
    wire M_this_ppu_vram_data_3;
    wire M_this_ppu_sprites_addr_1;
    wire M_this_sprites_address_q_3_ns_1_10;
    wire M_this_sprites_address_q_RNO_1Z0Z_10;
    wire M_this_sprites_address_qZ0Z_10;
    wire M_this_state_qZ0Z_5;
    wire M_this_sprites_address_q_3_sm0_0;
    wire M_this_sprites_address_q_3_ns_1_3_cascade_;
    wire M_this_sprites_address_q_RNO_1Z0Z_3;
    wire M_this_sprites_address_qZ0Z_3;
    wire \this_sprites_ram.mem_out_bus5_3 ;
    wire \this_sprites_ram.mem_out_bus1_3 ;
    wire \this_sprites_ram.mem_out_bus3_3 ;
    wire \this_sprites_ram.mem_out_bus7_3 ;
    wire \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_3 ;
    wire this_sprites_ram_mem_N_102;
    wire M_this_ppu_vram_data_1;
    wire \this_sprites_ram.mem_out_bus2_1 ;
    wire \this_sprites_ram.mem_out_bus6_1 ;
    wire this_sprites_ram_mem_N_91;
    wire \this_sprites_ram.mem_out_bus4_1 ;
    wire \this_sprites_ram.mem_out_bus0_1 ;
    wire \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_1 ;
    wire M_this_ppu_vram_addr_1;
    wire bfn_21_17_0_;
    wire M_this_ppu_vram_addr_2;
    wire M_this_ppu_sprites_addr_2;
    wire \this_ppu.sprites_addr_cry_1 ;
    wire M_this_ppu_vram_addr_3;
    wire M_this_ppu_sprites_addr_3;
    wire \this_ppu.sprites_addr_cry_2 ;
    wire M_this_ppu_vram_addr_4;
    wire M_this_ppu_sprites_addr_4;
    wire \this_ppu.sprites_addr_cry_3 ;
    wire M_this_ppu_vram_addr_5;
    wire M_this_ppu_sprites_addr_5;
    wire \this_ppu.sprites_addr_cry_4 ;
    wire M_this_ppu_vram_addr_6;
    wire M_this_ppu_sprites_addr_6;
    wire \this_ppu.sprites_addr_cry_5 ;
    wire M_this_ppu_vram_addr_7;
    wire M_this_ppu_sprites_addr_7;
    wire \this_ppu.sprites_addr_cry_6 ;
    wire \this_ppu.M_vaddress_qZ0Z_1 ;
    wire M_this_ppu_sprites_addr_8;
    wire \this_ppu.sprites_addr_cry_7 ;
    wire \this_ppu.sprites_addr_cry_8 ;
    wire \this_ppu.M_vaddress_qZ1Z_2 ;
    wire M_this_ppu_sprites_addr_9;
    wire bfn_21_18_0_;
    wire \this_ppu.M_vaddress_qZ0Z_3 ;
    wire M_this_ppu_sprites_addr_10;
    wire \this_ppu.sprites_addr_cry_9 ;
    wire \this_ppu.M_vaddress_qZ1Z_4 ;
    wire \this_ppu.sprites_addr_cry_10 ;
    wire \this_ppu.M_vaddress_qZ0Z_5 ;
    wire \this_ppu.sprites_addr_cry_11 ;
    wire \this_ppu.M_vaddress_qZ0Z_6 ;
    wire \this_ppu.sprites_addr_cry_12 ;
    wire M_this_ppu_vram_addr_0;
    wire M_this_ppu_vram_addr_i_0;
    wire \this_sprites_ram.mem_out_bus5_1 ;
    wire \this_sprites_ram.mem_out_bus1_1 ;
    wire \this_sprites_ram.mem_out_bus7_1 ;
    wire \this_sprites_ram.mem_out_bus3_1 ;
    wire \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_1_cascade_ ;
    wire this_sprites_ram_mem_N_88;
    wire \this_sprites_ram.mem_WE_14 ;
    wire \this_sprites_ram.mem_out_bus2_3 ;
    wire \this_sprites_ram.mem_out_bus6_3 ;
    wire this_sprites_ram_mem_N_105;
    wire N_200;
    wire M_this_ppu_vram_data_2;
    wire M_this_ppu_vram_en_0;
    wire this_sprites_ram_mem_radreg_11;
    wire M_this_ppu_vram_data_0;
    wire \this_sprites_ram.mem_out_bus4_3 ;
    wire \this_sprites_ram.mem_out_bus0_3 ;
    wire \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_3 ;
    wire M_this_state_qZ0Z_7;
    wire N_170_0;
    wire \this_sprites_ram.mem_WE_0 ;
    wire \this_sprites_ram.mem_out_bus4_2 ;
    wire \this_sprites_ram.mem_out_bus0_2 ;
    wire \this_sprites_ram.mem_out_bus6_2 ;
    wire \this_sprites_ram.mem_out_bus2_2 ;
    wire \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_2_cascade_ ;
    wire this_sprites_ram_mem_N_98;
    wire \this_sprites_ram.mem_out_bus5_0 ;
    wire \this_sprites_ram.mem_out_bus1_0 ;
    wire \this_sprites_ram.mem_out_bus3_0 ;
    wire \this_sprites_ram.mem_out_bus7_0 ;
    wire \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_0_cascade_ ;
    wire this_sprites_ram_mem_N_109;
    wire \this_sprites_ram.mem_out_bus0_0 ;
    wire \this_sprites_ram.mem_out_bus4_0 ;
    wire \this_sprites_ram.mem_out_bus6_0 ;
    wire \this_sprites_ram.mem_DOUT_3_i_m2_ns_1_0_cascade_ ;
    wire \this_sprites_ram.mem_out_bus2_0 ;
    wire this_sprites_ram_mem_N_112;
    wire \this_sprites_ram.mem_WE_10 ;
    wire \this_sprites_ram.mem_WE_8 ;
    wire \this_sprites_ram.mem_WE_12 ;
    wire \this_sprites_ram.mem_out_bus5_2 ;
    wire \this_sprites_ram.mem_radregZ0Z_13 ;
    wire \this_sprites_ram.mem_out_bus1_2 ;
    wire \this_sprites_ram.mem_out_bus7_2 ;
    wire \this_sprites_ram.mem_out_bus3_2 ;
    wire \this_sprites_ram.mem_DOUT_6_i_m2_ns_1_2_cascade_ ;
    wire \this_sprites_ram.mem_radregZ0Z_12 ;
    wire this_sprites_ram_mem_N_95;
    wire \this_sprites_ram.mem_WE_6 ;
    wire \this_sprites_ram.mem_WE_4 ;
    wire M_this_state_qZ0Z_2;
    wire M_this_start_data_delay_out_0;
    wire port_data_c_0;
    wire port_data_c_4;
    wire M_this_sprites_ram_write_data_0_sqmuxa_cascade_;
    wire M_this_sprites_ram_write_data_0_i_0;
    wire port_data_c_3;
    wire port_data_c_7;
    wire M_this_sprites_ram_write_data_0_i_3;
    wire port_data_c_2;
    wire port_data_c_6;
    wire M_this_sprites_ram_write_data_0_i_2;
    wire port_data_c_1;
    wire un1_M_this_state_q_2_0;
    wire port_data_c_5;
    wire M_this_sprites_ram_write_data_0_sqmuxa;
    wire M_this_sprites_ram_write_data_0_i_1;
    wire M_this_sprites_address_qZ0Z_12;
    wire M_this_sprites_ram_write_en_1_0_0;
    wire M_this_sprites_address_qZ0Z_13;
    wire M_this_sprites_address_qZ0Z_11;
    wire \this_sprites_ram.mem_WE_2 ;
    wire M_this_state_qZ0Z_3;
    wire M_this_external_address_qZ0Z_0;
    wire bfn_30_23_0_;
    wire M_this_external_address_qZ0Z_1;
    wire un1_M_this_external_address_q_cry_0;
    wire M_this_external_address_qZ0Z_2;
    wire un1_M_this_external_address_q_cry_1;
    wire M_this_external_address_qZ0Z_3;
    wire un1_M_this_external_address_q_cry_2;
    wire M_this_external_address_qZ0Z_4;
    wire un1_M_this_external_address_q_cry_3;
    wire M_this_external_address_qZ0Z_5;
    wire un1_M_this_external_address_q_cry_4;
    wire M_this_external_address_qZ0Z_6;
    wire un1_M_this_external_address_q_cry_5;
    wire M_this_external_address_qZ0Z_7;
    wire un1_M_this_external_address_q_cry_6;
    wire un1_M_this_external_address_q_cry_7;
    wire M_this_external_address_qZ0Z_8;
    wire bfn_30_24_0_;
    wire M_this_external_address_qZ0Z_9;
    wire un1_M_this_external_address_q_cry_8;
    wire M_this_external_address_qZ0Z_10;
    wire un1_M_this_external_address_q_cry_9;
    wire M_this_external_address_qZ0Z_11;
    wire un1_M_this_external_address_q_cry_10;
    wire M_this_external_address_qZ0Z_12;
    wire un1_M_this_external_address_q_cry_11;
    wire M_this_external_address_qZ0Z_13;
    wire un1_M_this_external_address_q_cry_12;
    wire M_this_external_address_qZ0Z_14;
    wire un1_M_this_external_address_q_cry_13;
    wire M_this_state_qZ0Z_0;
    wire un1_M_this_external_address_q_cry_14;
    wire M_this_external_address_qZ0Z_15;
    wire clk_0_c_g;
    wire M_this_state_q_nss_g_0;
    wire port_address_in_3;
    wire port_address_in_4;
    wire port_address_in_5;
    wire port_address_in_2;
    wire port_address_in_7;
    wire M_this_state_d36_2_0_3_cascade_;
    wire port_address_in_6;
    wire M_this_state_d37_1;
    wire _gnd_net_;

    defparam \this_sprites_ram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,\this_sprites_ram.mem_out_bus0_1 ,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,\this_sprites_ram.mem_out_bus0_0 ,dangling_wire_11,dangling_wire_12,dangling_wire_13}),
            .RADDR({N__19100,N__17630,N__17771,N__17918,N__18083,N__18242,N__18395,N__18557,N__16985,N__16664,N__18848}),
            .WADDR({N__16541,N__14810,N__14030,N__13604,N__14927,N__13742,N__13868,N__17417,N__16817,N__14672,N__15374}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,N__21410,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__20072,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .RCLKE(),
            .RCLK(N__22166),
            .RE(N__15906),
            .WCLKE(N__18677),
            .WCLK(N__22167),
            .WE(N__15908));
    defparam \this_sprites_ram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,\this_sprites_ram.mem_out_bus0_3 ,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,\this_sprites_ram.mem_out_bus0_2 ,dangling_wire_55,dangling_wire_56,dangling_wire_57}),
            .RADDR({N__19094,N__17624,N__17765,N__17912,N__18077,N__18236,N__18389,N__18551,N__16979,N__16658,N__18842}),
            .WADDR({N__16535,N__14804,N__14024,N__13598,N__14921,N__13736,N__13862,N__17411,N__16811,N__14666,N__15368}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,N__19922,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,N__19748,dangling_wire_85,dangling_wire_86,dangling_wire_87}),
            .RCLKE(),
            .RCLK(N__22168),
            .RE(N__15905),
            .WCLKE(N__18670),
            .WCLK(N__22169),
            .WE(N__15907));
    defparam \this_sprites_ram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,\this_sprites_ram.mem_out_bus1_1 ,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,\this_sprites_ram.mem_out_bus1_0 ,dangling_wire_99,dangling_wire_100,dangling_wire_101}),
            .RADDR({N__19088,N__17618,N__17759,N__17906,N__18071,N__18230,N__18383,N__18545,N__16973,N__16652,N__18836}),
            .WADDR({N__16529,N__14798,N__14018,N__13592,N__14915,N__13730,N__13856,N__17405,N__16805,N__14660,N__15362}),
            .MASK({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .WDATA({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__21406,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__20068,dangling_wire_129,dangling_wire_130,dangling_wire_131}),
            .RCLKE(),
            .RCLK(N__22170),
            .RE(N__15889),
            .WCLKE(N__19445),
            .WCLK(N__22171),
            .WE(N__15903));
    defparam \this_sprites_ram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,\this_sprites_ram.mem_out_bus1_3 ,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,\this_sprites_ram.mem_out_bus1_2 ,dangling_wire_143,dangling_wire_144,dangling_wire_145}),
            .RADDR({N__19082,N__17612,N__17753,N__17900,N__18065,N__18224,N__18377,N__18539,N__16967,N__16646,N__18830}),
            .WADDR({N__16523,N__14792,N__14012,N__13586,N__14909,N__13724,N__13850,N__17399,N__16799,N__14654,N__15356}),
            .MASK({dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161}),
            .WDATA({dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,N__19918,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,N__19744,dangling_wire_173,dangling_wire_174,dangling_wire_175}),
            .RCLKE(),
            .RCLK(N__22172),
            .RE(N__15888),
            .WCLKE(N__19441),
            .WCLK(N__22173),
            .WE(N__15902));
    defparam \this_sprites_ram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,\this_sprites_ram.mem_out_bus2_1 ,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,\this_sprites_ram.mem_out_bus2_0 ,dangling_wire_187,dangling_wire_188,dangling_wire_189}),
            .RADDR({N__19076,N__17606,N__17747,N__17894,N__18059,N__18218,N__18371,N__18533,N__16961,N__16640,N__18824}),
            .WADDR({N__16517,N__14786,N__14006,N__13580,N__14903,N__13718,N__13844,N__17393,N__16793,N__14648,N__15350}),
            .MASK({dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205}),
            .WDATA({dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,N__21399,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,N__20061,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .RCLKE(),
            .RCLK(N__22179),
            .RE(N__15854),
            .WCLKE(N__19487),
            .WCLK(N__22178),
            .WE(N__15876));
    defparam \this_sprites_ram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,\this_sprites_ram.mem_out_bus2_3 ,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,\this_sprites_ram.mem_out_bus2_2 ,dangling_wire_231,dangling_wire_232,dangling_wire_233}),
            .RADDR({N__19070,N__17600,N__17741,N__17888,N__18053,N__18212,N__18365,N__18527,N__16955,N__16634,N__18818}),
            .WADDR({N__16511,N__14780,N__14000,N__13574,N__14897,N__13712,N__13838,N__17387,N__16787,N__14642,N__15344}),
            .MASK({dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249}),
            .WDATA({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,N__19911,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,N__19736,dangling_wire_261,dangling_wire_262,dangling_wire_263}),
            .RCLKE(),
            .RCLK(N__22186),
            .RE(N__15853),
            .WCLKE(N__19486),
            .WCLK(N__22187),
            .WE(N__15875));
    defparam \this_sprites_ram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,\this_sprites_ram.mem_out_bus3_1 ,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,\this_sprites_ram.mem_out_bus3_0 ,dangling_wire_275,dangling_wire_276,dangling_wire_277}),
            .RADDR({N__19064,N__17594,N__17735,N__17882,N__18047,N__18206,N__18359,N__18521,N__16949,N__16628,N__18812}),
            .WADDR({N__16505,N__14774,N__13994,N__13568,N__14891,N__13706,N__13832,N__17381,N__16781,N__14636,N__15338}),
            .MASK({dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293}),
            .WDATA({dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,N__21390,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,N__20051,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .RCLKE(),
            .RCLK(N__22199),
            .RE(N__15799),
            .WCLKE(N__19459),
            .WCLK(N__22200),
            .WE(N__15848));
    defparam \this_sprites_ram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,\this_sprites_ram.mem_out_bus3_3 ,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,\this_sprites_ram.mem_out_bus3_2 ,dangling_wire_319,dangling_wire_320,dangling_wire_321}),
            .RADDR({N__19058,N__17588,N__17729,N__17876,N__18041,N__18200,N__18353,N__18515,N__16943,N__16622,N__18806}),
            .WADDR({N__16499,N__14768,N__13988,N__13562,N__14885,N__13700,N__13826,N__17375,N__16775,N__14630,N__15332}),
            .MASK({dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337}),
            .WDATA({dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,N__19902,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,N__19723,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .RCLKE(),
            .RCLK(N__22209),
            .RE(N__15798),
            .WCLKE(N__19463),
            .WCLK(N__22210),
            .WE(N__15790));
    defparam \this_sprites_ram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,\this_sprites_ram.mem_out_bus4_1 ,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,\this_sprites_ram.mem_out_bus4_0 ,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .RADDR({N__19052,N__17582,N__17723,N__17870,N__18035,N__18194,N__18347,N__18509,N__16937,N__16616,N__18800}),
            .WADDR({N__16493,N__14762,N__13982,N__13556,N__14879,N__13694,N__13820,N__17369,N__16769,N__14624,N__15326}),
            .MASK({dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381}),
            .WDATA({dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,N__21380,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,N__20038,dangling_wire_393,dangling_wire_394,dangling_wire_395}),
            .RCLKE(),
            .RCLK(N__22219),
            .RE(N__15734),
            .WCLKE(N__20431),
            .WCLK(N__22220),
            .WE(N__15786));
    defparam \this_sprites_ram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,\this_sprites_ram.mem_out_bus4_3 ,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,\this_sprites_ram.mem_out_bus4_2 ,dangling_wire_407,dangling_wire_408,dangling_wire_409}),
            .RADDR({N__19046,N__17576,N__17717,N__17864,N__18029,N__18188,N__18341,N__18503,N__16931,N__16610,N__18794}),
            .WADDR({N__16487,N__14756,N__13976,N__13550,N__14873,N__13688,N__13814,N__17363,N__16763,N__14618,N__15320}),
            .MASK({dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425}),
            .WDATA({dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,N__19888,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,N__19708,dangling_wire_437,dangling_wire_438,dangling_wire_439}),
            .RCLKE(),
            .RCLK(N__22225),
            .RE(N__15733),
            .WCLKE(N__20435),
            .WCLK(N__22226),
            .WE(N__15688));
    defparam \this_sprites_ram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,\this_sprites_ram.mem_out_bus5_1 ,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,\this_sprites_ram.mem_out_bus5_0 ,dangling_wire_451,dangling_wire_452,dangling_wire_453}),
            .RADDR({N__19040,N__17570,N__17711,N__17858,N__18023,N__18182,N__18335,N__18497,N__16925,N__16604,N__18788}),
            .WADDR({N__16481,N__14750,N__13970,N__13544,N__14867,N__13682,N__13808,N__17357,N__16757,N__14612,N__15314}),
            .MASK({dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469}),
            .WDATA({dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,N__21367,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,N__20003,dangling_wire_481,dangling_wire_482,dangling_wire_483}),
            .RCLKE(),
            .RCLK(N__22227),
            .RE(N__15758),
            .WCLKE(N__20413),
            .WCLK(N__22228),
            .WE(N__15774));
    defparam \this_sprites_ram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,\this_sprites_ram.mem_out_bus5_3 ,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,\this_sprites_ram.mem_out_bus5_2 ,dangling_wire_495,dangling_wire_496,dangling_wire_497}),
            .RADDR({N__19034,N__17564,N__17705,N__17852,N__18017,N__18176,N__18329,N__18491,N__16919,N__16598,N__18782}),
            .WADDR({N__16475,N__14744,N__13964,N__13538,N__14861,N__13676,N__13802,N__17351,N__16751,N__14606,N__15308}),
            .MASK({dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513}),
            .WDATA({dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,N__19862,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,N__19694,dangling_wire_525,dangling_wire_526,dangling_wire_527}),
            .RCLKE(),
            .RCLK(N__22233),
            .RE(N__15759),
            .WCLKE(N__20414),
            .WCLK(N__22234),
            .WE(N__15840));
    defparam \this_sprites_ram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,\this_sprites_ram.mem_out_bus6_1 ,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,\this_sprites_ram.mem_out_bus6_0 ,dangling_wire_539,dangling_wire_540,dangling_wire_541}),
            .RADDR({N__19028,N__17558,N__17699,N__17846,N__18011,N__18170,N__18323,N__18485,N__16913,N__16592,N__18776}),
            .WADDR({N__16469,N__14738,N__13958,N__13532,N__14855,N__13670,N__13796,N__17345,N__16745,N__14600,N__15302}),
            .MASK({dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557}),
            .WDATA({dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,N__21376,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,N__20034,dangling_wire_569,dangling_wire_570,dangling_wire_571}),
            .RCLKE(),
            .RCLK(N__22235),
            .RE(N__15829),
            .WCLKE(N__20989),
            .WCLK(N__22236),
            .WE(N__15841));
    defparam \this_sprites_ram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,\this_sprites_ram.mem_out_bus6_3 ,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,\this_sprites_ram.mem_out_bus6_2 ,dangling_wire_583,dangling_wire_584,dangling_wire_585}),
            .RADDR({N__19022,N__17552,N__17693,N__17840,N__18005,N__18164,N__18317,N__18479,N__16907,N__16586,N__18770}),
            .WADDR({N__16463,N__14732,N__13952,N__13526,N__14849,N__13664,N__13790,N__17339,N__16739,N__14594,N__15296}),
            .MASK({dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601}),
            .WDATA({dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,N__19889,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,N__19732,dangling_wire_613,dangling_wire_614,dangling_wire_615}),
            .RCLKE(),
            .RCLK(N__22237),
            .RE(N__15830),
            .WCLKE(N__20993),
            .WCLK(N__22238),
            .WE(N__15880));
    defparam \this_sprites_ram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,\this_sprites_ram.mem_out_bus7_1 ,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,\this_sprites_ram.mem_out_bus7_0 ,dangling_wire_627,dangling_wire_628,dangling_wire_629}),
            .RADDR({N__19016,N__17546,N__17687,N__17834,N__17999,N__18158,N__18311,N__18473,N__16901,N__16580,N__18764}),
            .WADDR({N__16457,N__14726,N__13946,N__13520,N__14843,N__13658,N__13784,N__17333,N__16733,N__14588,N__15290}),
            .MASK({dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645}),
            .WDATA({dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,N__21389,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,N__20050,dangling_wire_657,dangling_wire_658,dangling_wire_659}),
            .RCLKE(),
            .RCLK(N__22240),
            .RE(N__15881),
            .WCLKE(N__19147),
            .WCLK(N__22241),
            .WE(N__15883));
    defparam \this_sprites_ram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,\this_sprites_ram.mem_out_bus7_3 ,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,\this_sprites_ram.mem_out_bus7_2 ,dangling_wire_671,dangling_wire_672,dangling_wire_673}),
            .RADDR({N__19010,N__17540,N__17681,N__17828,N__17993,N__18152,N__18305,N__18467,N__16895,N__16574,N__18758}),
            .WADDR({N__16451,N__14720,N__13940,N__13514,N__14837,N__13652,N__13778,N__17327,N__16727,N__14582,N__15284}),
            .MASK({dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689}),
            .WDATA({dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,N__19901,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,N__19743,dangling_wire_701,dangling_wire_702,dangling_wire_703}),
            .RCLKE(),
            .RCLK(N__22243),
            .RE(N__15882),
            .WCLKE(N__19151),
            .WCLK(N__22244),
            .WE(N__15904));
    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,dangling_wire_709,dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,M_this_vram_read_data_3,M_this_vram_read_data_2,M_this_vram_read_data_1,M_this_vram_read_data_0}),
            .RADDR({dangling_wire_716,dangling_wire_717,dangling_wire_718,N__8381,N__8672,N__8243,N__8231,N__8630,N__8048,N__8036,N__8339}),
            .WADDR({dangling_wire_719,dangling_wire_720,dangling_wire_721,N__17966,N__18128,N__18281,N__18443,N__18602,N__17045,N__17114,N__18920}),
            .MASK({dangling_wire_722,dangling_wire_723,dangling_wire_724,dangling_wire_725,dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737}),
            .WDATA({dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741,dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,N__16676,N__19409,N__17210,N__19229}),
            .RCLKE(),
            .RCLK(N__22175),
            .RE(N__15887),
            .WCLKE(N__19386),
            .WCLK(N__22174),
            .WE(N__15849));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__22938),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__22940),
            .DIN(N__22939),
            .DOUT(N__22938),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__22940),
            .PADOUT(N__22939),
            .PADIN(N__22938),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__22929),
            .DIN(N__22928),
            .DOUT(N__22927),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__22929),
            .PADOUT(N__22928),
            .PADIN(N__22927),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__22920),
            .DIN(N__22919),
            .DOUT(N__22918),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__22920),
            .PADOUT(N__22919),
            .PADIN(N__22918),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__22911),
            .DIN(N__22910),
            .DOUT(N__22909),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__22911),
            .PADOUT(N__22910),
            .PADIN(N__22909),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__9443),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__22902),
            .DIN(N__22901),
            .DOUT(N__22900),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__22902),
            .PADOUT(N__22901),
            .PADIN(N__22900),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__10163),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__22893),
            .DIN(N__22892),
            .DOUT(N__22891),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__22893),
            .PADOUT(N__22892),
            .PADIN(N__22891),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__20837),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13042));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__22884),
            .DIN(N__22883),
            .DOUT(N__22882),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__22884),
            .PADOUT(N__22883),
            .PADIN(N__22882),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__20813),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13052));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__22875),
            .DIN(N__22874),
            .DOUT(N__22873),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__22875),
            .PADOUT(N__22874),
            .PADIN(N__22873),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__20789),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13099));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__22866),
            .DIN(N__22865),
            .DOUT(N__22864),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__22866),
            .PADOUT(N__22865),
            .PADIN(N__22864),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__20759),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13120));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__22857),
            .DIN(N__22856),
            .DOUT(N__22855),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__22857),
            .PADOUT(N__22856),
            .PADIN(N__22855),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__20735),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13035));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__22848),
            .DIN(N__22847),
            .DOUT(N__22846),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__22848),
            .PADOUT(N__22847),
            .PADIN(N__22846),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__20717),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13109));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__22839),
            .DIN(N__22838),
            .DOUT(N__22837),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__22839),
            .PADOUT(N__22838),
            .PADIN(N__22837),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__21734),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13124));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__22830),
            .DIN(N__22829),
            .DOUT(N__22828),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__22830),
            .PADOUT(N__22829),
            .PADIN(N__22828),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__21713),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13142));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__22821),
            .DIN(N__22820),
            .DOUT(N__22819),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__22821),
            .PADOUT(N__22820),
            .PADIN(N__22819),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21632),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13068));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__22812),
            .DIN(N__22811),
            .DOUT(N__22810),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__22812),
            .PADOUT(N__22811),
            .PADIN(N__22810),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21602),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13129));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__22803),
            .DIN(N__22802),
            .DOUT(N__22801),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__22803),
            .PADOUT(N__22802),
            .PADIN(N__22801),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21584),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13102));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__22794),
            .DIN(N__22793),
            .DOUT(N__22792),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__22794),
            .PADOUT(N__22793),
            .PADIN(N__22792),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21566),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13110));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__22785),
            .DIN(N__22784),
            .DOUT(N__22783),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__22785),
            .PADOUT(N__22784),
            .PADIN(N__22783),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22532),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13125));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__22776),
            .DIN(N__22775),
            .DOUT(N__22774),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__22776),
            .PADOUT(N__22775),
            .PADIN(N__22774),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22268),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13141));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__22767),
            .DIN(N__22766),
            .DOUT(N__22765),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__22767),
            .PADOUT(N__22766),
            .PADIN(N__22765),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21686),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13041));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__22758),
            .DIN(N__22757),
            .DOUT(N__22756),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__22758),
            .PADOUT(N__22757),
            .PADIN(N__22756),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21653),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13100));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__22749),
            .DIN(N__22748),
            .DOUT(N__22747),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__22749),
            .PADOUT(N__22748),
            .PADIN(N__22747),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__22740),
            .DIN(N__22739),
            .DOUT(N__22738),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__22740),
            .PADOUT(N__22739),
            .PADIN(N__22738),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__22731),
            .DIN(N__22730),
            .DOUT(N__22729),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__22731),
            .PADOUT(N__22730),
            .PADIN(N__22729),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__22722),
            .DIN(N__22721),
            .DOUT(N__22720),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__22722),
            .PADOUT(N__22721),
            .PADIN(N__22720),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__22713),
            .DIN(N__22712),
            .DOUT(N__22711),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__22713),
            .PADOUT(N__22712),
            .PADIN(N__22711),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__22704),
            .DIN(N__22703),
            .DOUT(N__22702),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__22704),
            .PADOUT(N__22703),
            .PADIN(N__22702),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__22695),
            .DIN(N__22694),
            .DOUT(N__22693),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__22695),
            .PADOUT(N__22694),
            .PADIN(N__22693),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__22686),
            .DIN(N__22685),
            .DOUT(N__22684),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__22686),
            .PADOUT(N__22685),
            .PADIN(N__22684),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_7_iopad (
            .OE(N__22677),
            .DIN(N__22676),
            .DOUT(N__22675),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_7_preio (
            .PADOEN(N__22677),
            .PADOUT(N__22676),
            .PADIN(N__22675),
            .CLOCKENABLE(),
            .DIN0(port_data_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__22668),
            .DIN(N__22667),
            .DOUT(N__22666),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__22668),
            .PADOUT(N__22667),
            .PADIN(N__22666),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7643),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__22659),
            .DIN(N__22658),
            .DOUT(N__22657),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__22659),
            .PADOUT(N__22658),
            .PADIN(N__22657),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13217),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__22650),
            .DIN(N__22649),
            .DOUT(N__22648),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__22650),
            .PADOUT(N__22649),
            .PADIN(N__22648),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__22641),
            .DIN(N__22640),
            .DOUT(N__22639),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__22641),
            .PADOUT(N__22640),
            .PADIN(N__22639),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7601),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__22632),
            .DIN(N__22631),
            .DOUT(N__22630),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__22632),
            .PADOUT(N__22631),
            .PADIN(N__22630),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__15797),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13101));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__22623),
            .DIN(N__22622),
            .DOUT(N__22621),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__22623),
            .PADOUT(N__22622),
            .PADIN(N__22621),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7637),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__22614),
            .DIN(N__22613),
            .DOUT(N__22612),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__22614),
            .PADOUT(N__22613),
            .PADIN(N__22612),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7814),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__22605),
            .DIN(N__22604),
            .DOUT(N__22603),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__22605),
            .PADOUT(N__22604),
            .PADIN(N__22603),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7829),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__22596),
            .DIN(N__22595),
            .DOUT(N__22594),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__22596),
            .PADOUT(N__22595),
            .PADIN(N__22594),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7589),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__22587),
            .DIN(N__22586),
            .DOUT(N__22585),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__22587),
            .PADOUT(N__22586),
            .PADIN(N__22585),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7619),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__22578),
            .DIN(N__22577),
            .DOUT(N__22576),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__22578),
            .PADOUT(N__22577),
            .PADIN(N__22576),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7577),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__22569),
            .DIN(N__22568),
            .DOUT(N__22567),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__22569),
            .PADOUT(N__22568),
            .PADIN(N__22567),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__22560),
            .DIN(N__22559),
            .DOUT(N__22558),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__22560),
            .PADOUT(N__22559),
            .PADIN(N__22558),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7841),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__22551),
            .DIN(N__22550),
            .DOUT(N__22549),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__22551),
            .PADOUT(N__22550),
            .PADIN(N__22549),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11210),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IoInMux I__5534 (
            .O(N__22532),
            .I(N__22529));
    LocalMux I__5533 (
            .O(N__22529),
            .I(N__22526));
    Span4Mux_s2_h I__5532 (
            .O(N__22526),
            .I(N__22523));
    Sp12to4 I__5531 (
            .O(N__22523),
            .I(N__22519));
    InMux I__5530 (
            .O(N__22522),
            .I(N__22516));
    Odrv12 I__5529 (
            .O(N__22519),
            .I(M_this_external_address_qZ0Z_14));
    LocalMux I__5528 (
            .O(N__22516),
            .I(M_this_external_address_qZ0Z_14));
    InMux I__5527 (
            .O(N__22511),
            .I(un1_M_this_external_address_q_cry_13));
    InMux I__5526 (
            .O(N__22508),
            .I(N__22493));
    InMux I__5525 (
            .O(N__22507),
            .I(N__22493));
    InMux I__5524 (
            .O(N__22506),
            .I(N__22493));
    InMux I__5523 (
            .O(N__22505),
            .I(N__22493));
    InMux I__5522 (
            .O(N__22504),
            .I(N__22493));
    LocalMux I__5521 (
            .O(N__22493),
            .I(N__22479));
    InMux I__5520 (
            .O(N__22492),
            .I(N__22472));
    InMux I__5519 (
            .O(N__22491),
            .I(N__22472));
    InMux I__5518 (
            .O(N__22490),
            .I(N__22472));
    InMux I__5517 (
            .O(N__22489),
            .I(N__22463));
    InMux I__5516 (
            .O(N__22488),
            .I(N__22463));
    InMux I__5515 (
            .O(N__22487),
            .I(N__22463));
    InMux I__5514 (
            .O(N__22486),
            .I(N__22463));
    InMux I__5513 (
            .O(N__22485),
            .I(N__22454));
    InMux I__5512 (
            .O(N__22484),
            .I(N__22454));
    InMux I__5511 (
            .O(N__22483),
            .I(N__22454));
    InMux I__5510 (
            .O(N__22482),
            .I(N__22454));
    Span4Mux_v I__5509 (
            .O(N__22479),
            .I(N__22444));
    LocalMux I__5508 (
            .O(N__22472),
            .I(N__22439));
    LocalMux I__5507 (
            .O(N__22463),
            .I(N__22439));
    LocalMux I__5506 (
            .O(N__22454),
            .I(N__22436));
    CascadeMux I__5505 (
            .O(N__22453),
            .I(N__22432));
    CascadeMux I__5504 (
            .O(N__22452),
            .I(N__22429));
    CascadeMux I__5503 (
            .O(N__22451),
            .I(N__22424));
    CascadeMux I__5502 (
            .O(N__22450),
            .I(N__22416));
    CascadeMux I__5501 (
            .O(N__22449),
            .I(N__22413));
    CascadeMux I__5500 (
            .O(N__22448),
            .I(N__22410));
    CascadeMux I__5499 (
            .O(N__22447),
            .I(N__22407));
    Span4Mux_s1_h I__5498 (
            .O(N__22444),
            .I(N__22400));
    Span4Mux_v I__5497 (
            .O(N__22439),
            .I(N__22400));
    Span4Mux_v I__5496 (
            .O(N__22436),
            .I(N__22400));
    InMux I__5495 (
            .O(N__22435),
            .I(N__22397));
    InMux I__5494 (
            .O(N__22432),
            .I(N__22392));
    InMux I__5493 (
            .O(N__22429),
            .I(N__22385));
    InMux I__5492 (
            .O(N__22428),
            .I(N__22385));
    InMux I__5491 (
            .O(N__22427),
            .I(N__22385));
    InMux I__5490 (
            .O(N__22424),
            .I(N__22382));
    InMux I__5489 (
            .O(N__22423),
            .I(N__22379));
    InMux I__5488 (
            .O(N__22422),
            .I(N__22376));
    CascadeMux I__5487 (
            .O(N__22421),
            .I(N__22372));
    CascadeMux I__5486 (
            .O(N__22420),
            .I(N__22369));
    CascadeMux I__5485 (
            .O(N__22419),
            .I(N__22366));
    InMux I__5484 (
            .O(N__22416),
            .I(N__22362));
    InMux I__5483 (
            .O(N__22413),
            .I(N__22357));
    InMux I__5482 (
            .O(N__22410),
            .I(N__22357));
    InMux I__5481 (
            .O(N__22407),
            .I(N__22354));
    Span4Mux_h I__5480 (
            .O(N__22400),
            .I(N__22351));
    LocalMux I__5479 (
            .O(N__22397),
            .I(N__22348));
    InMux I__5478 (
            .O(N__22396),
            .I(N__22343));
    InMux I__5477 (
            .O(N__22395),
            .I(N__22343));
    LocalMux I__5476 (
            .O(N__22392),
            .I(N__22338));
    LocalMux I__5475 (
            .O(N__22385),
            .I(N__22338));
    LocalMux I__5474 (
            .O(N__22382),
            .I(N__22333));
    LocalMux I__5473 (
            .O(N__22379),
            .I(N__22333));
    LocalMux I__5472 (
            .O(N__22376),
            .I(N__22330));
    InMux I__5471 (
            .O(N__22375),
            .I(N__22327));
    InMux I__5470 (
            .O(N__22372),
            .I(N__22324));
    InMux I__5469 (
            .O(N__22369),
            .I(N__22321));
    InMux I__5468 (
            .O(N__22366),
            .I(N__22316));
    InMux I__5467 (
            .O(N__22365),
            .I(N__22316));
    LocalMux I__5466 (
            .O(N__22362),
            .I(N__22309));
    LocalMux I__5465 (
            .O(N__22357),
            .I(N__22309));
    LocalMux I__5464 (
            .O(N__22354),
            .I(N__22309));
    Span4Mux_h I__5463 (
            .O(N__22351),
            .I(N__22306));
    Span4Mux_h I__5462 (
            .O(N__22348),
            .I(N__22301));
    LocalMux I__5461 (
            .O(N__22343),
            .I(N__22301));
    Span4Mux_v I__5460 (
            .O(N__22338),
            .I(N__22296));
    Span4Mux_v I__5459 (
            .O(N__22333),
            .I(N__22296));
    Span4Mux_h I__5458 (
            .O(N__22330),
            .I(N__22291));
    LocalMux I__5457 (
            .O(N__22327),
            .I(N__22291));
    LocalMux I__5456 (
            .O(N__22324),
            .I(N__22278));
    LocalMux I__5455 (
            .O(N__22321),
            .I(N__22278));
    LocalMux I__5454 (
            .O(N__22316),
            .I(N__22278));
    Span4Mux_v I__5453 (
            .O(N__22309),
            .I(N__22278));
    Span4Mux_h I__5452 (
            .O(N__22306),
            .I(N__22278));
    Span4Mux_v I__5451 (
            .O(N__22301),
            .I(N__22278));
    Odrv4 I__5450 (
            .O(N__22296),
            .I(M_this_state_qZ0Z_0));
    Odrv4 I__5449 (
            .O(N__22291),
            .I(M_this_state_qZ0Z_0));
    Odrv4 I__5448 (
            .O(N__22278),
            .I(M_this_state_qZ0Z_0));
    InMux I__5447 (
            .O(N__22271),
            .I(un1_M_this_external_address_q_cry_14));
    IoInMux I__5446 (
            .O(N__22268),
            .I(N__22265));
    LocalMux I__5445 (
            .O(N__22265),
            .I(N__22262));
    Span4Mux_s2_h I__5444 (
            .O(N__22262),
            .I(N__22259));
    Sp12to4 I__5443 (
            .O(N__22259),
            .I(N__22256));
    Span12Mux_v I__5442 (
            .O(N__22256),
            .I(N__22252));
    InMux I__5441 (
            .O(N__22255),
            .I(N__22249));
    Odrv12 I__5440 (
            .O(N__22252),
            .I(M_this_external_address_qZ0Z_15));
    LocalMux I__5439 (
            .O(N__22249),
            .I(M_this_external_address_qZ0Z_15));
    ClkMux I__5438 (
            .O(N__22244),
            .I(N__22007));
    ClkMux I__5437 (
            .O(N__22243),
            .I(N__22007));
    ClkMux I__5436 (
            .O(N__22242),
            .I(N__22007));
    ClkMux I__5435 (
            .O(N__22241),
            .I(N__22007));
    ClkMux I__5434 (
            .O(N__22240),
            .I(N__22007));
    ClkMux I__5433 (
            .O(N__22239),
            .I(N__22007));
    ClkMux I__5432 (
            .O(N__22238),
            .I(N__22007));
    ClkMux I__5431 (
            .O(N__22237),
            .I(N__22007));
    ClkMux I__5430 (
            .O(N__22236),
            .I(N__22007));
    ClkMux I__5429 (
            .O(N__22235),
            .I(N__22007));
    ClkMux I__5428 (
            .O(N__22234),
            .I(N__22007));
    ClkMux I__5427 (
            .O(N__22233),
            .I(N__22007));
    ClkMux I__5426 (
            .O(N__22232),
            .I(N__22007));
    ClkMux I__5425 (
            .O(N__22231),
            .I(N__22007));
    ClkMux I__5424 (
            .O(N__22230),
            .I(N__22007));
    ClkMux I__5423 (
            .O(N__22229),
            .I(N__22007));
    ClkMux I__5422 (
            .O(N__22228),
            .I(N__22007));
    ClkMux I__5421 (
            .O(N__22227),
            .I(N__22007));
    ClkMux I__5420 (
            .O(N__22226),
            .I(N__22007));
    ClkMux I__5419 (
            .O(N__22225),
            .I(N__22007));
    ClkMux I__5418 (
            .O(N__22224),
            .I(N__22007));
    ClkMux I__5417 (
            .O(N__22223),
            .I(N__22007));
    ClkMux I__5416 (
            .O(N__22222),
            .I(N__22007));
    ClkMux I__5415 (
            .O(N__22221),
            .I(N__22007));
    ClkMux I__5414 (
            .O(N__22220),
            .I(N__22007));
    ClkMux I__5413 (
            .O(N__22219),
            .I(N__22007));
    ClkMux I__5412 (
            .O(N__22218),
            .I(N__22007));
    ClkMux I__5411 (
            .O(N__22217),
            .I(N__22007));
    ClkMux I__5410 (
            .O(N__22216),
            .I(N__22007));
    ClkMux I__5409 (
            .O(N__22215),
            .I(N__22007));
    ClkMux I__5408 (
            .O(N__22214),
            .I(N__22007));
    ClkMux I__5407 (
            .O(N__22213),
            .I(N__22007));
    ClkMux I__5406 (
            .O(N__22212),
            .I(N__22007));
    ClkMux I__5405 (
            .O(N__22211),
            .I(N__22007));
    ClkMux I__5404 (
            .O(N__22210),
            .I(N__22007));
    ClkMux I__5403 (
            .O(N__22209),
            .I(N__22007));
    ClkMux I__5402 (
            .O(N__22208),
            .I(N__22007));
    ClkMux I__5401 (
            .O(N__22207),
            .I(N__22007));
    ClkMux I__5400 (
            .O(N__22206),
            .I(N__22007));
    ClkMux I__5399 (
            .O(N__22205),
            .I(N__22007));
    ClkMux I__5398 (
            .O(N__22204),
            .I(N__22007));
    ClkMux I__5397 (
            .O(N__22203),
            .I(N__22007));
    ClkMux I__5396 (
            .O(N__22202),
            .I(N__22007));
    ClkMux I__5395 (
            .O(N__22201),
            .I(N__22007));
    ClkMux I__5394 (
            .O(N__22200),
            .I(N__22007));
    ClkMux I__5393 (
            .O(N__22199),
            .I(N__22007));
    ClkMux I__5392 (
            .O(N__22198),
            .I(N__22007));
    ClkMux I__5391 (
            .O(N__22197),
            .I(N__22007));
    ClkMux I__5390 (
            .O(N__22196),
            .I(N__22007));
    ClkMux I__5389 (
            .O(N__22195),
            .I(N__22007));
    ClkMux I__5388 (
            .O(N__22194),
            .I(N__22007));
    ClkMux I__5387 (
            .O(N__22193),
            .I(N__22007));
    ClkMux I__5386 (
            .O(N__22192),
            .I(N__22007));
    ClkMux I__5385 (
            .O(N__22191),
            .I(N__22007));
    ClkMux I__5384 (
            .O(N__22190),
            .I(N__22007));
    ClkMux I__5383 (
            .O(N__22189),
            .I(N__22007));
    ClkMux I__5382 (
            .O(N__22188),
            .I(N__22007));
    ClkMux I__5381 (
            .O(N__22187),
            .I(N__22007));
    ClkMux I__5380 (
            .O(N__22186),
            .I(N__22007));
    ClkMux I__5379 (
            .O(N__22185),
            .I(N__22007));
    ClkMux I__5378 (
            .O(N__22184),
            .I(N__22007));
    ClkMux I__5377 (
            .O(N__22183),
            .I(N__22007));
    ClkMux I__5376 (
            .O(N__22182),
            .I(N__22007));
    ClkMux I__5375 (
            .O(N__22181),
            .I(N__22007));
    ClkMux I__5374 (
            .O(N__22180),
            .I(N__22007));
    ClkMux I__5373 (
            .O(N__22179),
            .I(N__22007));
    ClkMux I__5372 (
            .O(N__22178),
            .I(N__22007));
    ClkMux I__5371 (
            .O(N__22177),
            .I(N__22007));
    ClkMux I__5370 (
            .O(N__22176),
            .I(N__22007));
    ClkMux I__5369 (
            .O(N__22175),
            .I(N__22007));
    ClkMux I__5368 (
            .O(N__22174),
            .I(N__22007));
    ClkMux I__5367 (
            .O(N__22173),
            .I(N__22007));
    ClkMux I__5366 (
            .O(N__22172),
            .I(N__22007));
    ClkMux I__5365 (
            .O(N__22171),
            .I(N__22007));
    ClkMux I__5364 (
            .O(N__22170),
            .I(N__22007));
    ClkMux I__5363 (
            .O(N__22169),
            .I(N__22007));
    ClkMux I__5362 (
            .O(N__22168),
            .I(N__22007));
    ClkMux I__5361 (
            .O(N__22167),
            .I(N__22007));
    ClkMux I__5360 (
            .O(N__22166),
            .I(N__22007));
    GlobalMux I__5359 (
            .O(N__22007),
            .I(N__22004));
    gio2CtrlBuf I__5358 (
            .O(N__22004),
            .I(clk_0_c_g));
    InMux I__5357 (
            .O(N__22001),
            .I(N__21984));
    InMux I__5356 (
            .O(N__22000),
            .I(N__21981));
    InMux I__5355 (
            .O(N__21999),
            .I(N__21976));
    InMux I__5354 (
            .O(N__21998),
            .I(N__21976));
    InMux I__5353 (
            .O(N__21997),
            .I(N__21973));
    InMux I__5352 (
            .O(N__21996),
            .I(N__21970));
    InMux I__5351 (
            .O(N__21995),
            .I(N__21967));
    InMux I__5350 (
            .O(N__21994),
            .I(N__21964));
    InMux I__5349 (
            .O(N__21993),
            .I(N__21957));
    InMux I__5348 (
            .O(N__21992),
            .I(N__21957));
    InMux I__5347 (
            .O(N__21991),
            .I(N__21957));
    InMux I__5346 (
            .O(N__21990),
            .I(N__21954));
    InMux I__5345 (
            .O(N__21989),
            .I(N__21951));
    InMux I__5344 (
            .O(N__21988),
            .I(N__21946));
    InMux I__5343 (
            .O(N__21987),
            .I(N__21946));
    LocalMux I__5342 (
            .O(N__21984),
            .I(N__21934));
    LocalMux I__5341 (
            .O(N__21981),
            .I(N__21931));
    LocalMux I__5340 (
            .O(N__21976),
            .I(N__21928));
    LocalMux I__5339 (
            .O(N__21973),
            .I(N__21925));
    LocalMux I__5338 (
            .O(N__21970),
            .I(N__21922));
    LocalMux I__5337 (
            .O(N__21967),
            .I(N__21919));
    LocalMux I__5336 (
            .O(N__21964),
            .I(N__21916));
    LocalMux I__5335 (
            .O(N__21957),
            .I(N__21913));
    LocalMux I__5334 (
            .O(N__21954),
            .I(N__21910));
    LocalMux I__5333 (
            .O(N__21951),
            .I(N__21907));
    LocalMux I__5332 (
            .O(N__21946),
            .I(N__21904));
    SRMux I__5331 (
            .O(N__21945),
            .I(N__21863));
    SRMux I__5330 (
            .O(N__21944),
            .I(N__21863));
    SRMux I__5329 (
            .O(N__21943),
            .I(N__21863));
    SRMux I__5328 (
            .O(N__21942),
            .I(N__21863));
    SRMux I__5327 (
            .O(N__21941),
            .I(N__21863));
    SRMux I__5326 (
            .O(N__21940),
            .I(N__21863));
    SRMux I__5325 (
            .O(N__21939),
            .I(N__21863));
    SRMux I__5324 (
            .O(N__21938),
            .I(N__21863));
    SRMux I__5323 (
            .O(N__21937),
            .I(N__21863));
    Glb2LocalMux I__5322 (
            .O(N__21934),
            .I(N__21863));
    Glb2LocalMux I__5321 (
            .O(N__21931),
            .I(N__21863));
    Glb2LocalMux I__5320 (
            .O(N__21928),
            .I(N__21863));
    Glb2LocalMux I__5319 (
            .O(N__21925),
            .I(N__21863));
    Glb2LocalMux I__5318 (
            .O(N__21922),
            .I(N__21863));
    Glb2LocalMux I__5317 (
            .O(N__21919),
            .I(N__21863));
    Glb2LocalMux I__5316 (
            .O(N__21916),
            .I(N__21863));
    Glb2LocalMux I__5315 (
            .O(N__21913),
            .I(N__21863));
    Glb2LocalMux I__5314 (
            .O(N__21910),
            .I(N__21863));
    Glb2LocalMux I__5313 (
            .O(N__21907),
            .I(N__21863));
    Glb2LocalMux I__5312 (
            .O(N__21904),
            .I(N__21863));
    GlobalMux I__5311 (
            .O(N__21863),
            .I(N__21860));
    gio2CtrlBuf I__5310 (
            .O(N__21860),
            .I(M_this_state_q_nss_g_0));
    InMux I__5309 (
            .O(N__21857),
            .I(N__21854));
    LocalMux I__5308 (
            .O(N__21854),
            .I(N__21851));
    Span12Mux_v I__5307 (
            .O(N__21851),
            .I(N__21848));
    Odrv12 I__5306 (
            .O(N__21848),
            .I(port_address_in_3));
    InMux I__5305 (
            .O(N__21845),
            .I(N__21842));
    LocalMux I__5304 (
            .O(N__21842),
            .I(port_address_in_4));
    CascadeMux I__5303 (
            .O(N__21839),
            .I(N__21836));
    InMux I__5302 (
            .O(N__21836),
            .I(N__21833));
    LocalMux I__5301 (
            .O(N__21833),
            .I(port_address_in_5));
    InMux I__5300 (
            .O(N__21830),
            .I(N__21827));
    LocalMux I__5299 (
            .O(N__21827),
            .I(N__21824));
    Span4Mux_s3_h I__5298 (
            .O(N__21824),
            .I(N__21821));
    Span4Mux_v I__5297 (
            .O(N__21821),
            .I(N__21818));
    Span4Mux_v I__5296 (
            .O(N__21818),
            .I(N__21815));
    IoSpan4Mux I__5295 (
            .O(N__21815),
            .I(N__21812));
    IoSpan4Mux I__5294 (
            .O(N__21812),
            .I(N__21809));
    Odrv4 I__5293 (
            .O(N__21809),
            .I(port_address_in_2));
    InMux I__5292 (
            .O(N__21806),
            .I(N__21803));
    LocalMux I__5291 (
            .O(N__21803),
            .I(N__21800));
    Span4Mux_v I__5290 (
            .O(N__21800),
            .I(N__21797));
    Span4Mux_v I__5289 (
            .O(N__21797),
            .I(N__21794));
    Span4Mux_v I__5288 (
            .O(N__21794),
            .I(N__21791));
    Span4Mux_v I__5287 (
            .O(N__21791),
            .I(N__21788));
    Span4Mux_v I__5286 (
            .O(N__21788),
            .I(N__21785));
    Odrv4 I__5285 (
            .O(N__21785),
            .I(port_address_in_7));
    CascadeMux I__5284 (
            .O(N__21782),
            .I(M_this_state_d36_2_0_3_cascade_));
    InMux I__5283 (
            .O(N__21779),
            .I(N__21776));
    LocalMux I__5282 (
            .O(N__21776),
            .I(N__21773));
    Span12Mux_v I__5281 (
            .O(N__21773),
            .I(N__21770));
    Odrv12 I__5280 (
            .O(N__21770),
            .I(port_address_in_6));
    CascadeMux I__5279 (
            .O(N__21767),
            .I(N__21761));
    CascadeMux I__5278 (
            .O(N__21766),
            .I(N__21758));
    CascadeMux I__5277 (
            .O(N__21765),
            .I(N__21755));
    InMux I__5276 (
            .O(N__21764),
            .I(N__21752));
    InMux I__5275 (
            .O(N__21761),
            .I(N__21745));
    InMux I__5274 (
            .O(N__21758),
            .I(N__21745));
    InMux I__5273 (
            .O(N__21755),
            .I(N__21745));
    LocalMux I__5272 (
            .O(N__21752),
            .I(N__21740));
    LocalMux I__5271 (
            .O(N__21745),
            .I(N__21740));
    Span12Mux_h I__5270 (
            .O(N__21740),
            .I(N__21737));
    Odrv12 I__5269 (
            .O(N__21737),
            .I(M_this_state_d37_1));
    IoInMux I__5268 (
            .O(N__21734),
            .I(N__21731));
    LocalMux I__5267 (
            .O(N__21731),
            .I(N__21728));
    Span12Mux_s2_h I__5266 (
            .O(N__21728),
            .I(N__21724));
    InMux I__5265 (
            .O(N__21727),
            .I(N__21721));
    Odrv12 I__5264 (
            .O(N__21724),
            .I(M_this_external_address_qZ0Z_6));
    LocalMux I__5263 (
            .O(N__21721),
            .I(M_this_external_address_qZ0Z_6));
    InMux I__5262 (
            .O(N__21716),
            .I(un1_M_this_external_address_q_cry_5));
    IoInMux I__5261 (
            .O(N__21713),
            .I(N__21710));
    LocalMux I__5260 (
            .O(N__21710),
            .I(N__21707));
    Span4Mux_s2_h I__5259 (
            .O(N__21707),
            .I(N__21704));
    Sp12to4 I__5258 (
            .O(N__21704),
            .I(N__21701));
    Span12Mux_v I__5257 (
            .O(N__21701),
            .I(N__21697));
    InMux I__5256 (
            .O(N__21700),
            .I(N__21694));
    Odrv12 I__5255 (
            .O(N__21697),
            .I(M_this_external_address_qZ0Z_7));
    LocalMux I__5254 (
            .O(N__21694),
            .I(M_this_external_address_qZ0Z_7));
    InMux I__5253 (
            .O(N__21689),
            .I(un1_M_this_external_address_q_cry_6));
    IoInMux I__5252 (
            .O(N__21686),
            .I(N__21683));
    LocalMux I__5251 (
            .O(N__21683),
            .I(N__21680));
    IoSpan4Mux I__5250 (
            .O(N__21680),
            .I(N__21677));
    Span4Mux_s0_v I__5249 (
            .O(N__21677),
            .I(N__21674));
    Sp12to4 I__5248 (
            .O(N__21674),
            .I(N__21671));
    Span12Mux_v I__5247 (
            .O(N__21671),
            .I(N__21668));
    Span12Mux_h I__5246 (
            .O(N__21668),
            .I(N__21664));
    InMux I__5245 (
            .O(N__21667),
            .I(N__21661));
    Odrv12 I__5244 (
            .O(N__21664),
            .I(M_this_external_address_qZ0Z_8));
    LocalMux I__5243 (
            .O(N__21661),
            .I(M_this_external_address_qZ0Z_8));
    InMux I__5242 (
            .O(N__21656),
            .I(bfn_30_24_0_));
    IoInMux I__5241 (
            .O(N__21653),
            .I(N__21650));
    LocalMux I__5240 (
            .O(N__21650),
            .I(N__21647));
    Span12Mux_s8_v I__5239 (
            .O(N__21647),
            .I(N__21643));
    InMux I__5238 (
            .O(N__21646),
            .I(N__21640));
    Odrv12 I__5237 (
            .O(N__21643),
            .I(M_this_external_address_qZ0Z_9));
    LocalMux I__5236 (
            .O(N__21640),
            .I(M_this_external_address_qZ0Z_9));
    InMux I__5235 (
            .O(N__21635),
            .I(un1_M_this_external_address_q_cry_8));
    IoInMux I__5234 (
            .O(N__21632),
            .I(N__21629));
    LocalMux I__5233 (
            .O(N__21629),
            .I(N__21626));
    IoSpan4Mux I__5232 (
            .O(N__21626),
            .I(N__21623));
    Span4Mux_s2_v I__5231 (
            .O(N__21623),
            .I(N__21620));
    Sp12to4 I__5230 (
            .O(N__21620),
            .I(N__21617));
    Span12Mux_s8_v I__5229 (
            .O(N__21617),
            .I(N__21613));
    InMux I__5228 (
            .O(N__21616),
            .I(N__21610));
    Odrv12 I__5227 (
            .O(N__21613),
            .I(M_this_external_address_qZ0Z_10));
    LocalMux I__5226 (
            .O(N__21610),
            .I(M_this_external_address_qZ0Z_10));
    InMux I__5225 (
            .O(N__21605),
            .I(un1_M_this_external_address_q_cry_9));
    IoInMux I__5224 (
            .O(N__21602),
            .I(N__21599));
    LocalMux I__5223 (
            .O(N__21599),
            .I(N__21595));
    InMux I__5222 (
            .O(N__21598),
            .I(N__21592));
    Odrv12 I__5221 (
            .O(N__21595),
            .I(M_this_external_address_qZ0Z_11));
    LocalMux I__5220 (
            .O(N__21592),
            .I(M_this_external_address_qZ0Z_11));
    InMux I__5219 (
            .O(N__21587),
            .I(un1_M_this_external_address_q_cry_10));
    IoInMux I__5218 (
            .O(N__21584),
            .I(N__21581));
    LocalMux I__5217 (
            .O(N__21581),
            .I(N__21577));
    InMux I__5216 (
            .O(N__21580),
            .I(N__21574));
    Odrv4 I__5215 (
            .O(N__21577),
            .I(M_this_external_address_qZ0Z_12));
    LocalMux I__5214 (
            .O(N__21574),
            .I(M_this_external_address_qZ0Z_12));
    InMux I__5213 (
            .O(N__21569),
            .I(un1_M_this_external_address_q_cry_11));
    IoInMux I__5212 (
            .O(N__21566),
            .I(N__21563));
    LocalMux I__5211 (
            .O(N__21563),
            .I(N__21560));
    IoSpan4Mux I__5210 (
            .O(N__21560),
            .I(N__21557));
    Sp12to4 I__5209 (
            .O(N__21557),
            .I(N__21553));
    InMux I__5208 (
            .O(N__21556),
            .I(N__21550));
    Odrv12 I__5207 (
            .O(N__21553),
            .I(M_this_external_address_qZ0Z_13));
    LocalMux I__5206 (
            .O(N__21550),
            .I(M_this_external_address_qZ0Z_13));
    InMux I__5205 (
            .O(N__21545),
            .I(un1_M_this_external_address_q_cry_12));
    CascadeMux I__5204 (
            .O(N__21542),
            .I(N__21539));
    InMux I__5203 (
            .O(N__21539),
            .I(N__21535));
    CascadeMux I__5202 (
            .O(N__21538),
            .I(N__21532));
    LocalMux I__5201 (
            .O(N__21535),
            .I(N__21528));
    InMux I__5200 (
            .O(N__21532),
            .I(N__21525));
    InMux I__5199 (
            .O(N__21531),
            .I(N__21522));
    Span4Mux_h I__5198 (
            .O(N__21528),
            .I(N__21519));
    LocalMux I__5197 (
            .O(N__21525),
            .I(N__21516));
    LocalMux I__5196 (
            .O(N__21522),
            .I(N__21513));
    Span4Mux_v I__5195 (
            .O(N__21519),
            .I(N__21510));
    Span4Mux_h I__5194 (
            .O(N__21516),
            .I(N__21507));
    Span12Mux_h I__5193 (
            .O(N__21513),
            .I(N__21504));
    Span4Mux_v I__5192 (
            .O(N__21510),
            .I(N__21501));
    Span4Mux_v I__5191 (
            .O(N__21507),
            .I(N__21498));
    Odrv12 I__5190 (
            .O(N__21504),
            .I(port_data_c_1));
    Odrv4 I__5189 (
            .O(N__21501),
            .I(port_data_c_1));
    Odrv4 I__5188 (
            .O(N__21498),
            .I(port_data_c_1));
    InMux I__5187 (
            .O(N__21491),
            .I(N__21483));
    InMux I__5186 (
            .O(N__21490),
            .I(N__21483));
    InMux I__5185 (
            .O(N__21489),
            .I(N__21478));
    InMux I__5184 (
            .O(N__21488),
            .I(N__21478));
    LocalMux I__5183 (
            .O(N__21483),
            .I(un1_M_this_state_q_2_0));
    LocalMux I__5182 (
            .O(N__21478),
            .I(un1_M_this_state_q_2_0));
    CascadeMux I__5181 (
            .O(N__21473),
            .I(N__21469));
    CascadeMux I__5180 (
            .O(N__21472),
            .I(N__21466));
    InMux I__5179 (
            .O(N__21469),
            .I(N__21462));
    InMux I__5178 (
            .O(N__21466),
            .I(N__21459));
    CascadeMux I__5177 (
            .O(N__21465),
            .I(N__21456));
    LocalMux I__5176 (
            .O(N__21462),
            .I(N__21451));
    LocalMux I__5175 (
            .O(N__21459),
            .I(N__21451));
    InMux I__5174 (
            .O(N__21456),
            .I(N__21448));
    Span4Mux_v I__5173 (
            .O(N__21451),
            .I(N__21445));
    LocalMux I__5172 (
            .O(N__21448),
            .I(N__21442));
    Sp12to4 I__5171 (
            .O(N__21445),
            .I(N__21439));
    Span4Mux_v I__5170 (
            .O(N__21442),
            .I(N__21436));
    Span12Mux_h I__5169 (
            .O(N__21439),
            .I(N__21433));
    Span4Mux_h I__5168 (
            .O(N__21436),
            .I(N__21430));
    Odrv12 I__5167 (
            .O(N__21433),
            .I(port_data_c_5));
    Odrv4 I__5166 (
            .O(N__21430),
            .I(port_data_c_5));
    InMux I__5165 (
            .O(N__21425),
            .I(N__21418));
    InMux I__5164 (
            .O(N__21424),
            .I(N__21418));
    InMux I__5163 (
            .O(N__21423),
            .I(N__21415));
    LocalMux I__5162 (
            .O(N__21418),
            .I(M_this_sprites_ram_write_data_0_sqmuxa));
    LocalMux I__5161 (
            .O(N__21415),
            .I(M_this_sprites_ram_write_data_0_sqmuxa));
    InMux I__5160 (
            .O(N__21410),
            .I(N__21407));
    LocalMux I__5159 (
            .O(N__21407),
            .I(N__21403));
    InMux I__5158 (
            .O(N__21406),
            .I(N__21400));
    Span4Mux_s2_v I__5157 (
            .O(N__21403),
            .I(N__21394));
    LocalMux I__5156 (
            .O(N__21400),
            .I(N__21394));
    InMux I__5155 (
            .O(N__21399),
            .I(N__21391));
    Span4Mux_v I__5154 (
            .O(N__21394),
            .I(N__21384));
    LocalMux I__5153 (
            .O(N__21391),
            .I(N__21384));
    InMux I__5152 (
            .O(N__21390),
            .I(N__21381));
    InMux I__5151 (
            .O(N__21389),
            .I(N__21377));
    Span4Mux_v I__5150 (
            .O(N__21384),
            .I(N__21371));
    LocalMux I__5149 (
            .O(N__21381),
            .I(N__21371));
    InMux I__5148 (
            .O(N__21380),
            .I(N__21368));
    LocalMux I__5147 (
            .O(N__21377),
            .I(N__21364));
    InMux I__5146 (
            .O(N__21376),
            .I(N__21361));
    Span4Mux_v I__5145 (
            .O(N__21371),
            .I(N__21356));
    LocalMux I__5144 (
            .O(N__21368),
            .I(N__21356));
    InMux I__5143 (
            .O(N__21367),
            .I(N__21353));
    Span4Mux_v I__5142 (
            .O(N__21364),
            .I(N__21348));
    LocalMux I__5141 (
            .O(N__21361),
            .I(N__21348));
    Span4Mux_v I__5140 (
            .O(N__21356),
            .I(N__21343));
    LocalMux I__5139 (
            .O(N__21353),
            .I(N__21343));
    Odrv4 I__5138 (
            .O(N__21348),
            .I(M_this_sprites_ram_write_data_0_i_1));
    Odrv4 I__5137 (
            .O(N__21343),
            .I(M_this_sprites_ram_write_data_0_i_1));
    InMux I__5136 (
            .O(N__21338),
            .I(N__21335));
    LocalMux I__5135 (
            .O(N__21335),
            .I(N__21332));
    Span4Mux_v I__5134 (
            .O(N__21332),
            .I(N__21328));
    InMux I__5133 (
            .O(N__21331),
            .I(N__21321));
    Span4Mux_v I__5132 (
            .O(N__21328),
            .I(N__21317));
    InMux I__5131 (
            .O(N__21327),
            .I(N__21310));
    InMux I__5130 (
            .O(N__21326),
            .I(N__21310));
    InMux I__5129 (
            .O(N__21325),
            .I(N__21310));
    InMux I__5128 (
            .O(N__21324),
            .I(N__21307));
    LocalMux I__5127 (
            .O(N__21321),
            .I(N__21304));
    InMux I__5126 (
            .O(N__21320),
            .I(N__21301));
    Span4Mux_v I__5125 (
            .O(N__21317),
            .I(N__21297));
    LocalMux I__5124 (
            .O(N__21310),
            .I(N__21292));
    LocalMux I__5123 (
            .O(N__21307),
            .I(N__21292));
    Span4Mux_v I__5122 (
            .O(N__21304),
            .I(N__21289));
    LocalMux I__5121 (
            .O(N__21301),
            .I(N__21286));
    InMux I__5120 (
            .O(N__21300),
            .I(N__21283));
    Sp12to4 I__5119 (
            .O(N__21297),
            .I(N__21270));
    Span12Mux_v I__5118 (
            .O(N__21292),
            .I(N__21270));
    Sp12to4 I__5117 (
            .O(N__21289),
            .I(N__21270));
    Span12Mux_s8_h I__5116 (
            .O(N__21286),
            .I(N__21270));
    LocalMux I__5115 (
            .O(N__21283),
            .I(N__21270));
    InMux I__5114 (
            .O(N__21282),
            .I(N__21265));
    InMux I__5113 (
            .O(N__21281),
            .I(N__21265));
    Odrv12 I__5112 (
            .O(N__21270),
            .I(M_this_sprites_address_qZ0Z_12));
    LocalMux I__5111 (
            .O(N__21265),
            .I(M_this_sprites_address_qZ0Z_12));
    InMux I__5110 (
            .O(N__21260),
            .I(N__21250));
    InMux I__5109 (
            .O(N__21259),
            .I(N__21250));
    InMux I__5108 (
            .O(N__21258),
            .I(N__21250));
    InMux I__5107 (
            .O(N__21257),
            .I(N__21244));
    LocalMux I__5106 (
            .O(N__21250),
            .I(N__21241));
    InMux I__5105 (
            .O(N__21249),
            .I(N__21238));
    InMux I__5104 (
            .O(N__21248),
            .I(N__21235));
    InMux I__5103 (
            .O(N__21247),
            .I(N__21231));
    LocalMux I__5102 (
            .O(N__21244),
            .I(N__21228));
    Span4Mux_h I__5101 (
            .O(N__21241),
            .I(N__21225));
    LocalMux I__5100 (
            .O(N__21238),
            .I(N__21222));
    LocalMux I__5099 (
            .O(N__21235),
            .I(N__21219));
    InMux I__5098 (
            .O(N__21234),
            .I(N__21216));
    LocalMux I__5097 (
            .O(N__21231),
            .I(N__21213));
    Sp12to4 I__5096 (
            .O(N__21228),
            .I(N__21210));
    Span4Mux_v I__5095 (
            .O(N__21225),
            .I(N__21205));
    Span4Mux_h I__5094 (
            .O(N__21222),
            .I(N__21205));
    Span4Mux_v I__5093 (
            .O(N__21219),
            .I(N__21202));
    LocalMux I__5092 (
            .O(N__21216),
            .I(N__21199));
    Span4Mux_h I__5091 (
            .O(N__21213),
            .I(N__21196));
    Odrv12 I__5090 (
            .O(N__21210),
            .I(M_this_sprites_ram_write_en_1_0_0));
    Odrv4 I__5089 (
            .O(N__21205),
            .I(M_this_sprites_ram_write_en_1_0_0));
    Odrv4 I__5088 (
            .O(N__21202),
            .I(M_this_sprites_ram_write_en_1_0_0));
    Odrv4 I__5087 (
            .O(N__21199),
            .I(M_this_sprites_ram_write_en_1_0_0));
    Odrv4 I__5086 (
            .O(N__21196),
            .I(M_this_sprites_ram_write_en_1_0_0));
    CascadeMux I__5085 (
            .O(N__21185),
            .I(N__21179));
    CascadeMux I__5084 (
            .O(N__21184),
            .I(N__21176));
    CascadeMux I__5083 (
            .O(N__21183),
            .I(N__21172));
    InMux I__5082 (
            .O(N__21182),
            .I(N__21165));
    InMux I__5081 (
            .O(N__21179),
            .I(N__21165));
    InMux I__5080 (
            .O(N__21176),
            .I(N__21165));
    CascadeMux I__5079 (
            .O(N__21175),
            .I(N__21162));
    InMux I__5078 (
            .O(N__21172),
            .I(N__21157));
    LocalMux I__5077 (
            .O(N__21165),
            .I(N__21153));
    InMux I__5076 (
            .O(N__21162),
            .I(N__21150));
    CascadeMux I__5075 (
            .O(N__21161),
            .I(N__21147));
    CascadeMux I__5074 (
            .O(N__21160),
            .I(N__21144));
    LocalMux I__5073 (
            .O(N__21157),
            .I(N__21141));
    CascadeMux I__5072 (
            .O(N__21156),
            .I(N__21138));
    Span4Mux_v I__5071 (
            .O(N__21153),
            .I(N__21133));
    LocalMux I__5070 (
            .O(N__21150),
            .I(N__21133));
    InMux I__5069 (
            .O(N__21147),
            .I(N__21130));
    InMux I__5068 (
            .O(N__21144),
            .I(N__21127));
    Span4Mux_v I__5067 (
            .O(N__21141),
            .I(N__21124));
    InMux I__5066 (
            .O(N__21138),
            .I(N__21121));
    Span4Mux_v I__5065 (
            .O(N__21133),
            .I(N__21116));
    LocalMux I__5064 (
            .O(N__21130),
            .I(N__21116));
    LocalMux I__5063 (
            .O(N__21127),
            .I(N__21113));
    Span4Mux_v I__5062 (
            .O(N__21124),
            .I(N__21110));
    LocalMux I__5061 (
            .O(N__21121),
            .I(N__21107));
    Span4Mux_v I__5060 (
            .O(N__21116),
            .I(N__21101));
    Span4Mux_v I__5059 (
            .O(N__21113),
            .I(N__21101));
    Span4Mux_v I__5058 (
            .O(N__21110),
            .I(N__21096));
    Span4Mux_v I__5057 (
            .O(N__21107),
            .I(N__21096));
    InMux I__5056 (
            .O(N__21106),
            .I(N__21093));
    Sp12to4 I__5055 (
            .O(N__21101),
            .I(N__21085));
    Sp12to4 I__5054 (
            .O(N__21096),
            .I(N__21085));
    LocalMux I__5053 (
            .O(N__21093),
            .I(N__21085));
    InMux I__5052 (
            .O(N__21092),
            .I(N__21082));
    Odrv12 I__5051 (
            .O(N__21085),
            .I(M_this_sprites_address_qZ0Z_13));
    LocalMux I__5050 (
            .O(N__21082),
            .I(M_this_sprites_address_qZ0Z_13));
    CascadeMux I__5049 (
            .O(N__21077),
            .I(N__21073));
    InMux I__5048 (
            .O(N__21076),
            .I(N__21068));
    InMux I__5047 (
            .O(N__21073),
            .I(N__21061));
    InMux I__5046 (
            .O(N__21072),
            .I(N__21061));
    InMux I__5045 (
            .O(N__21071),
            .I(N__21061));
    LocalMux I__5044 (
            .O(N__21068),
            .I(N__21057));
    LocalMux I__5043 (
            .O(N__21061),
            .I(N__21054));
    InMux I__5042 (
            .O(N__21060),
            .I(N__21051));
    Span4Mux_v I__5041 (
            .O(N__21057),
            .I(N__21047));
    Span4Mux_v I__5040 (
            .O(N__21054),
            .I(N__21042));
    LocalMux I__5039 (
            .O(N__21051),
            .I(N__21042));
    InMux I__5038 (
            .O(N__21050),
            .I(N__21039));
    Span4Mux_v I__5037 (
            .O(N__21047),
            .I(N__21036));
    Span4Mux_v I__5036 (
            .O(N__21042),
            .I(N__21031));
    LocalMux I__5035 (
            .O(N__21039),
            .I(N__21031));
    Span4Mux_v I__5034 (
            .O(N__21036),
            .I(N__21026));
    Span4Mux_v I__5033 (
            .O(N__21031),
            .I(N__21023));
    InMux I__5032 (
            .O(N__21030),
            .I(N__21020));
    InMux I__5031 (
            .O(N__21029),
            .I(N__21017));
    Sp12to4 I__5030 (
            .O(N__21026),
            .I(N__21006));
    Sp12to4 I__5029 (
            .O(N__21023),
            .I(N__21006));
    LocalMux I__5028 (
            .O(N__21020),
            .I(N__21006));
    LocalMux I__5027 (
            .O(N__21017),
            .I(N__21006));
    InMux I__5026 (
            .O(N__21016),
            .I(N__21003));
    InMux I__5025 (
            .O(N__21015),
            .I(N__21000));
    Odrv12 I__5024 (
            .O(N__21006),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__5023 (
            .O(N__21003),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__5022 (
            .O(N__21000),
            .I(M_this_sprites_address_qZ0Z_11));
    CEMux I__5021 (
            .O(N__20993),
            .I(N__20990));
    LocalMux I__5020 (
            .O(N__20990),
            .I(N__20986));
    CEMux I__5019 (
            .O(N__20989),
            .I(N__20983));
    Span4Mux_v I__5018 (
            .O(N__20986),
            .I(N__20978));
    LocalMux I__5017 (
            .O(N__20983),
            .I(N__20978));
    Odrv4 I__5016 (
            .O(N__20978),
            .I(\this_sprites_ram.mem_WE_2 ));
    CascadeMux I__5015 (
            .O(N__20975),
            .I(N__20970));
    CascadeMux I__5014 (
            .O(N__20974),
            .I(N__20966));
    CascadeMux I__5013 (
            .O(N__20973),
            .I(N__20963));
    InMux I__5012 (
            .O(N__20970),
            .I(N__20955));
    InMux I__5011 (
            .O(N__20969),
            .I(N__20949));
    InMux I__5010 (
            .O(N__20966),
            .I(N__20946));
    InMux I__5009 (
            .O(N__20963),
            .I(N__20943));
    InMux I__5008 (
            .O(N__20962),
            .I(N__20938));
    InMux I__5007 (
            .O(N__20961),
            .I(N__20938));
    InMux I__5006 (
            .O(N__20960),
            .I(N__20931));
    InMux I__5005 (
            .O(N__20959),
            .I(N__20931));
    InMux I__5004 (
            .O(N__20958),
            .I(N__20931));
    LocalMux I__5003 (
            .O(N__20955),
            .I(N__20919));
    InMux I__5002 (
            .O(N__20954),
            .I(N__20916));
    InMux I__5001 (
            .O(N__20953),
            .I(N__20913));
    InMux I__5000 (
            .O(N__20952),
            .I(N__20910));
    LocalMux I__4999 (
            .O(N__20949),
            .I(N__20907));
    LocalMux I__4998 (
            .O(N__20946),
            .I(N__20904));
    LocalMux I__4997 (
            .O(N__20943),
            .I(N__20897));
    LocalMux I__4996 (
            .O(N__20938),
            .I(N__20897));
    LocalMux I__4995 (
            .O(N__20931),
            .I(N__20897));
    InMux I__4994 (
            .O(N__20930),
            .I(N__20888));
    InMux I__4993 (
            .O(N__20929),
            .I(N__20888));
    InMux I__4992 (
            .O(N__20928),
            .I(N__20888));
    InMux I__4991 (
            .O(N__20927),
            .I(N__20888));
    InMux I__4990 (
            .O(N__20926),
            .I(N__20879));
    InMux I__4989 (
            .O(N__20925),
            .I(N__20879));
    InMux I__4988 (
            .O(N__20924),
            .I(N__20879));
    InMux I__4987 (
            .O(N__20923),
            .I(N__20879));
    InMux I__4986 (
            .O(N__20922),
            .I(N__20876));
    Span4Mux_h I__4985 (
            .O(N__20919),
            .I(N__20873));
    LocalMux I__4984 (
            .O(N__20916),
            .I(N__20868));
    LocalMux I__4983 (
            .O(N__20913),
            .I(N__20868));
    LocalMux I__4982 (
            .O(N__20910),
            .I(N__20861));
    Sp12to4 I__4981 (
            .O(N__20907),
            .I(N__20861));
    Span12Mux_s2_h I__4980 (
            .O(N__20904),
            .I(N__20861));
    Span4Mux_v I__4979 (
            .O(N__20897),
            .I(N__20854));
    LocalMux I__4978 (
            .O(N__20888),
            .I(N__20854));
    LocalMux I__4977 (
            .O(N__20879),
            .I(N__20854));
    LocalMux I__4976 (
            .O(N__20876),
            .I(N__20851));
    Span4Mux_h I__4975 (
            .O(N__20873),
            .I(N__20846));
    Span4Mux_h I__4974 (
            .O(N__20868),
            .I(N__20846));
    Odrv12 I__4973 (
            .O(N__20861),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__4972 (
            .O(N__20854),
            .I(M_this_state_qZ0Z_3));
    Odrv12 I__4971 (
            .O(N__20851),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__4970 (
            .O(N__20846),
            .I(M_this_state_qZ0Z_3));
    IoInMux I__4969 (
            .O(N__20837),
            .I(N__20834));
    LocalMux I__4968 (
            .O(N__20834),
            .I(N__20831));
    Span4Mux_s1_v I__4967 (
            .O(N__20831),
            .I(N__20828));
    Sp12to4 I__4966 (
            .O(N__20828),
            .I(N__20825));
    Span12Mux_h I__4965 (
            .O(N__20825),
            .I(N__20821));
    InMux I__4964 (
            .O(N__20824),
            .I(N__20818));
    Odrv12 I__4963 (
            .O(N__20821),
            .I(M_this_external_address_qZ0Z_0));
    LocalMux I__4962 (
            .O(N__20818),
            .I(M_this_external_address_qZ0Z_0));
    IoInMux I__4961 (
            .O(N__20813),
            .I(N__20810));
    LocalMux I__4960 (
            .O(N__20810),
            .I(N__20807));
    IoSpan4Mux I__4959 (
            .O(N__20807),
            .I(N__20804));
    Sp12to4 I__4958 (
            .O(N__20804),
            .I(N__20800));
    InMux I__4957 (
            .O(N__20803),
            .I(N__20797));
    Odrv12 I__4956 (
            .O(N__20800),
            .I(M_this_external_address_qZ0Z_1));
    LocalMux I__4955 (
            .O(N__20797),
            .I(M_this_external_address_qZ0Z_1));
    InMux I__4954 (
            .O(N__20792),
            .I(un1_M_this_external_address_q_cry_0));
    IoInMux I__4953 (
            .O(N__20789),
            .I(N__20786));
    LocalMux I__4952 (
            .O(N__20786),
            .I(N__20783));
    IoSpan4Mux I__4951 (
            .O(N__20783),
            .I(N__20780));
    IoSpan4Mux I__4950 (
            .O(N__20780),
            .I(N__20777));
    Span4Mux_s2_v I__4949 (
            .O(N__20777),
            .I(N__20774));
    Span4Mux_v I__4948 (
            .O(N__20774),
            .I(N__20770));
    InMux I__4947 (
            .O(N__20773),
            .I(N__20767));
    Odrv4 I__4946 (
            .O(N__20770),
            .I(M_this_external_address_qZ0Z_2));
    LocalMux I__4945 (
            .O(N__20767),
            .I(M_this_external_address_qZ0Z_2));
    InMux I__4944 (
            .O(N__20762),
            .I(un1_M_this_external_address_q_cry_1));
    IoInMux I__4943 (
            .O(N__20759),
            .I(N__20756));
    LocalMux I__4942 (
            .O(N__20756),
            .I(N__20753));
    Span4Mux_s2_h I__4941 (
            .O(N__20753),
            .I(N__20750));
    Span4Mux_v I__4940 (
            .O(N__20750),
            .I(N__20746));
    InMux I__4939 (
            .O(N__20749),
            .I(N__20743));
    Odrv4 I__4938 (
            .O(N__20746),
            .I(M_this_external_address_qZ0Z_3));
    LocalMux I__4937 (
            .O(N__20743),
            .I(M_this_external_address_qZ0Z_3));
    InMux I__4936 (
            .O(N__20738),
            .I(un1_M_this_external_address_q_cry_2));
    IoInMux I__4935 (
            .O(N__20735),
            .I(N__20732));
    LocalMux I__4934 (
            .O(N__20732),
            .I(N__20728));
    InMux I__4933 (
            .O(N__20731),
            .I(N__20725));
    Odrv4 I__4932 (
            .O(N__20728),
            .I(M_this_external_address_qZ0Z_4));
    LocalMux I__4931 (
            .O(N__20725),
            .I(M_this_external_address_qZ0Z_4));
    InMux I__4930 (
            .O(N__20720),
            .I(un1_M_this_external_address_q_cry_3));
    IoInMux I__4929 (
            .O(N__20717),
            .I(N__20714));
    LocalMux I__4928 (
            .O(N__20714),
            .I(N__20711));
    Span4Mux_s2_h I__4927 (
            .O(N__20711),
            .I(N__20707));
    InMux I__4926 (
            .O(N__20710),
            .I(N__20704));
    Odrv4 I__4925 (
            .O(N__20707),
            .I(M_this_external_address_qZ0Z_5));
    LocalMux I__4924 (
            .O(N__20704),
            .I(M_this_external_address_qZ0Z_5));
    InMux I__4923 (
            .O(N__20699),
            .I(un1_M_this_external_address_q_cry_4));
    InMux I__4922 (
            .O(N__20696),
            .I(N__20693));
    LocalMux I__4921 (
            .O(N__20693),
            .I(N__20690));
    Sp12to4 I__4920 (
            .O(N__20690),
            .I(N__20687));
    Odrv12 I__4919 (
            .O(N__20687),
            .I(\this_sprites_ram.mem_out_bus5_2 ));
    CascadeMux I__4918 (
            .O(N__20684),
            .I(N__20679));
    CascadeMux I__4917 (
            .O(N__20683),
            .I(N__20675));
    InMux I__4916 (
            .O(N__20682),
            .I(N__20667));
    InMux I__4915 (
            .O(N__20679),
            .I(N__20667));
    CascadeMux I__4914 (
            .O(N__20678),
            .I(N__20664));
    InMux I__4913 (
            .O(N__20675),
            .I(N__20661));
    CascadeMux I__4912 (
            .O(N__20674),
            .I(N__20658));
    CascadeMux I__4911 (
            .O(N__20673),
            .I(N__20654));
    CascadeMux I__4910 (
            .O(N__20672),
            .I(N__20651));
    LocalMux I__4909 (
            .O(N__20667),
            .I(N__20648));
    InMux I__4908 (
            .O(N__20664),
            .I(N__20645));
    LocalMux I__4907 (
            .O(N__20661),
            .I(N__20642));
    InMux I__4906 (
            .O(N__20658),
            .I(N__20639));
    CascadeMux I__4905 (
            .O(N__20657),
            .I(N__20636));
    InMux I__4904 (
            .O(N__20654),
            .I(N__20633));
    InMux I__4903 (
            .O(N__20651),
            .I(N__20630));
    Span4Mux_v I__4902 (
            .O(N__20648),
            .I(N__20625));
    LocalMux I__4901 (
            .O(N__20645),
            .I(N__20625));
    Span4Mux_v I__4900 (
            .O(N__20642),
            .I(N__20620));
    LocalMux I__4899 (
            .O(N__20639),
            .I(N__20620));
    InMux I__4898 (
            .O(N__20636),
            .I(N__20617));
    LocalMux I__4897 (
            .O(N__20633),
            .I(N__20614));
    LocalMux I__4896 (
            .O(N__20630),
            .I(N__20611));
    Span4Mux_v I__4895 (
            .O(N__20625),
            .I(N__20608));
    Span4Mux_v I__4894 (
            .O(N__20620),
            .I(N__20605));
    LocalMux I__4893 (
            .O(N__20617),
            .I(N__20602));
    Span12Mux_s11_h I__4892 (
            .O(N__20614),
            .I(N__20597));
    Sp12to4 I__4891 (
            .O(N__20611),
            .I(N__20597));
    Odrv4 I__4890 (
            .O(N__20608),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__4889 (
            .O(N__20605),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__4888 (
            .O(N__20602),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv12 I__4887 (
            .O(N__20597),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    InMux I__4886 (
            .O(N__20588),
            .I(N__20585));
    LocalMux I__4885 (
            .O(N__20585),
            .I(N__20582));
    Span4Mux_v I__4884 (
            .O(N__20582),
            .I(N__20579));
    Odrv4 I__4883 (
            .O(N__20579),
            .I(\this_sprites_ram.mem_out_bus1_2 ));
    InMux I__4882 (
            .O(N__20576),
            .I(N__20573));
    LocalMux I__4881 (
            .O(N__20573),
            .I(N__20570));
    Sp12to4 I__4880 (
            .O(N__20570),
            .I(N__20567));
    Span12Mux_v I__4879 (
            .O(N__20567),
            .I(N__20564));
    Odrv12 I__4878 (
            .O(N__20564),
            .I(\this_sprites_ram.mem_out_bus7_2 ));
    InMux I__4877 (
            .O(N__20561),
            .I(N__20558));
    LocalMux I__4876 (
            .O(N__20558),
            .I(\this_sprites_ram.mem_out_bus3_2 ));
    CascadeMux I__4875 (
            .O(N__20555),
            .I(\this_sprites_ram.mem_DOUT_6_i_m2_ns_1_2_cascade_ ));
    InMux I__4874 (
            .O(N__20552),
            .I(N__20537));
    InMux I__4873 (
            .O(N__20551),
            .I(N__20537));
    InMux I__4872 (
            .O(N__20550),
            .I(N__20537));
    InMux I__4871 (
            .O(N__20549),
            .I(N__20537));
    InMux I__4870 (
            .O(N__20548),
            .I(N__20525));
    InMux I__4869 (
            .O(N__20547),
            .I(N__20525));
    InMux I__4868 (
            .O(N__20546),
            .I(N__20522));
    LocalMux I__4867 (
            .O(N__20537),
            .I(N__20519));
    InMux I__4866 (
            .O(N__20536),
            .I(N__20514));
    InMux I__4865 (
            .O(N__20535),
            .I(N__20514));
    InMux I__4864 (
            .O(N__20534),
            .I(N__20511));
    InMux I__4863 (
            .O(N__20533),
            .I(N__20506));
    InMux I__4862 (
            .O(N__20532),
            .I(N__20506));
    InMux I__4861 (
            .O(N__20531),
            .I(N__20503));
    InMux I__4860 (
            .O(N__20530),
            .I(N__20500));
    LocalMux I__4859 (
            .O(N__20525),
            .I(N__20497));
    LocalMux I__4858 (
            .O(N__20522),
            .I(N__20488));
    Span4Mux_h I__4857 (
            .O(N__20519),
            .I(N__20488));
    LocalMux I__4856 (
            .O(N__20514),
            .I(N__20488));
    LocalMux I__4855 (
            .O(N__20511),
            .I(N__20481));
    LocalMux I__4854 (
            .O(N__20506),
            .I(N__20481));
    LocalMux I__4853 (
            .O(N__20503),
            .I(N__20481));
    LocalMux I__4852 (
            .O(N__20500),
            .I(N__20476));
    Span4Mux_h I__4851 (
            .O(N__20497),
            .I(N__20476));
    InMux I__4850 (
            .O(N__20496),
            .I(N__20473));
    InMux I__4849 (
            .O(N__20495),
            .I(N__20470));
    Span4Mux_v I__4848 (
            .O(N__20488),
            .I(N__20467));
    Span4Mux_h I__4847 (
            .O(N__20481),
            .I(N__20464));
    Span4Mux_v I__4846 (
            .O(N__20476),
            .I(N__20459));
    LocalMux I__4845 (
            .O(N__20473),
            .I(N__20459));
    LocalMux I__4844 (
            .O(N__20470),
            .I(N__20456));
    Odrv4 I__4843 (
            .O(N__20467),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    Odrv4 I__4842 (
            .O(N__20464),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    Odrv4 I__4841 (
            .O(N__20459),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    Odrv12 I__4840 (
            .O(N__20456),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    InMux I__4839 (
            .O(N__20447),
            .I(N__20444));
    LocalMux I__4838 (
            .O(N__20444),
            .I(N__20441));
    Span4Mux_v I__4837 (
            .O(N__20441),
            .I(N__20438));
    Odrv4 I__4836 (
            .O(N__20438),
            .I(this_sprites_ram_mem_N_95));
    CEMux I__4835 (
            .O(N__20435),
            .I(N__20432));
    LocalMux I__4834 (
            .O(N__20432),
            .I(N__20428));
    CEMux I__4833 (
            .O(N__20431),
            .I(N__20425));
    Span4Mux_h I__4832 (
            .O(N__20428),
            .I(N__20422));
    LocalMux I__4831 (
            .O(N__20425),
            .I(N__20419));
    Odrv4 I__4830 (
            .O(N__20422),
            .I(\this_sprites_ram.mem_WE_6 ));
    Odrv12 I__4829 (
            .O(N__20419),
            .I(\this_sprites_ram.mem_WE_6 ));
    CEMux I__4828 (
            .O(N__20414),
            .I(N__20410));
    CEMux I__4827 (
            .O(N__20413),
            .I(N__20407));
    LocalMux I__4826 (
            .O(N__20410),
            .I(N__20404));
    LocalMux I__4825 (
            .O(N__20407),
            .I(N__20401));
    Span4Mux_h I__4824 (
            .O(N__20404),
            .I(N__20398));
    Span4Mux_h I__4823 (
            .O(N__20401),
            .I(N__20395));
    Odrv4 I__4822 (
            .O(N__20398),
            .I(\this_sprites_ram.mem_WE_4 ));
    Odrv4 I__4821 (
            .O(N__20395),
            .I(\this_sprites_ram.mem_WE_4 ));
    InMux I__4820 (
            .O(N__20390),
            .I(N__20384));
    InMux I__4819 (
            .O(N__20389),
            .I(N__20381));
    InMux I__4818 (
            .O(N__20388),
            .I(N__20378));
    InMux I__4817 (
            .O(N__20387),
            .I(N__20374));
    LocalMux I__4816 (
            .O(N__20384),
            .I(N__20370));
    LocalMux I__4815 (
            .O(N__20381),
            .I(N__20365));
    LocalMux I__4814 (
            .O(N__20378),
            .I(N__20365));
    InMux I__4813 (
            .O(N__20377),
            .I(N__20362));
    LocalMux I__4812 (
            .O(N__20374),
            .I(N__20359));
    InMux I__4811 (
            .O(N__20373),
            .I(N__20356));
    Span4Mux_h I__4810 (
            .O(N__20370),
            .I(N__20353));
    Span4Mux_h I__4809 (
            .O(N__20365),
            .I(N__20350));
    LocalMux I__4808 (
            .O(N__20362),
            .I(N__20343));
    Span12Mux_s8_h I__4807 (
            .O(N__20359),
            .I(N__20343));
    LocalMux I__4806 (
            .O(N__20356),
            .I(N__20343));
    Odrv4 I__4805 (
            .O(N__20353),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__4804 (
            .O(N__20350),
            .I(M_this_state_qZ0Z_2));
    Odrv12 I__4803 (
            .O(N__20343),
            .I(M_this_state_qZ0Z_2));
    CascadeMux I__4802 (
            .O(N__20336),
            .I(N__20332));
    InMux I__4801 (
            .O(N__20335),
            .I(N__20328));
    InMux I__4800 (
            .O(N__20332),
            .I(N__20318));
    InMux I__4799 (
            .O(N__20331),
            .I(N__20315));
    LocalMux I__4798 (
            .O(N__20328),
            .I(N__20312));
    InMux I__4797 (
            .O(N__20327),
            .I(N__20309));
    InMux I__4796 (
            .O(N__20326),
            .I(N__20306));
    InMux I__4795 (
            .O(N__20325),
            .I(N__20303));
    InMux I__4794 (
            .O(N__20324),
            .I(N__20298));
    InMux I__4793 (
            .O(N__20323),
            .I(N__20298));
    InMux I__4792 (
            .O(N__20322),
            .I(N__20295));
    InMux I__4791 (
            .O(N__20321),
            .I(N__20292));
    LocalMux I__4790 (
            .O(N__20318),
            .I(N__20283));
    LocalMux I__4789 (
            .O(N__20315),
            .I(N__20270));
    Span4Mux_v I__4788 (
            .O(N__20312),
            .I(N__20270));
    LocalMux I__4787 (
            .O(N__20309),
            .I(N__20270));
    LocalMux I__4786 (
            .O(N__20306),
            .I(N__20270));
    LocalMux I__4785 (
            .O(N__20303),
            .I(N__20270));
    LocalMux I__4784 (
            .O(N__20298),
            .I(N__20263));
    LocalMux I__4783 (
            .O(N__20295),
            .I(N__20263));
    LocalMux I__4782 (
            .O(N__20292),
            .I(N__20263));
    InMux I__4781 (
            .O(N__20291),
            .I(N__20259));
    InMux I__4780 (
            .O(N__20290),
            .I(N__20251));
    InMux I__4779 (
            .O(N__20289),
            .I(N__20244));
    InMux I__4778 (
            .O(N__20288),
            .I(N__20244));
    InMux I__4777 (
            .O(N__20287),
            .I(N__20244));
    InMux I__4776 (
            .O(N__20286),
            .I(N__20241));
    Span4Mux_v I__4775 (
            .O(N__20283),
            .I(N__20238));
    InMux I__4774 (
            .O(N__20282),
            .I(N__20235));
    InMux I__4773 (
            .O(N__20281),
            .I(N__20232));
    Span4Mux_v I__4772 (
            .O(N__20270),
            .I(N__20227));
    Span4Mux_v I__4771 (
            .O(N__20263),
            .I(N__20227));
    InMux I__4770 (
            .O(N__20262),
            .I(N__20224));
    LocalMux I__4769 (
            .O(N__20259),
            .I(N__20221));
    InMux I__4768 (
            .O(N__20258),
            .I(N__20216));
    InMux I__4767 (
            .O(N__20257),
            .I(N__20216));
    InMux I__4766 (
            .O(N__20256),
            .I(N__20213));
    InMux I__4765 (
            .O(N__20255),
            .I(N__20208));
    InMux I__4764 (
            .O(N__20254),
            .I(N__20208));
    LocalMux I__4763 (
            .O(N__20251),
            .I(N__20205));
    LocalMux I__4762 (
            .O(N__20244),
            .I(N__20202));
    LocalMux I__4761 (
            .O(N__20241),
            .I(N__20185));
    Sp12to4 I__4760 (
            .O(N__20238),
            .I(N__20185));
    LocalMux I__4759 (
            .O(N__20235),
            .I(N__20185));
    LocalMux I__4758 (
            .O(N__20232),
            .I(N__20185));
    Sp12to4 I__4757 (
            .O(N__20227),
            .I(N__20185));
    LocalMux I__4756 (
            .O(N__20224),
            .I(N__20185));
    Sp12to4 I__4755 (
            .O(N__20221),
            .I(N__20185));
    LocalMux I__4754 (
            .O(N__20216),
            .I(N__20185));
    LocalMux I__4753 (
            .O(N__20213),
            .I(M_this_start_data_delay_out_0));
    LocalMux I__4752 (
            .O(N__20208),
            .I(M_this_start_data_delay_out_0));
    Odrv4 I__4751 (
            .O(N__20205),
            .I(M_this_start_data_delay_out_0));
    Odrv4 I__4750 (
            .O(N__20202),
            .I(M_this_start_data_delay_out_0));
    Odrv12 I__4749 (
            .O(N__20185),
            .I(M_this_start_data_delay_out_0));
    CascadeMux I__4748 (
            .O(N__20174),
            .I(N__20170));
    InMux I__4747 (
            .O(N__20173),
            .I(N__20167));
    InMux I__4746 (
            .O(N__20170),
            .I(N__20164));
    LocalMux I__4745 (
            .O(N__20167),
            .I(N__20160));
    LocalMux I__4744 (
            .O(N__20164),
            .I(N__20157));
    CascadeMux I__4743 (
            .O(N__20163),
            .I(N__20154));
    Span4Mux_v I__4742 (
            .O(N__20160),
            .I(N__20151));
    Span4Mux_v I__4741 (
            .O(N__20157),
            .I(N__20148));
    InMux I__4740 (
            .O(N__20154),
            .I(N__20145));
    Sp12to4 I__4739 (
            .O(N__20151),
            .I(N__20142));
    Span4Mux_h I__4738 (
            .O(N__20148),
            .I(N__20137));
    LocalMux I__4737 (
            .O(N__20145),
            .I(N__20137));
    Span12Mux_h I__4736 (
            .O(N__20142),
            .I(N__20134));
    Span4Mux_h I__4735 (
            .O(N__20137),
            .I(N__20131));
    Span12Mux_v I__4734 (
            .O(N__20134),
            .I(N__20128));
    Sp12to4 I__4733 (
            .O(N__20131),
            .I(N__20125));
    Odrv12 I__4732 (
            .O(N__20128),
            .I(port_data_c_0));
    Odrv12 I__4731 (
            .O(N__20125),
            .I(port_data_c_0));
    CascadeMux I__4730 (
            .O(N__20120),
            .I(N__20115));
    CascadeMux I__4729 (
            .O(N__20119),
            .I(N__20112));
    InMux I__4728 (
            .O(N__20118),
            .I(N__20109));
    InMux I__4727 (
            .O(N__20115),
            .I(N__20106));
    InMux I__4726 (
            .O(N__20112),
            .I(N__20103));
    LocalMux I__4725 (
            .O(N__20109),
            .I(N__20100));
    LocalMux I__4724 (
            .O(N__20106),
            .I(N__20095));
    LocalMux I__4723 (
            .O(N__20103),
            .I(N__20095));
    Span4Mux_v I__4722 (
            .O(N__20100),
            .I(N__20092));
    Span12Mux_v I__4721 (
            .O(N__20095),
            .I(N__20089));
    Span4Mux_h I__4720 (
            .O(N__20092),
            .I(N__20086));
    Span12Mux_h I__4719 (
            .O(N__20089),
            .I(N__20083));
    IoSpan4Mux I__4718 (
            .O(N__20086),
            .I(N__20080));
    Odrv12 I__4717 (
            .O(N__20083),
            .I(port_data_c_4));
    Odrv4 I__4716 (
            .O(N__20080),
            .I(port_data_c_4));
    CascadeMux I__4715 (
            .O(N__20075),
            .I(M_this_sprites_ram_write_data_0_sqmuxa_cascade_));
    InMux I__4714 (
            .O(N__20072),
            .I(N__20069));
    LocalMux I__4713 (
            .O(N__20069),
            .I(N__20065));
    InMux I__4712 (
            .O(N__20068),
            .I(N__20062));
    Span4Mux_h I__4711 (
            .O(N__20065),
            .I(N__20058));
    LocalMux I__4710 (
            .O(N__20062),
            .I(N__20055));
    InMux I__4709 (
            .O(N__20061),
            .I(N__20052));
    Span4Mux_v I__4708 (
            .O(N__20058),
            .I(N__20045));
    Span4Mux_h I__4707 (
            .O(N__20055),
            .I(N__20045));
    LocalMux I__4706 (
            .O(N__20052),
            .I(N__20042));
    InMux I__4705 (
            .O(N__20051),
            .I(N__20039));
    InMux I__4704 (
            .O(N__20050),
            .I(N__20035));
    Span4Mux_v I__4703 (
            .O(N__20045),
            .I(N__20029));
    Span4Mux_h I__4702 (
            .O(N__20042),
            .I(N__20029));
    LocalMux I__4701 (
            .O(N__20039),
            .I(N__20026));
    InMux I__4700 (
            .O(N__20038),
            .I(N__20023));
    LocalMux I__4699 (
            .O(N__20035),
            .I(N__20020));
    InMux I__4698 (
            .O(N__20034),
            .I(N__20017));
    Span4Mux_v I__4697 (
            .O(N__20029),
            .I(N__20012));
    Span4Mux_h I__4696 (
            .O(N__20026),
            .I(N__20012));
    LocalMux I__4695 (
            .O(N__20023),
            .I(N__20009));
    Span4Mux_v I__4694 (
            .O(N__20020),
            .I(N__20004));
    LocalMux I__4693 (
            .O(N__20017),
            .I(N__20004));
    Span4Mux_v I__4692 (
            .O(N__20012),
            .I(N__19998));
    Span4Mux_h I__4691 (
            .O(N__20009),
            .I(N__19998));
    Span4Mux_v I__4690 (
            .O(N__20004),
            .I(N__19995));
    InMux I__4689 (
            .O(N__20003),
            .I(N__19992));
    Odrv4 I__4688 (
            .O(N__19998),
            .I(M_this_sprites_ram_write_data_0_i_0));
    Odrv4 I__4687 (
            .O(N__19995),
            .I(M_this_sprites_ram_write_data_0_i_0));
    LocalMux I__4686 (
            .O(N__19992),
            .I(M_this_sprites_ram_write_data_0_i_0));
    CascadeMux I__4685 (
            .O(N__19985),
            .I(N__19982));
    InMux I__4684 (
            .O(N__19982),
            .I(N__19979));
    LocalMux I__4683 (
            .O(N__19979),
            .I(N__19975));
    InMux I__4682 (
            .O(N__19978),
            .I(N__19972));
    Span4Mux_v I__4681 (
            .O(N__19975),
            .I(N__19968));
    LocalMux I__4680 (
            .O(N__19972),
            .I(N__19965));
    InMux I__4679 (
            .O(N__19971),
            .I(N__19962));
    Span4Mux_h I__4678 (
            .O(N__19968),
            .I(N__19957));
    Span4Mux_v I__4677 (
            .O(N__19965),
            .I(N__19957));
    LocalMux I__4676 (
            .O(N__19962),
            .I(N__19954));
    Span4Mux_v I__4675 (
            .O(N__19957),
            .I(N__19951));
    Span12Mux_h I__4674 (
            .O(N__19954),
            .I(N__19948));
    Span4Mux_h I__4673 (
            .O(N__19951),
            .I(N__19945));
    Odrv12 I__4672 (
            .O(N__19948),
            .I(port_data_c_3));
    Odrv4 I__4671 (
            .O(N__19945),
            .I(port_data_c_3));
    CascadeMux I__4670 (
            .O(N__19940),
            .I(N__19937));
    InMux I__4669 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__4668 (
            .O(N__19934),
            .I(N__19931));
    Span12Mux_h I__4667 (
            .O(N__19931),
            .I(N__19928));
    Span12Mux_v I__4666 (
            .O(N__19928),
            .I(N__19925));
    Odrv12 I__4665 (
            .O(N__19925),
            .I(port_data_c_7));
    InMux I__4664 (
            .O(N__19922),
            .I(N__19919));
    LocalMux I__4663 (
            .O(N__19919),
            .I(N__19915));
    InMux I__4662 (
            .O(N__19918),
            .I(N__19912));
    Span4Mux_v I__4661 (
            .O(N__19915),
            .I(N__19906));
    LocalMux I__4660 (
            .O(N__19912),
            .I(N__19906));
    InMux I__4659 (
            .O(N__19911),
            .I(N__19903));
    Span4Mux_v I__4658 (
            .O(N__19906),
            .I(N__19896));
    LocalMux I__4657 (
            .O(N__19903),
            .I(N__19896));
    InMux I__4656 (
            .O(N__19902),
            .I(N__19893));
    InMux I__4655 (
            .O(N__19901),
            .I(N__19890));
    Span4Mux_v I__4654 (
            .O(N__19896),
            .I(N__19883));
    LocalMux I__4653 (
            .O(N__19893),
            .I(N__19883));
    LocalMux I__4652 (
            .O(N__19890),
            .I(N__19880));
    InMux I__4651 (
            .O(N__19889),
            .I(N__19877));
    InMux I__4650 (
            .O(N__19888),
            .I(N__19874));
    Span4Mux_v I__4649 (
            .O(N__19883),
            .I(N__19871));
    Span4Mux_s3_v I__4648 (
            .O(N__19880),
            .I(N__19866));
    LocalMux I__4647 (
            .O(N__19877),
            .I(N__19866));
    LocalMux I__4646 (
            .O(N__19874),
            .I(N__19863));
    Span4Mux_v I__4645 (
            .O(N__19871),
            .I(N__19857));
    Span4Mux_v I__4644 (
            .O(N__19866),
            .I(N__19857));
    Span4Mux_h I__4643 (
            .O(N__19863),
            .I(N__19854));
    InMux I__4642 (
            .O(N__19862),
            .I(N__19851));
    Odrv4 I__4641 (
            .O(N__19857),
            .I(M_this_sprites_ram_write_data_0_i_3));
    Odrv4 I__4640 (
            .O(N__19854),
            .I(M_this_sprites_ram_write_data_0_i_3));
    LocalMux I__4639 (
            .O(N__19851),
            .I(M_this_sprites_ram_write_data_0_i_3));
    CascadeMux I__4638 (
            .O(N__19844),
            .I(N__19840));
    CascadeMux I__4637 (
            .O(N__19843),
            .I(N__19837));
    InMux I__4636 (
            .O(N__19840),
            .I(N__19834));
    InMux I__4635 (
            .O(N__19837),
            .I(N__19831));
    LocalMux I__4634 (
            .O(N__19834),
            .I(N__19828));
    LocalMux I__4633 (
            .O(N__19831),
            .I(N__19824));
    Span4Mux_v I__4632 (
            .O(N__19828),
            .I(N__19821));
    InMux I__4631 (
            .O(N__19827),
            .I(N__19818));
    Span4Mux_v I__4630 (
            .O(N__19824),
            .I(N__19815));
    Span4Mux_h I__4629 (
            .O(N__19821),
            .I(N__19810));
    LocalMux I__4628 (
            .O(N__19818),
            .I(N__19810));
    Sp12to4 I__4627 (
            .O(N__19815),
            .I(N__19807));
    Span4Mux_h I__4626 (
            .O(N__19810),
            .I(N__19804));
    Span12Mux_h I__4625 (
            .O(N__19807),
            .I(N__19799));
    Sp12to4 I__4624 (
            .O(N__19804),
            .I(N__19799));
    Odrv12 I__4623 (
            .O(N__19799),
            .I(port_data_c_2));
    CascadeMux I__4622 (
            .O(N__19796),
            .I(N__19792));
    CascadeMux I__4621 (
            .O(N__19795),
            .I(N__19789));
    InMux I__4620 (
            .O(N__19792),
            .I(N__19785));
    InMux I__4619 (
            .O(N__19789),
            .I(N__19782));
    CascadeMux I__4618 (
            .O(N__19788),
            .I(N__19779));
    LocalMux I__4617 (
            .O(N__19785),
            .I(N__19776));
    LocalMux I__4616 (
            .O(N__19782),
            .I(N__19773));
    InMux I__4615 (
            .O(N__19779),
            .I(N__19770));
    Span12Mux_v I__4614 (
            .O(N__19776),
            .I(N__19767));
    Span12Mux_h I__4613 (
            .O(N__19773),
            .I(N__19764));
    LocalMux I__4612 (
            .O(N__19770),
            .I(N__19761));
    Span12Mux_h I__4611 (
            .O(N__19767),
            .I(N__19756));
    Span12Mux_v I__4610 (
            .O(N__19764),
            .I(N__19756));
    Span12Mux_v I__4609 (
            .O(N__19761),
            .I(N__19753));
    Odrv12 I__4608 (
            .O(N__19756),
            .I(port_data_c_6));
    Odrv12 I__4607 (
            .O(N__19753),
            .I(port_data_c_6));
    InMux I__4606 (
            .O(N__19748),
            .I(N__19745));
    LocalMux I__4605 (
            .O(N__19745),
            .I(N__19740));
    InMux I__4604 (
            .O(N__19744),
            .I(N__19737));
    InMux I__4603 (
            .O(N__19743),
            .I(N__19733));
    Span4Mux_v I__4602 (
            .O(N__19740),
            .I(N__19727));
    LocalMux I__4601 (
            .O(N__19737),
            .I(N__19727));
    InMux I__4600 (
            .O(N__19736),
            .I(N__19724));
    LocalMux I__4599 (
            .O(N__19733),
            .I(N__19720));
    InMux I__4598 (
            .O(N__19732),
            .I(N__19717));
    Span4Mux_v I__4597 (
            .O(N__19727),
            .I(N__19712));
    LocalMux I__4596 (
            .O(N__19724),
            .I(N__19712));
    InMux I__4595 (
            .O(N__19723),
            .I(N__19709));
    Span4Mux_s3_v I__4594 (
            .O(N__19720),
            .I(N__19703));
    LocalMux I__4593 (
            .O(N__19717),
            .I(N__19703));
    Span4Mux_v I__4592 (
            .O(N__19712),
            .I(N__19698));
    LocalMux I__4591 (
            .O(N__19709),
            .I(N__19698));
    InMux I__4590 (
            .O(N__19708),
            .I(N__19695));
    Span4Mux_v I__4589 (
            .O(N__19703),
            .I(N__19691));
    Span4Mux_v I__4588 (
            .O(N__19698),
            .I(N__19686));
    LocalMux I__4587 (
            .O(N__19695),
            .I(N__19686));
    InMux I__4586 (
            .O(N__19694),
            .I(N__19683));
    Odrv4 I__4585 (
            .O(N__19691),
            .I(M_this_sprites_ram_write_data_0_i_2));
    Odrv4 I__4584 (
            .O(N__19686),
            .I(M_this_sprites_ram_write_data_0_i_2));
    LocalMux I__4583 (
            .O(N__19683),
            .I(M_this_sprites_ram_write_data_0_i_2));
    InMux I__4582 (
            .O(N__19676),
            .I(N__19673));
    LocalMux I__4581 (
            .O(N__19673),
            .I(N__19670));
    Span4Mux_v I__4580 (
            .O(N__19670),
            .I(N__19667));
    Span4Mux_v I__4579 (
            .O(N__19667),
            .I(N__19664));
    Odrv4 I__4578 (
            .O(N__19664),
            .I(\this_sprites_ram.mem_out_bus4_2 ));
    InMux I__4577 (
            .O(N__19661),
            .I(N__19658));
    LocalMux I__4576 (
            .O(N__19658),
            .I(N__19655));
    Span4Mux_v I__4575 (
            .O(N__19655),
            .I(N__19652));
    Odrv4 I__4574 (
            .O(N__19652),
            .I(\this_sprites_ram.mem_out_bus0_2 ));
    InMux I__4573 (
            .O(N__19649),
            .I(N__19646));
    LocalMux I__4572 (
            .O(N__19646),
            .I(N__19643));
    Span4Mux_h I__4571 (
            .O(N__19643),
            .I(N__19640));
    Sp12to4 I__4570 (
            .O(N__19640),
            .I(N__19637));
    Span12Mux_v I__4569 (
            .O(N__19637),
            .I(N__19634));
    Odrv12 I__4568 (
            .O(N__19634),
            .I(\this_sprites_ram.mem_out_bus6_2 ));
    InMux I__4567 (
            .O(N__19631),
            .I(N__19628));
    LocalMux I__4566 (
            .O(N__19628),
            .I(N__19625));
    Odrv4 I__4565 (
            .O(N__19625),
            .I(\this_sprites_ram.mem_out_bus2_2 ));
    CascadeMux I__4564 (
            .O(N__19622),
            .I(\this_sprites_ram.mem_DOUT_3_i_m2_ns_1_2_cascade_ ));
    InMux I__4563 (
            .O(N__19619),
            .I(N__19616));
    LocalMux I__4562 (
            .O(N__19616),
            .I(this_sprites_ram_mem_N_98));
    InMux I__4561 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__4560 (
            .O(N__19610),
            .I(N__19607));
    Span4Mux_v I__4559 (
            .O(N__19607),
            .I(N__19604));
    Span4Mux_v I__4558 (
            .O(N__19604),
            .I(N__19601));
    Odrv4 I__4557 (
            .O(N__19601),
            .I(\this_sprites_ram.mem_out_bus5_0 ));
    InMux I__4556 (
            .O(N__19598),
            .I(N__19595));
    LocalMux I__4555 (
            .O(N__19595),
            .I(N__19592));
    Span4Mux_v I__4554 (
            .O(N__19592),
            .I(N__19589));
    Odrv4 I__4553 (
            .O(N__19589),
            .I(\this_sprites_ram.mem_out_bus1_0 ));
    InMux I__4552 (
            .O(N__19586),
            .I(N__19583));
    LocalMux I__4551 (
            .O(N__19583),
            .I(N__19580));
    Odrv4 I__4550 (
            .O(N__19580),
            .I(\this_sprites_ram.mem_out_bus3_0 ));
    InMux I__4549 (
            .O(N__19577),
            .I(N__19574));
    LocalMux I__4548 (
            .O(N__19574),
            .I(N__19571));
    Span4Mux_v I__4547 (
            .O(N__19571),
            .I(N__19568));
    Sp12to4 I__4546 (
            .O(N__19568),
            .I(N__19565));
    Span12Mux_v I__4545 (
            .O(N__19565),
            .I(N__19562));
    Odrv12 I__4544 (
            .O(N__19562),
            .I(\this_sprites_ram.mem_out_bus7_0 ));
    CascadeMux I__4543 (
            .O(N__19559),
            .I(\this_sprites_ram.mem_DOUT_6_i_m2_ns_1_0_cascade_ ));
    InMux I__4542 (
            .O(N__19556),
            .I(N__19553));
    LocalMux I__4541 (
            .O(N__19553),
            .I(this_sprites_ram_mem_N_109));
    InMux I__4540 (
            .O(N__19550),
            .I(N__19547));
    LocalMux I__4539 (
            .O(N__19547),
            .I(N__19544));
    Span4Mux_v I__4538 (
            .O(N__19544),
            .I(N__19541));
    Span4Mux_v I__4537 (
            .O(N__19541),
            .I(N__19538));
    Odrv4 I__4536 (
            .O(N__19538),
            .I(\this_sprites_ram.mem_out_bus0_0 ));
    CascadeMux I__4535 (
            .O(N__19535),
            .I(N__19532));
    InMux I__4534 (
            .O(N__19532),
            .I(N__19529));
    LocalMux I__4533 (
            .O(N__19529),
            .I(N__19526));
    Span4Mux_v I__4532 (
            .O(N__19526),
            .I(N__19523));
    Span4Mux_h I__4531 (
            .O(N__19523),
            .I(N__19520));
    Odrv4 I__4530 (
            .O(N__19520),
            .I(\this_sprites_ram.mem_out_bus4_0 ));
    InMux I__4529 (
            .O(N__19517),
            .I(N__19514));
    LocalMux I__4528 (
            .O(N__19514),
            .I(N__19511));
    Sp12to4 I__4527 (
            .O(N__19511),
            .I(N__19508));
    Span12Mux_v I__4526 (
            .O(N__19508),
            .I(N__19505));
    Odrv12 I__4525 (
            .O(N__19505),
            .I(\this_sprites_ram.mem_out_bus6_0 ));
    CascadeMux I__4524 (
            .O(N__19502),
            .I(\this_sprites_ram.mem_DOUT_3_i_m2_ns_1_0_cascade_ ));
    InMux I__4523 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__4522 (
            .O(N__19496),
            .I(\this_sprites_ram.mem_out_bus2_0 ));
    InMux I__4521 (
            .O(N__19493),
            .I(N__19490));
    LocalMux I__4520 (
            .O(N__19490),
            .I(this_sprites_ram_mem_N_112));
    CEMux I__4519 (
            .O(N__19487),
            .I(N__19483));
    CEMux I__4518 (
            .O(N__19486),
            .I(N__19480));
    LocalMux I__4517 (
            .O(N__19483),
            .I(N__19477));
    LocalMux I__4516 (
            .O(N__19480),
            .I(N__19474));
    Span12Mux_s8_h I__4515 (
            .O(N__19477),
            .I(N__19471));
    Span4Mux_h I__4514 (
            .O(N__19474),
            .I(N__19468));
    Odrv12 I__4513 (
            .O(N__19471),
            .I(\this_sprites_ram.mem_WE_10 ));
    Odrv4 I__4512 (
            .O(N__19468),
            .I(\this_sprites_ram.mem_WE_10 ));
    CEMux I__4511 (
            .O(N__19463),
            .I(N__19460));
    LocalMux I__4510 (
            .O(N__19460),
            .I(N__19456));
    CEMux I__4509 (
            .O(N__19459),
            .I(N__19453));
    Span4Mux_v I__4508 (
            .O(N__19456),
            .I(N__19448));
    LocalMux I__4507 (
            .O(N__19453),
            .I(N__19448));
    Odrv4 I__4506 (
            .O(N__19448),
            .I(\this_sprites_ram.mem_WE_8 ));
    CEMux I__4505 (
            .O(N__19445),
            .I(N__19442));
    LocalMux I__4504 (
            .O(N__19442),
            .I(N__19438));
    CEMux I__4503 (
            .O(N__19441),
            .I(N__19435));
    Span4Mux_v I__4502 (
            .O(N__19438),
            .I(N__19430));
    LocalMux I__4501 (
            .O(N__19435),
            .I(N__19430));
    Span4Mux_v I__4500 (
            .O(N__19430),
            .I(N__19427));
    Span4Mux_h I__4499 (
            .O(N__19427),
            .I(N__19424));
    Odrv4 I__4498 (
            .O(N__19424),
            .I(\this_sprites_ram.mem_WE_12 ));
    CascadeMux I__4497 (
            .O(N__19421),
            .I(N__19418));
    InMux I__4496 (
            .O(N__19418),
            .I(N__19415));
    LocalMux I__4495 (
            .O(N__19415),
            .I(N__19412));
    Odrv12 I__4494 (
            .O(N__19412),
            .I(N_200));
    InMux I__4493 (
            .O(N__19409),
            .I(N__19406));
    LocalMux I__4492 (
            .O(N__19406),
            .I(N__19403));
    Span4Mux_v I__4491 (
            .O(N__19403),
            .I(N__19400));
    Sp12to4 I__4490 (
            .O(N__19400),
            .I(N__19397));
    Span12Mux_h I__4489 (
            .O(N__19397),
            .I(N__19394));
    Odrv12 I__4488 (
            .O(N__19394),
            .I(M_this_ppu_vram_data_2));
    InMux I__4487 (
            .O(N__19391),
            .I(N__19388));
    LocalMux I__4486 (
            .O(N__19388),
            .I(N__19382));
    InMux I__4485 (
            .O(N__19387),
            .I(N__19379));
    CEMux I__4484 (
            .O(N__19386),
            .I(N__19375));
    CascadeMux I__4483 (
            .O(N__19385),
            .I(N__19369));
    Span4Mux_v I__4482 (
            .O(N__19382),
            .I(N__19362));
    LocalMux I__4481 (
            .O(N__19379),
            .I(N__19362));
    InMux I__4480 (
            .O(N__19378),
            .I(N__19359));
    LocalMux I__4479 (
            .O(N__19375),
            .I(N__19356));
    InMux I__4478 (
            .O(N__19374),
            .I(N__19353));
    InMux I__4477 (
            .O(N__19373),
            .I(N__19350));
    InMux I__4476 (
            .O(N__19372),
            .I(N__19347));
    InMux I__4475 (
            .O(N__19369),
            .I(N__19344));
    InMux I__4474 (
            .O(N__19368),
            .I(N__19341));
    InMux I__4473 (
            .O(N__19367),
            .I(N__19338));
    Span4Mux_h I__4472 (
            .O(N__19362),
            .I(N__19333));
    LocalMux I__4471 (
            .O(N__19359),
            .I(N__19333));
    Sp12to4 I__4470 (
            .O(N__19356),
            .I(N__19330));
    LocalMux I__4469 (
            .O(N__19353),
            .I(N__19327));
    LocalMux I__4468 (
            .O(N__19350),
            .I(N__19322));
    LocalMux I__4467 (
            .O(N__19347),
            .I(N__19322));
    LocalMux I__4466 (
            .O(N__19344),
            .I(N__19319));
    LocalMux I__4465 (
            .O(N__19341),
            .I(N__19314));
    LocalMux I__4464 (
            .O(N__19338),
            .I(N__19314));
    Span4Mux_v I__4463 (
            .O(N__19333),
            .I(N__19311));
    Span12Mux_v I__4462 (
            .O(N__19330),
            .I(N__19306));
    Span12Mux_v I__4461 (
            .O(N__19327),
            .I(N__19306));
    Span4Mux_h I__4460 (
            .O(N__19322),
            .I(N__19303));
    Span4Mux_h I__4459 (
            .O(N__19319),
            .I(N__19298));
    Span4Mux_h I__4458 (
            .O(N__19314),
            .I(N__19298));
    Odrv4 I__4457 (
            .O(N__19311),
            .I(M_this_ppu_vram_en_0));
    Odrv12 I__4456 (
            .O(N__19306),
            .I(M_this_ppu_vram_en_0));
    Odrv4 I__4455 (
            .O(N__19303),
            .I(M_this_ppu_vram_en_0));
    Odrv4 I__4454 (
            .O(N__19298),
            .I(M_this_ppu_vram_en_0));
    CascadeMux I__4453 (
            .O(N__19289),
            .I(N__19286));
    InMux I__4452 (
            .O(N__19286),
            .I(N__19282));
    CascadeMux I__4451 (
            .O(N__19285),
            .I(N__19279));
    LocalMux I__4450 (
            .O(N__19282),
            .I(N__19275));
    InMux I__4449 (
            .O(N__19279),
            .I(N__19272));
    CascadeMux I__4448 (
            .O(N__19278),
            .I(N__19269));
    Span4Mux_h I__4447 (
            .O(N__19275),
            .I(N__19265));
    LocalMux I__4446 (
            .O(N__19272),
            .I(N__19262));
    InMux I__4445 (
            .O(N__19269),
            .I(N__19259));
    CascadeMux I__4444 (
            .O(N__19268),
            .I(N__19256));
    Span4Mux_v I__4443 (
            .O(N__19265),
            .I(N__19253));
    Span4Mux_h I__4442 (
            .O(N__19262),
            .I(N__19248));
    LocalMux I__4441 (
            .O(N__19259),
            .I(N__19248));
    InMux I__4440 (
            .O(N__19256),
            .I(N__19245));
    Span4Mux_v I__4439 (
            .O(N__19253),
            .I(N__19242));
    Span4Mux_v I__4438 (
            .O(N__19248),
            .I(N__19239));
    LocalMux I__4437 (
            .O(N__19245),
            .I(N__19236));
    Odrv4 I__4436 (
            .O(N__19242),
            .I(this_sprites_ram_mem_radreg_11));
    Odrv4 I__4435 (
            .O(N__19239),
            .I(this_sprites_ram_mem_radreg_11));
    Odrv12 I__4434 (
            .O(N__19236),
            .I(this_sprites_ram_mem_radreg_11));
    InMux I__4433 (
            .O(N__19229),
            .I(N__19226));
    LocalMux I__4432 (
            .O(N__19226),
            .I(N__19223));
    Span12Mux_h I__4431 (
            .O(N__19223),
            .I(N__19220));
    Odrv12 I__4430 (
            .O(N__19220),
            .I(M_this_ppu_vram_data_0));
    InMux I__4429 (
            .O(N__19217),
            .I(N__19214));
    LocalMux I__4428 (
            .O(N__19214),
            .I(N__19211));
    Span4Mux_h I__4427 (
            .O(N__19211),
            .I(N__19208));
    Odrv4 I__4426 (
            .O(N__19208),
            .I(\this_sprites_ram.mem_out_bus4_3 ));
    InMux I__4425 (
            .O(N__19205),
            .I(N__19202));
    LocalMux I__4424 (
            .O(N__19202),
            .I(N__19199));
    Span12Mux_h I__4423 (
            .O(N__19199),
            .I(N__19196));
    Span12Mux_v I__4422 (
            .O(N__19196),
            .I(N__19193));
    Odrv12 I__4421 (
            .O(N__19193),
            .I(\this_sprites_ram.mem_out_bus0_3 ));
    InMux I__4420 (
            .O(N__19190),
            .I(N__19187));
    LocalMux I__4419 (
            .O(N__19187),
            .I(\this_sprites_ram.mem_DOUT_3_i_m2_ns_1_3 ));
    InMux I__4418 (
            .O(N__19184),
            .I(N__19179));
    InMux I__4417 (
            .O(N__19183),
            .I(N__19174));
    InMux I__4416 (
            .O(N__19182),
            .I(N__19174));
    LocalMux I__4415 (
            .O(N__19179),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__4414 (
            .O(N__19174),
            .I(M_this_state_qZ0Z_7));
    InMux I__4413 (
            .O(N__19169),
            .I(N__19166));
    LocalMux I__4412 (
            .O(N__19166),
            .I(N__19162));
    InMux I__4411 (
            .O(N__19165),
            .I(N__19159));
    Span4Mux_h I__4410 (
            .O(N__19162),
            .I(N__19156));
    LocalMux I__4409 (
            .O(N__19159),
            .I(N_170_0));
    Odrv4 I__4408 (
            .O(N__19156),
            .I(N_170_0));
    CEMux I__4407 (
            .O(N__19151),
            .I(N__19148));
    LocalMux I__4406 (
            .O(N__19148),
            .I(N__19144));
    CEMux I__4405 (
            .O(N__19147),
            .I(N__19141));
    Span4Mux_h I__4404 (
            .O(N__19144),
            .I(N__19136));
    LocalMux I__4403 (
            .O(N__19141),
            .I(N__19136));
    Span4Mux_v I__4402 (
            .O(N__19136),
            .I(N__19133));
    Span4Mux_v I__4401 (
            .O(N__19133),
            .I(N__19130));
    Odrv4 I__4400 (
            .O(N__19130),
            .I(\this_sprites_ram.mem_WE_0 ));
    InMux I__4399 (
            .O(N__19127),
            .I(N__19121));
    InMux I__4398 (
            .O(N__19126),
            .I(N__19118));
    InMux I__4397 (
            .O(N__19125),
            .I(N__19115));
    InMux I__4396 (
            .O(N__19124),
            .I(N__19112));
    LocalMux I__4395 (
            .O(N__19121),
            .I(N__19105));
    LocalMux I__4394 (
            .O(N__19118),
            .I(N__19105));
    LocalMux I__4393 (
            .O(N__19115),
            .I(N__19105));
    LocalMux I__4392 (
            .O(N__19112),
            .I(\this_ppu.M_vaddress_qZ0Z_3 ));
    Odrv4 I__4391 (
            .O(N__19105),
            .I(\this_ppu.M_vaddress_qZ0Z_3 ));
    CascadeMux I__4390 (
            .O(N__19100),
            .I(N__19097));
    CascadeBuf I__4389 (
            .O(N__19097),
            .I(N__19094));
    CascadeMux I__4388 (
            .O(N__19094),
            .I(N__19091));
    CascadeBuf I__4387 (
            .O(N__19091),
            .I(N__19088));
    CascadeMux I__4386 (
            .O(N__19088),
            .I(N__19085));
    CascadeBuf I__4385 (
            .O(N__19085),
            .I(N__19082));
    CascadeMux I__4384 (
            .O(N__19082),
            .I(N__19079));
    CascadeBuf I__4383 (
            .O(N__19079),
            .I(N__19076));
    CascadeMux I__4382 (
            .O(N__19076),
            .I(N__19073));
    CascadeBuf I__4381 (
            .O(N__19073),
            .I(N__19070));
    CascadeMux I__4380 (
            .O(N__19070),
            .I(N__19067));
    CascadeBuf I__4379 (
            .O(N__19067),
            .I(N__19064));
    CascadeMux I__4378 (
            .O(N__19064),
            .I(N__19061));
    CascadeBuf I__4377 (
            .O(N__19061),
            .I(N__19058));
    CascadeMux I__4376 (
            .O(N__19058),
            .I(N__19055));
    CascadeBuf I__4375 (
            .O(N__19055),
            .I(N__19052));
    CascadeMux I__4374 (
            .O(N__19052),
            .I(N__19049));
    CascadeBuf I__4373 (
            .O(N__19049),
            .I(N__19046));
    CascadeMux I__4372 (
            .O(N__19046),
            .I(N__19043));
    CascadeBuf I__4371 (
            .O(N__19043),
            .I(N__19040));
    CascadeMux I__4370 (
            .O(N__19040),
            .I(N__19037));
    CascadeBuf I__4369 (
            .O(N__19037),
            .I(N__19034));
    CascadeMux I__4368 (
            .O(N__19034),
            .I(N__19031));
    CascadeBuf I__4367 (
            .O(N__19031),
            .I(N__19028));
    CascadeMux I__4366 (
            .O(N__19028),
            .I(N__19025));
    CascadeBuf I__4365 (
            .O(N__19025),
            .I(N__19022));
    CascadeMux I__4364 (
            .O(N__19022),
            .I(N__19019));
    CascadeBuf I__4363 (
            .O(N__19019),
            .I(N__19016));
    CascadeMux I__4362 (
            .O(N__19016),
            .I(N__19013));
    CascadeBuf I__4361 (
            .O(N__19013),
            .I(N__19010));
    CascadeMux I__4360 (
            .O(N__19010),
            .I(N__19007));
    InMux I__4359 (
            .O(N__19007),
            .I(N__19004));
    LocalMux I__4358 (
            .O(N__19004),
            .I(N__19001));
    Span12Mux_s11_h I__4357 (
            .O(N__19001),
            .I(N__18998));
    Span12Mux_v I__4356 (
            .O(N__18998),
            .I(N__18995));
    Odrv12 I__4355 (
            .O(N__18995),
            .I(M_this_ppu_sprites_addr_10));
    InMux I__4354 (
            .O(N__18992),
            .I(\this_ppu.sprites_addr_cry_9 ));
    CascadeMux I__4353 (
            .O(N__18989),
            .I(N__18985));
    InMux I__4352 (
            .O(N__18988),
            .I(N__18982));
    InMux I__4351 (
            .O(N__18985),
            .I(N__18978));
    LocalMux I__4350 (
            .O(N__18982),
            .I(N__18975));
    InMux I__4349 (
            .O(N__18981),
            .I(N__18972));
    LocalMux I__4348 (
            .O(N__18978),
            .I(\this_ppu.M_vaddress_qZ1Z_4 ));
    Odrv4 I__4347 (
            .O(N__18975),
            .I(\this_ppu.M_vaddress_qZ1Z_4 ));
    LocalMux I__4346 (
            .O(N__18972),
            .I(\this_ppu.M_vaddress_qZ1Z_4 ));
    InMux I__4345 (
            .O(N__18965),
            .I(\this_ppu.sprites_addr_cry_10 ));
    InMux I__4344 (
            .O(N__18962),
            .I(N__18955));
    InMux I__4343 (
            .O(N__18961),
            .I(N__18955));
    InMux I__4342 (
            .O(N__18960),
            .I(N__18952));
    LocalMux I__4341 (
            .O(N__18955),
            .I(N__18947));
    LocalMux I__4340 (
            .O(N__18952),
            .I(N__18947));
    Odrv4 I__4339 (
            .O(N__18947),
            .I(\this_ppu.M_vaddress_qZ0Z_5 ));
    InMux I__4338 (
            .O(N__18944),
            .I(\this_ppu.sprites_addr_cry_11 ));
    CascadeMux I__4337 (
            .O(N__18941),
            .I(N__18938));
    InMux I__4336 (
            .O(N__18938),
            .I(N__18934));
    InMux I__4335 (
            .O(N__18937),
            .I(N__18931));
    LocalMux I__4334 (
            .O(N__18934),
            .I(N__18926));
    LocalMux I__4333 (
            .O(N__18931),
            .I(N__18926));
    Odrv4 I__4332 (
            .O(N__18926),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    InMux I__4331 (
            .O(N__18923),
            .I(\this_ppu.sprites_addr_cry_12 ));
    CascadeMux I__4330 (
            .O(N__18920),
            .I(N__18917));
    InMux I__4329 (
            .O(N__18917),
            .I(N__18914));
    LocalMux I__4328 (
            .O(N__18914),
            .I(N__18911));
    Span4Mux_h I__4327 (
            .O(N__18911),
            .I(N__18907));
    InMux I__4326 (
            .O(N__18910),
            .I(N__18904));
    Sp12to4 I__4325 (
            .O(N__18907),
            .I(N__18897));
    LocalMux I__4324 (
            .O(N__18904),
            .I(N__18891));
    InMux I__4323 (
            .O(N__18903),
            .I(N__18888));
    InMux I__4322 (
            .O(N__18902),
            .I(N__18885));
    InMux I__4321 (
            .O(N__18901),
            .I(N__18880));
    InMux I__4320 (
            .O(N__18900),
            .I(N__18880));
    Span12Mux_v I__4319 (
            .O(N__18897),
            .I(N__18877));
    InMux I__4318 (
            .O(N__18896),
            .I(N__18872));
    InMux I__4317 (
            .O(N__18895),
            .I(N__18872));
    InMux I__4316 (
            .O(N__18894),
            .I(N__18869));
    Span4Mux_v I__4315 (
            .O(N__18891),
            .I(N__18862));
    LocalMux I__4314 (
            .O(N__18888),
            .I(N__18862));
    LocalMux I__4313 (
            .O(N__18885),
            .I(N__18862));
    LocalMux I__4312 (
            .O(N__18880),
            .I(N__18859));
    Odrv12 I__4311 (
            .O(N__18877),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__4310 (
            .O(N__18872),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__4309 (
            .O(N__18869),
            .I(M_this_ppu_vram_addr_0));
    Odrv4 I__4308 (
            .O(N__18862),
            .I(M_this_ppu_vram_addr_0));
    Odrv4 I__4307 (
            .O(N__18859),
            .I(M_this_ppu_vram_addr_0));
    CascadeMux I__4306 (
            .O(N__18848),
            .I(N__18845));
    CascadeBuf I__4305 (
            .O(N__18845),
            .I(N__18842));
    CascadeMux I__4304 (
            .O(N__18842),
            .I(N__18839));
    CascadeBuf I__4303 (
            .O(N__18839),
            .I(N__18836));
    CascadeMux I__4302 (
            .O(N__18836),
            .I(N__18833));
    CascadeBuf I__4301 (
            .O(N__18833),
            .I(N__18830));
    CascadeMux I__4300 (
            .O(N__18830),
            .I(N__18827));
    CascadeBuf I__4299 (
            .O(N__18827),
            .I(N__18824));
    CascadeMux I__4298 (
            .O(N__18824),
            .I(N__18821));
    CascadeBuf I__4297 (
            .O(N__18821),
            .I(N__18818));
    CascadeMux I__4296 (
            .O(N__18818),
            .I(N__18815));
    CascadeBuf I__4295 (
            .O(N__18815),
            .I(N__18812));
    CascadeMux I__4294 (
            .O(N__18812),
            .I(N__18809));
    CascadeBuf I__4293 (
            .O(N__18809),
            .I(N__18806));
    CascadeMux I__4292 (
            .O(N__18806),
            .I(N__18803));
    CascadeBuf I__4291 (
            .O(N__18803),
            .I(N__18800));
    CascadeMux I__4290 (
            .O(N__18800),
            .I(N__18797));
    CascadeBuf I__4289 (
            .O(N__18797),
            .I(N__18794));
    CascadeMux I__4288 (
            .O(N__18794),
            .I(N__18791));
    CascadeBuf I__4287 (
            .O(N__18791),
            .I(N__18788));
    CascadeMux I__4286 (
            .O(N__18788),
            .I(N__18785));
    CascadeBuf I__4285 (
            .O(N__18785),
            .I(N__18782));
    CascadeMux I__4284 (
            .O(N__18782),
            .I(N__18779));
    CascadeBuf I__4283 (
            .O(N__18779),
            .I(N__18776));
    CascadeMux I__4282 (
            .O(N__18776),
            .I(N__18773));
    CascadeBuf I__4281 (
            .O(N__18773),
            .I(N__18770));
    CascadeMux I__4280 (
            .O(N__18770),
            .I(N__18767));
    CascadeBuf I__4279 (
            .O(N__18767),
            .I(N__18764));
    CascadeMux I__4278 (
            .O(N__18764),
            .I(N__18761));
    CascadeBuf I__4277 (
            .O(N__18761),
            .I(N__18758));
    CascadeMux I__4276 (
            .O(N__18758),
            .I(N__18755));
    InMux I__4275 (
            .O(N__18755),
            .I(N__18752));
    LocalMux I__4274 (
            .O(N__18752),
            .I(N__18749));
    Span12Mux_v I__4273 (
            .O(N__18749),
            .I(N__18746));
    Odrv12 I__4272 (
            .O(N__18746),
            .I(M_this_ppu_vram_addr_i_0));
    InMux I__4271 (
            .O(N__18743),
            .I(N__18740));
    LocalMux I__4270 (
            .O(N__18740),
            .I(N__18737));
    Span12Mux_h I__4269 (
            .O(N__18737),
            .I(N__18734));
    Odrv12 I__4268 (
            .O(N__18734),
            .I(\this_sprites_ram.mem_out_bus5_1 ));
    InMux I__4267 (
            .O(N__18731),
            .I(N__18728));
    LocalMux I__4266 (
            .O(N__18728),
            .I(N__18725));
    Span4Mux_v I__4265 (
            .O(N__18725),
            .I(N__18722));
    Span4Mux_v I__4264 (
            .O(N__18722),
            .I(N__18719));
    Odrv4 I__4263 (
            .O(N__18719),
            .I(\this_sprites_ram.mem_out_bus1_1 ));
    InMux I__4262 (
            .O(N__18716),
            .I(N__18713));
    LocalMux I__4261 (
            .O(N__18713),
            .I(N__18710));
    Span4Mux_h I__4260 (
            .O(N__18710),
            .I(N__18707));
    Span4Mux_v I__4259 (
            .O(N__18707),
            .I(N__18704));
    Span4Mux_v I__4258 (
            .O(N__18704),
            .I(N__18701));
    Span4Mux_v I__4257 (
            .O(N__18701),
            .I(N__18698));
    Odrv4 I__4256 (
            .O(N__18698),
            .I(\this_sprites_ram.mem_out_bus7_1 ));
    InMux I__4255 (
            .O(N__18695),
            .I(N__18692));
    LocalMux I__4254 (
            .O(N__18692),
            .I(N__18689));
    Odrv4 I__4253 (
            .O(N__18689),
            .I(\this_sprites_ram.mem_out_bus3_1 ));
    CascadeMux I__4252 (
            .O(N__18686),
            .I(\this_sprites_ram.mem_DOUT_6_i_m2_ns_1_1_cascade_ ));
    InMux I__4251 (
            .O(N__18683),
            .I(N__18680));
    LocalMux I__4250 (
            .O(N__18680),
            .I(this_sprites_ram_mem_N_88));
    CEMux I__4249 (
            .O(N__18677),
            .I(N__18674));
    LocalMux I__4248 (
            .O(N__18674),
            .I(N__18671));
    Span4Mux_s3_v I__4247 (
            .O(N__18671),
            .I(N__18667));
    CEMux I__4246 (
            .O(N__18670),
            .I(N__18664));
    Span4Mux_h I__4245 (
            .O(N__18667),
            .I(N__18659));
    LocalMux I__4244 (
            .O(N__18664),
            .I(N__18659));
    Span4Mux_h I__4243 (
            .O(N__18659),
            .I(N__18656));
    Span4Mux_v I__4242 (
            .O(N__18656),
            .I(N__18653));
    Span4Mux_v I__4241 (
            .O(N__18653),
            .I(N__18650));
    Odrv4 I__4240 (
            .O(N__18650),
            .I(\this_sprites_ram.mem_WE_14 ));
    InMux I__4239 (
            .O(N__18647),
            .I(N__18644));
    LocalMux I__4238 (
            .O(N__18644),
            .I(N__18641));
    Span4Mux_v I__4237 (
            .O(N__18641),
            .I(N__18638));
    Odrv4 I__4236 (
            .O(N__18638),
            .I(\this_sprites_ram.mem_out_bus2_3 ));
    CascadeMux I__4235 (
            .O(N__18635),
            .I(N__18632));
    InMux I__4234 (
            .O(N__18632),
            .I(N__18629));
    LocalMux I__4233 (
            .O(N__18629),
            .I(N__18626));
    Span12Mux_h I__4232 (
            .O(N__18626),
            .I(N__18623));
    Span12Mux_v I__4231 (
            .O(N__18623),
            .I(N__18620));
    Odrv12 I__4230 (
            .O(N__18620),
            .I(\this_sprites_ram.mem_out_bus6_3 ));
    InMux I__4229 (
            .O(N__18617),
            .I(N__18614));
    LocalMux I__4228 (
            .O(N__18614),
            .I(N__18611));
    Span4Mux_h I__4227 (
            .O(N__18611),
            .I(N__18608));
    Odrv4 I__4226 (
            .O(N__18608),
            .I(this_sprites_ram_mem_N_105));
    InMux I__4225 (
            .O(N__18605),
            .I(\this_ppu.sprites_addr_cry_1 ));
    CascadeMux I__4224 (
            .O(N__18602),
            .I(N__18599));
    InMux I__4223 (
            .O(N__18599),
            .I(N__18596));
    LocalMux I__4222 (
            .O(N__18596),
            .I(N__18592));
    InMux I__4221 (
            .O(N__18595),
            .I(N__18587));
    Span12Mux_v I__4220 (
            .O(N__18592),
            .I(N__18582));
    InMux I__4219 (
            .O(N__18591),
            .I(N__18579));
    InMux I__4218 (
            .O(N__18590),
            .I(N__18576));
    LocalMux I__4217 (
            .O(N__18587),
            .I(N__18573));
    InMux I__4216 (
            .O(N__18586),
            .I(N__18568));
    InMux I__4215 (
            .O(N__18585),
            .I(N__18568));
    Odrv12 I__4214 (
            .O(N__18582),
            .I(M_this_ppu_vram_addr_3));
    LocalMux I__4213 (
            .O(N__18579),
            .I(M_this_ppu_vram_addr_3));
    LocalMux I__4212 (
            .O(N__18576),
            .I(M_this_ppu_vram_addr_3));
    Odrv12 I__4211 (
            .O(N__18573),
            .I(M_this_ppu_vram_addr_3));
    LocalMux I__4210 (
            .O(N__18568),
            .I(M_this_ppu_vram_addr_3));
    CascadeMux I__4209 (
            .O(N__18557),
            .I(N__18554));
    CascadeBuf I__4208 (
            .O(N__18554),
            .I(N__18551));
    CascadeMux I__4207 (
            .O(N__18551),
            .I(N__18548));
    CascadeBuf I__4206 (
            .O(N__18548),
            .I(N__18545));
    CascadeMux I__4205 (
            .O(N__18545),
            .I(N__18542));
    CascadeBuf I__4204 (
            .O(N__18542),
            .I(N__18539));
    CascadeMux I__4203 (
            .O(N__18539),
            .I(N__18536));
    CascadeBuf I__4202 (
            .O(N__18536),
            .I(N__18533));
    CascadeMux I__4201 (
            .O(N__18533),
            .I(N__18530));
    CascadeBuf I__4200 (
            .O(N__18530),
            .I(N__18527));
    CascadeMux I__4199 (
            .O(N__18527),
            .I(N__18524));
    CascadeBuf I__4198 (
            .O(N__18524),
            .I(N__18521));
    CascadeMux I__4197 (
            .O(N__18521),
            .I(N__18518));
    CascadeBuf I__4196 (
            .O(N__18518),
            .I(N__18515));
    CascadeMux I__4195 (
            .O(N__18515),
            .I(N__18512));
    CascadeBuf I__4194 (
            .O(N__18512),
            .I(N__18509));
    CascadeMux I__4193 (
            .O(N__18509),
            .I(N__18506));
    CascadeBuf I__4192 (
            .O(N__18506),
            .I(N__18503));
    CascadeMux I__4191 (
            .O(N__18503),
            .I(N__18500));
    CascadeBuf I__4190 (
            .O(N__18500),
            .I(N__18497));
    CascadeMux I__4189 (
            .O(N__18497),
            .I(N__18494));
    CascadeBuf I__4188 (
            .O(N__18494),
            .I(N__18491));
    CascadeMux I__4187 (
            .O(N__18491),
            .I(N__18488));
    CascadeBuf I__4186 (
            .O(N__18488),
            .I(N__18485));
    CascadeMux I__4185 (
            .O(N__18485),
            .I(N__18482));
    CascadeBuf I__4184 (
            .O(N__18482),
            .I(N__18479));
    CascadeMux I__4183 (
            .O(N__18479),
            .I(N__18476));
    CascadeBuf I__4182 (
            .O(N__18476),
            .I(N__18473));
    CascadeMux I__4181 (
            .O(N__18473),
            .I(N__18470));
    CascadeBuf I__4180 (
            .O(N__18470),
            .I(N__18467));
    CascadeMux I__4179 (
            .O(N__18467),
            .I(N__18464));
    InMux I__4178 (
            .O(N__18464),
            .I(N__18461));
    LocalMux I__4177 (
            .O(N__18461),
            .I(N__18458));
    Span4Mux_v I__4176 (
            .O(N__18458),
            .I(N__18455));
    Span4Mux_h I__4175 (
            .O(N__18455),
            .I(N__18452));
    Sp12to4 I__4174 (
            .O(N__18452),
            .I(N__18449));
    Odrv12 I__4173 (
            .O(N__18449),
            .I(M_this_ppu_sprites_addr_3));
    InMux I__4172 (
            .O(N__18446),
            .I(\this_ppu.sprites_addr_cry_2 ));
    CascadeMux I__4171 (
            .O(N__18443),
            .I(N__18440));
    InMux I__4170 (
            .O(N__18440),
            .I(N__18437));
    LocalMux I__4169 (
            .O(N__18437),
            .I(N__18434));
    Sp12to4 I__4168 (
            .O(N__18434),
            .I(N__18427));
    InMux I__4167 (
            .O(N__18433),
            .I(N__18424));
    InMux I__4166 (
            .O(N__18432),
            .I(N__18421));
    InMux I__4165 (
            .O(N__18431),
            .I(N__18418));
    CascadeMux I__4164 (
            .O(N__18430),
            .I(N__18415));
    Span12Mux_h I__4163 (
            .O(N__18427),
            .I(N__18412));
    LocalMux I__4162 (
            .O(N__18424),
            .I(N__18405));
    LocalMux I__4161 (
            .O(N__18421),
            .I(N__18405));
    LocalMux I__4160 (
            .O(N__18418),
            .I(N__18405));
    InMux I__4159 (
            .O(N__18415),
            .I(N__18402));
    Odrv12 I__4158 (
            .O(N__18412),
            .I(M_this_ppu_vram_addr_4));
    Odrv12 I__4157 (
            .O(N__18405),
            .I(M_this_ppu_vram_addr_4));
    LocalMux I__4156 (
            .O(N__18402),
            .I(M_this_ppu_vram_addr_4));
    CascadeMux I__4155 (
            .O(N__18395),
            .I(N__18392));
    CascadeBuf I__4154 (
            .O(N__18392),
            .I(N__18389));
    CascadeMux I__4153 (
            .O(N__18389),
            .I(N__18386));
    CascadeBuf I__4152 (
            .O(N__18386),
            .I(N__18383));
    CascadeMux I__4151 (
            .O(N__18383),
            .I(N__18380));
    CascadeBuf I__4150 (
            .O(N__18380),
            .I(N__18377));
    CascadeMux I__4149 (
            .O(N__18377),
            .I(N__18374));
    CascadeBuf I__4148 (
            .O(N__18374),
            .I(N__18371));
    CascadeMux I__4147 (
            .O(N__18371),
            .I(N__18368));
    CascadeBuf I__4146 (
            .O(N__18368),
            .I(N__18365));
    CascadeMux I__4145 (
            .O(N__18365),
            .I(N__18362));
    CascadeBuf I__4144 (
            .O(N__18362),
            .I(N__18359));
    CascadeMux I__4143 (
            .O(N__18359),
            .I(N__18356));
    CascadeBuf I__4142 (
            .O(N__18356),
            .I(N__18353));
    CascadeMux I__4141 (
            .O(N__18353),
            .I(N__18350));
    CascadeBuf I__4140 (
            .O(N__18350),
            .I(N__18347));
    CascadeMux I__4139 (
            .O(N__18347),
            .I(N__18344));
    CascadeBuf I__4138 (
            .O(N__18344),
            .I(N__18341));
    CascadeMux I__4137 (
            .O(N__18341),
            .I(N__18338));
    CascadeBuf I__4136 (
            .O(N__18338),
            .I(N__18335));
    CascadeMux I__4135 (
            .O(N__18335),
            .I(N__18332));
    CascadeBuf I__4134 (
            .O(N__18332),
            .I(N__18329));
    CascadeMux I__4133 (
            .O(N__18329),
            .I(N__18326));
    CascadeBuf I__4132 (
            .O(N__18326),
            .I(N__18323));
    CascadeMux I__4131 (
            .O(N__18323),
            .I(N__18320));
    CascadeBuf I__4130 (
            .O(N__18320),
            .I(N__18317));
    CascadeMux I__4129 (
            .O(N__18317),
            .I(N__18314));
    CascadeBuf I__4128 (
            .O(N__18314),
            .I(N__18311));
    CascadeMux I__4127 (
            .O(N__18311),
            .I(N__18308));
    CascadeBuf I__4126 (
            .O(N__18308),
            .I(N__18305));
    CascadeMux I__4125 (
            .O(N__18305),
            .I(N__18302));
    InMux I__4124 (
            .O(N__18302),
            .I(N__18299));
    LocalMux I__4123 (
            .O(N__18299),
            .I(N__18296));
    Span4Mux_s3_v I__4122 (
            .O(N__18296),
            .I(N__18293));
    Span4Mux_h I__4121 (
            .O(N__18293),
            .I(N__18290));
    Sp12to4 I__4120 (
            .O(N__18290),
            .I(N__18287));
    Odrv12 I__4119 (
            .O(N__18287),
            .I(M_this_ppu_sprites_addr_4));
    InMux I__4118 (
            .O(N__18284),
            .I(\this_ppu.sprites_addr_cry_3 ));
    CascadeMux I__4117 (
            .O(N__18281),
            .I(N__18278));
    InMux I__4116 (
            .O(N__18278),
            .I(N__18275));
    LocalMux I__4115 (
            .O(N__18275),
            .I(N__18271));
    InMux I__4114 (
            .O(N__18274),
            .I(N__18266));
    Span12Mux_h I__4113 (
            .O(N__18271),
            .I(N__18262));
    InMux I__4112 (
            .O(N__18270),
            .I(N__18257));
    InMux I__4111 (
            .O(N__18269),
            .I(N__18257));
    LocalMux I__4110 (
            .O(N__18266),
            .I(N__18254));
    InMux I__4109 (
            .O(N__18265),
            .I(N__18251));
    Odrv12 I__4108 (
            .O(N__18262),
            .I(M_this_ppu_vram_addr_5));
    LocalMux I__4107 (
            .O(N__18257),
            .I(M_this_ppu_vram_addr_5));
    Odrv4 I__4106 (
            .O(N__18254),
            .I(M_this_ppu_vram_addr_5));
    LocalMux I__4105 (
            .O(N__18251),
            .I(M_this_ppu_vram_addr_5));
    CascadeMux I__4104 (
            .O(N__18242),
            .I(N__18239));
    CascadeBuf I__4103 (
            .O(N__18239),
            .I(N__18236));
    CascadeMux I__4102 (
            .O(N__18236),
            .I(N__18233));
    CascadeBuf I__4101 (
            .O(N__18233),
            .I(N__18230));
    CascadeMux I__4100 (
            .O(N__18230),
            .I(N__18227));
    CascadeBuf I__4099 (
            .O(N__18227),
            .I(N__18224));
    CascadeMux I__4098 (
            .O(N__18224),
            .I(N__18221));
    CascadeBuf I__4097 (
            .O(N__18221),
            .I(N__18218));
    CascadeMux I__4096 (
            .O(N__18218),
            .I(N__18215));
    CascadeBuf I__4095 (
            .O(N__18215),
            .I(N__18212));
    CascadeMux I__4094 (
            .O(N__18212),
            .I(N__18209));
    CascadeBuf I__4093 (
            .O(N__18209),
            .I(N__18206));
    CascadeMux I__4092 (
            .O(N__18206),
            .I(N__18203));
    CascadeBuf I__4091 (
            .O(N__18203),
            .I(N__18200));
    CascadeMux I__4090 (
            .O(N__18200),
            .I(N__18197));
    CascadeBuf I__4089 (
            .O(N__18197),
            .I(N__18194));
    CascadeMux I__4088 (
            .O(N__18194),
            .I(N__18191));
    CascadeBuf I__4087 (
            .O(N__18191),
            .I(N__18188));
    CascadeMux I__4086 (
            .O(N__18188),
            .I(N__18185));
    CascadeBuf I__4085 (
            .O(N__18185),
            .I(N__18182));
    CascadeMux I__4084 (
            .O(N__18182),
            .I(N__18179));
    CascadeBuf I__4083 (
            .O(N__18179),
            .I(N__18176));
    CascadeMux I__4082 (
            .O(N__18176),
            .I(N__18173));
    CascadeBuf I__4081 (
            .O(N__18173),
            .I(N__18170));
    CascadeMux I__4080 (
            .O(N__18170),
            .I(N__18167));
    CascadeBuf I__4079 (
            .O(N__18167),
            .I(N__18164));
    CascadeMux I__4078 (
            .O(N__18164),
            .I(N__18161));
    CascadeBuf I__4077 (
            .O(N__18161),
            .I(N__18158));
    CascadeMux I__4076 (
            .O(N__18158),
            .I(N__18155));
    CascadeBuf I__4075 (
            .O(N__18155),
            .I(N__18152));
    CascadeMux I__4074 (
            .O(N__18152),
            .I(N__18149));
    InMux I__4073 (
            .O(N__18149),
            .I(N__18146));
    LocalMux I__4072 (
            .O(N__18146),
            .I(N__18143));
    Sp12to4 I__4071 (
            .O(N__18143),
            .I(N__18140));
    Span12Mux_s3_v I__4070 (
            .O(N__18140),
            .I(N__18137));
    Span12Mux_v I__4069 (
            .O(N__18137),
            .I(N__18134));
    Odrv12 I__4068 (
            .O(N__18134),
            .I(M_this_ppu_sprites_addr_5));
    InMux I__4067 (
            .O(N__18131),
            .I(\this_ppu.sprites_addr_cry_4 ));
    CascadeMux I__4066 (
            .O(N__18128),
            .I(N__18125));
    InMux I__4065 (
            .O(N__18125),
            .I(N__18122));
    LocalMux I__4064 (
            .O(N__18122),
            .I(N__18119));
    Span4Mux_h I__4063 (
            .O(N__18119),
            .I(N__18116));
    Sp12to4 I__4062 (
            .O(N__18116),
            .I(N__18110));
    CascadeMux I__4061 (
            .O(N__18115),
            .I(N__18107));
    InMux I__4060 (
            .O(N__18114),
            .I(N__18104));
    InMux I__4059 (
            .O(N__18113),
            .I(N__18101));
    Span12Mux_v I__4058 (
            .O(N__18110),
            .I(N__18098));
    InMux I__4057 (
            .O(N__18107),
            .I(N__18095));
    LocalMux I__4056 (
            .O(N__18104),
            .I(N__18090));
    LocalMux I__4055 (
            .O(N__18101),
            .I(N__18090));
    Odrv12 I__4054 (
            .O(N__18098),
            .I(M_this_ppu_vram_addr_6));
    LocalMux I__4053 (
            .O(N__18095),
            .I(M_this_ppu_vram_addr_6));
    Odrv4 I__4052 (
            .O(N__18090),
            .I(M_this_ppu_vram_addr_6));
    CascadeMux I__4051 (
            .O(N__18083),
            .I(N__18080));
    CascadeBuf I__4050 (
            .O(N__18080),
            .I(N__18077));
    CascadeMux I__4049 (
            .O(N__18077),
            .I(N__18074));
    CascadeBuf I__4048 (
            .O(N__18074),
            .I(N__18071));
    CascadeMux I__4047 (
            .O(N__18071),
            .I(N__18068));
    CascadeBuf I__4046 (
            .O(N__18068),
            .I(N__18065));
    CascadeMux I__4045 (
            .O(N__18065),
            .I(N__18062));
    CascadeBuf I__4044 (
            .O(N__18062),
            .I(N__18059));
    CascadeMux I__4043 (
            .O(N__18059),
            .I(N__18056));
    CascadeBuf I__4042 (
            .O(N__18056),
            .I(N__18053));
    CascadeMux I__4041 (
            .O(N__18053),
            .I(N__18050));
    CascadeBuf I__4040 (
            .O(N__18050),
            .I(N__18047));
    CascadeMux I__4039 (
            .O(N__18047),
            .I(N__18044));
    CascadeBuf I__4038 (
            .O(N__18044),
            .I(N__18041));
    CascadeMux I__4037 (
            .O(N__18041),
            .I(N__18038));
    CascadeBuf I__4036 (
            .O(N__18038),
            .I(N__18035));
    CascadeMux I__4035 (
            .O(N__18035),
            .I(N__18032));
    CascadeBuf I__4034 (
            .O(N__18032),
            .I(N__18029));
    CascadeMux I__4033 (
            .O(N__18029),
            .I(N__18026));
    CascadeBuf I__4032 (
            .O(N__18026),
            .I(N__18023));
    CascadeMux I__4031 (
            .O(N__18023),
            .I(N__18020));
    CascadeBuf I__4030 (
            .O(N__18020),
            .I(N__18017));
    CascadeMux I__4029 (
            .O(N__18017),
            .I(N__18014));
    CascadeBuf I__4028 (
            .O(N__18014),
            .I(N__18011));
    CascadeMux I__4027 (
            .O(N__18011),
            .I(N__18008));
    CascadeBuf I__4026 (
            .O(N__18008),
            .I(N__18005));
    CascadeMux I__4025 (
            .O(N__18005),
            .I(N__18002));
    CascadeBuf I__4024 (
            .O(N__18002),
            .I(N__17999));
    CascadeMux I__4023 (
            .O(N__17999),
            .I(N__17996));
    CascadeBuf I__4022 (
            .O(N__17996),
            .I(N__17993));
    CascadeMux I__4021 (
            .O(N__17993),
            .I(N__17990));
    InMux I__4020 (
            .O(N__17990),
            .I(N__17987));
    LocalMux I__4019 (
            .O(N__17987),
            .I(N__17984));
    Span4Mux_v I__4018 (
            .O(N__17984),
            .I(N__17981));
    Span4Mux_h I__4017 (
            .O(N__17981),
            .I(N__17978));
    Span4Mux_v I__4016 (
            .O(N__17978),
            .I(N__17975));
    Span4Mux_v I__4015 (
            .O(N__17975),
            .I(N__17972));
    Odrv4 I__4014 (
            .O(N__17972),
            .I(M_this_ppu_sprites_addr_6));
    InMux I__4013 (
            .O(N__17969),
            .I(\this_ppu.sprites_addr_cry_5 ));
    CascadeMux I__4012 (
            .O(N__17966),
            .I(N__17963));
    InMux I__4011 (
            .O(N__17963),
            .I(N__17960));
    LocalMux I__4010 (
            .O(N__17960),
            .I(N__17956));
    InMux I__4009 (
            .O(N__17959),
            .I(N__17953));
    Span4Mux_h I__4008 (
            .O(N__17956),
            .I(N__17950));
    LocalMux I__4007 (
            .O(N__17953),
            .I(N__17947));
    Span4Mux_v I__4006 (
            .O(N__17950),
            .I(N__17944));
    Span4Mux_h I__4005 (
            .O(N__17947),
            .I(N__17940));
    Span4Mux_h I__4004 (
            .O(N__17944),
            .I(N__17936));
    InMux I__4003 (
            .O(N__17943),
            .I(N__17933));
    Span4Mux_h I__4002 (
            .O(N__17940),
            .I(N__17930));
    InMux I__4001 (
            .O(N__17939),
            .I(N__17927));
    Odrv4 I__4000 (
            .O(N__17936),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__3999 (
            .O(N__17933),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__3998 (
            .O(N__17930),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__3997 (
            .O(N__17927),
            .I(M_this_ppu_vram_addr_7));
    CascadeMux I__3996 (
            .O(N__17918),
            .I(N__17915));
    CascadeBuf I__3995 (
            .O(N__17915),
            .I(N__17912));
    CascadeMux I__3994 (
            .O(N__17912),
            .I(N__17909));
    CascadeBuf I__3993 (
            .O(N__17909),
            .I(N__17906));
    CascadeMux I__3992 (
            .O(N__17906),
            .I(N__17903));
    CascadeBuf I__3991 (
            .O(N__17903),
            .I(N__17900));
    CascadeMux I__3990 (
            .O(N__17900),
            .I(N__17897));
    CascadeBuf I__3989 (
            .O(N__17897),
            .I(N__17894));
    CascadeMux I__3988 (
            .O(N__17894),
            .I(N__17891));
    CascadeBuf I__3987 (
            .O(N__17891),
            .I(N__17888));
    CascadeMux I__3986 (
            .O(N__17888),
            .I(N__17885));
    CascadeBuf I__3985 (
            .O(N__17885),
            .I(N__17882));
    CascadeMux I__3984 (
            .O(N__17882),
            .I(N__17879));
    CascadeBuf I__3983 (
            .O(N__17879),
            .I(N__17876));
    CascadeMux I__3982 (
            .O(N__17876),
            .I(N__17873));
    CascadeBuf I__3981 (
            .O(N__17873),
            .I(N__17870));
    CascadeMux I__3980 (
            .O(N__17870),
            .I(N__17867));
    CascadeBuf I__3979 (
            .O(N__17867),
            .I(N__17864));
    CascadeMux I__3978 (
            .O(N__17864),
            .I(N__17861));
    CascadeBuf I__3977 (
            .O(N__17861),
            .I(N__17858));
    CascadeMux I__3976 (
            .O(N__17858),
            .I(N__17855));
    CascadeBuf I__3975 (
            .O(N__17855),
            .I(N__17852));
    CascadeMux I__3974 (
            .O(N__17852),
            .I(N__17849));
    CascadeBuf I__3973 (
            .O(N__17849),
            .I(N__17846));
    CascadeMux I__3972 (
            .O(N__17846),
            .I(N__17843));
    CascadeBuf I__3971 (
            .O(N__17843),
            .I(N__17840));
    CascadeMux I__3970 (
            .O(N__17840),
            .I(N__17837));
    CascadeBuf I__3969 (
            .O(N__17837),
            .I(N__17834));
    CascadeMux I__3968 (
            .O(N__17834),
            .I(N__17831));
    CascadeBuf I__3967 (
            .O(N__17831),
            .I(N__17828));
    CascadeMux I__3966 (
            .O(N__17828),
            .I(N__17825));
    InMux I__3965 (
            .O(N__17825),
            .I(N__17822));
    LocalMux I__3964 (
            .O(N__17822),
            .I(N__17819));
    Span4Mux_v I__3963 (
            .O(N__17819),
            .I(N__17816));
    Span4Mux_h I__3962 (
            .O(N__17816),
            .I(N__17813));
    Span4Mux_v I__3961 (
            .O(N__17813),
            .I(N__17810));
    Span4Mux_v I__3960 (
            .O(N__17810),
            .I(N__17807));
    Odrv4 I__3959 (
            .O(N__17807),
            .I(M_this_ppu_sprites_addr_7));
    InMux I__3958 (
            .O(N__17804),
            .I(\this_ppu.sprites_addr_cry_6 ));
    InMux I__3957 (
            .O(N__17801),
            .I(N__17798));
    LocalMux I__3956 (
            .O(N__17798),
            .I(N__17793));
    InMux I__3955 (
            .O(N__17797),
            .I(N__17789));
    InMux I__3954 (
            .O(N__17796),
            .I(N__17786));
    Span4Mux_v I__3953 (
            .O(N__17793),
            .I(N__17783));
    InMux I__3952 (
            .O(N__17792),
            .I(N__17780));
    LocalMux I__3951 (
            .O(N__17789),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    LocalMux I__3950 (
            .O(N__17786),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv4 I__3949 (
            .O(N__17783),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    LocalMux I__3948 (
            .O(N__17780),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    CascadeMux I__3947 (
            .O(N__17771),
            .I(N__17768));
    CascadeBuf I__3946 (
            .O(N__17768),
            .I(N__17765));
    CascadeMux I__3945 (
            .O(N__17765),
            .I(N__17762));
    CascadeBuf I__3944 (
            .O(N__17762),
            .I(N__17759));
    CascadeMux I__3943 (
            .O(N__17759),
            .I(N__17756));
    CascadeBuf I__3942 (
            .O(N__17756),
            .I(N__17753));
    CascadeMux I__3941 (
            .O(N__17753),
            .I(N__17750));
    CascadeBuf I__3940 (
            .O(N__17750),
            .I(N__17747));
    CascadeMux I__3939 (
            .O(N__17747),
            .I(N__17744));
    CascadeBuf I__3938 (
            .O(N__17744),
            .I(N__17741));
    CascadeMux I__3937 (
            .O(N__17741),
            .I(N__17738));
    CascadeBuf I__3936 (
            .O(N__17738),
            .I(N__17735));
    CascadeMux I__3935 (
            .O(N__17735),
            .I(N__17732));
    CascadeBuf I__3934 (
            .O(N__17732),
            .I(N__17729));
    CascadeMux I__3933 (
            .O(N__17729),
            .I(N__17726));
    CascadeBuf I__3932 (
            .O(N__17726),
            .I(N__17723));
    CascadeMux I__3931 (
            .O(N__17723),
            .I(N__17720));
    CascadeBuf I__3930 (
            .O(N__17720),
            .I(N__17717));
    CascadeMux I__3929 (
            .O(N__17717),
            .I(N__17714));
    CascadeBuf I__3928 (
            .O(N__17714),
            .I(N__17711));
    CascadeMux I__3927 (
            .O(N__17711),
            .I(N__17708));
    CascadeBuf I__3926 (
            .O(N__17708),
            .I(N__17705));
    CascadeMux I__3925 (
            .O(N__17705),
            .I(N__17702));
    CascadeBuf I__3924 (
            .O(N__17702),
            .I(N__17699));
    CascadeMux I__3923 (
            .O(N__17699),
            .I(N__17696));
    CascadeBuf I__3922 (
            .O(N__17696),
            .I(N__17693));
    CascadeMux I__3921 (
            .O(N__17693),
            .I(N__17690));
    CascadeBuf I__3920 (
            .O(N__17690),
            .I(N__17687));
    CascadeMux I__3919 (
            .O(N__17687),
            .I(N__17684));
    CascadeBuf I__3918 (
            .O(N__17684),
            .I(N__17681));
    CascadeMux I__3917 (
            .O(N__17681),
            .I(N__17678));
    InMux I__3916 (
            .O(N__17678),
            .I(N__17675));
    LocalMux I__3915 (
            .O(N__17675),
            .I(N__17672));
    Span4Mux_v I__3914 (
            .O(N__17672),
            .I(N__17669));
    Span4Mux_h I__3913 (
            .O(N__17669),
            .I(N__17666));
    Span4Mux_v I__3912 (
            .O(N__17666),
            .I(N__17663));
    Span4Mux_v I__3911 (
            .O(N__17663),
            .I(N__17660));
    Odrv4 I__3910 (
            .O(N__17660),
            .I(M_this_ppu_sprites_addr_8));
    InMux I__3909 (
            .O(N__17657),
            .I(\this_ppu.sprites_addr_cry_7 ));
    CascadeMux I__3908 (
            .O(N__17654),
            .I(N__17650));
    InMux I__3907 (
            .O(N__17653),
            .I(N__17647));
    InMux I__3906 (
            .O(N__17650),
            .I(N__17643));
    LocalMux I__3905 (
            .O(N__17647),
            .I(N__17640));
    InMux I__3904 (
            .O(N__17646),
            .I(N__17637));
    LocalMux I__3903 (
            .O(N__17643),
            .I(\this_ppu.M_vaddress_qZ1Z_2 ));
    Odrv12 I__3902 (
            .O(N__17640),
            .I(\this_ppu.M_vaddress_qZ1Z_2 ));
    LocalMux I__3901 (
            .O(N__17637),
            .I(\this_ppu.M_vaddress_qZ1Z_2 ));
    CascadeMux I__3900 (
            .O(N__17630),
            .I(N__17627));
    CascadeBuf I__3899 (
            .O(N__17627),
            .I(N__17624));
    CascadeMux I__3898 (
            .O(N__17624),
            .I(N__17621));
    CascadeBuf I__3897 (
            .O(N__17621),
            .I(N__17618));
    CascadeMux I__3896 (
            .O(N__17618),
            .I(N__17615));
    CascadeBuf I__3895 (
            .O(N__17615),
            .I(N__17612));
    CascadeMux I__3894 (
            .O(N__17612),
            .I(N__17609));
    CascadeBuf I__3893 (
            .O(N__17609),
            .I(N__17606));
    CascadeMux I__3892 (
            .O(N__17606),
            .I(N__17603));
    CascadeBuf I__3891 (
            .O(N__17603),
            .I(N__17600));
    CascadeMux I__3890 (
            .O(N__17600),
            .I(N__17597));
    CascadeBuf I__3889 (
            .O(N__17597),
            .I(N__17594));
    CascadeMux I__3888 (
            .O(N__17594),
            .I(N__17591));
    CascadeBuf I__3887 (
            .O(N__17591),
            .I(N__17588));
    CascadeMux I__3886 (
            .O(N__17588),
            .I(N__17585));
    CascadeBuf I__3885 (
            .O(N__17585),
            .I(N__17582));
    CascadeMux I__3884 (
            .O(N__17582),
            .I(N__17579));
    CascadeBuf I__3883 (
            .O(N__17579),
            .I(N__17576));
    CascadeMux I__3882 (
            .O(N__17576),
            .I(N__17573));
    CascadeBuf I__3881 (
            .O(N__17573),
            .I(N__17570));
    CascadeMux I__3880 (
            .O(N__17570),
            .I(N__17567));
    CascadeBuf I__3879 (
            .O(N__17567),
            .I(N__17564));
    CascadeMux I__3878 (
            .O(N__17564),
            .I(N__17561));
    CascadeBuf I__3877 (
            .O(N__17561),
            .I(N__17558));
    CascadeMux I__3876 (
            .O(N__17558),
            .I(N__17555));
    CascadeBuf I__3875 (
            .O(N__17555),
            .I(N__17552));
    CascadeMux I__3874 (
            .O(N__17552),
            .I(N__17549));
    CascadeBuf I__3873 (
            .O(N__17549),
            .I(N__17546));
    CascadeMux I__3872 (
            .O(N__17546),
            .I(N__17543));
    CascadeBuf I__3871 (
            .O(N__17543),
            .I(N__17540));
    CascadeMux I__3870 (
            .O(N__17540),
            .I(N__17537));
    InMux I__3869 (
            .O(N__17537),
            .I(N__17534));
    LocalMux I__3868 (
            .O(N__17534),
            .I(N__17531));
    Span4Mux_s2_v I__3867 (
            .O(N__17531),
            .I(N__17528));
    Span4Mux_v I__3866 (
            .O(N__17528),
            .I(N__17525));
    Span4Mux_v I__3865 (
            .O(N__17525),
            .I(N__17522));
    Span4Mux_v I__3864 (
            .O(N__17522),
            .I(N__17519));
    Odrv4 I__3863 (
            .O(N__17519),
            .I(M_this_ppu_sprites_addr_9));
    InMux I__3862 (
            .O(N__17516),
            .I(bfn_21_18_0_));
    InMux I__3861 (
            .O(N__17513),
            .I(N__17499));
    InMux I__3860 (
            .O(N__17512),
            .I(N__17499));
    InMux I__3859 (
            .O(N__17511),
            .I(N__17496));
    InMux I__3858 (
            .O(N__17510),
            .I(N__17491));
    InMux I__3857 (
            .O(N__17509),
            .I(N__17484));
    InMux I__3856 (
            .O(N__17508),
            .I(N__17484));
    InMux I__3855 (
            .O(N__17507),
            .I(N__17484));
    InMux I__3854 (
            .O(N__17506),
            .I(N__17479));
    InMux I__3853 (
            .O(N__17505),
            .I(N__17474));
    InMux I__3852 (
            .O(N__17504),
            .I(N__17474));
    LocalMux I__3851 (
            .O(N__17499),
            .I(N__17469));
    LocalMux I__3850 (
            .O(N__17496),
            .I(N__17469));
    InMux I__3849 (
            .O(N__17495),
            .I(N__17464));
    InMux I__3848 (
            .O(N__17494),
            .I(N__17464));
    LocalMux I__3847 (
            .O(N__17491),
            .I(N__17459));
    LocalMux I__3846 (
            .O(N__17484),
            .I(N__17459));
    InMux I__3845 (
            .O(N__17483),
            .I(N__17454));
    InMux I__3844 (
            .O(N__17482),
            .I(N__17454));
    LocalMux I__3843 (
            .O(N__17479),
            .I(N__17451));
    LocalMux I__3842 (
            .O(N__17474),
            .I(N__17448));
    Span4Mux_v I__3841 (
            .O(N__17469),
            .I(N__17439));
    LocalMux I__3840 (
            .O(N__17464),
            .I(N__17439));
    Span4Mux_v I__3839 (
            .O(N__17459),
            .I(N__17439));
    LocalMux I__3838 (
            .O(N__17454),
            .I(N__17439));
    Odrv4 I__3837 (
            .O(N__17451),
            .I(M_this_sprites_address_q_3_sm0_0));
    Odrv4 I__3836 (
            .O(N__17448),
            .I(M_this_sprites_address_q_3_sm0_0));
    Odrv4 I__3835 (
            .O(N__17439),
            .I(M_this_sprites_address_q_3_sm0_0));
    CascadeMux I__3834 (
            .O(N__17432),
            .I(M_this_sprites_address_q_3_ns_1_3_cascade_));
    InMux I__3833 (
            .O(N__17429),
            .I(N__17426));
    LocalMux I__3832 (
            .O(N__17426),
            .I(N__17423));
    Span12Mux_s10_v I__3831 (
            .O(N__17423),
            .I(N__17420));
    Odrv12 I__3830 (
            .O(N__17420),
            .I(M_this_sprites_address_q_RNO_1Z0Z_3));
    CascadeMux I__3829 (
            .O(N__17417),
            .I(N__17414));
    CascadeBuf I__3828 (
            .O(N__17414),
            .I(N__17411));
    CascadeMux I__3827 (
            .O(N__17411),
            .I(N__17408));
    CascadeBuf I__3826 (
            .O(N__17408),
            .I(N__17405));
    CascadeMux I__3825 (
            .O(N__17405),
            .I(N__17402));
    CascadeBuf I__3824 (
            .O(N__17402),
            .I(N__17399));
    CascadeMux I__3823 (
            .O(N__17399),
            .I(N__17396));
    CascadeBuf I__3822 (
            .O(N__17396),
            .I(N__17393));
    CascadeMux I__3821 (
            .O(N__17393),
            .I(N__17390));
    CascadeBuf I__3820 (
            .O(N__17390),
            .I(N__17387));
    CascadeMux I__3819 (
            .O(N__17387),
            .I(N__17384));
    CascadeBuf I__3818 (
            .O(N__17384),
            .I(N__17381));
    CascadeMux I__3817 (
            .O(N__17381),
            .I(N__17378));
    CascadeBuf I__3816 (
            .O(N__17378),
            .I(N__17375));
    CascadeMux I__3815 (
            .O(N__17375),
            .I(N__17372));
    CascadeBuf I__3814 (
            .O(N__17372),
            .I(N__17369));
    CascadeMux I__3813 (
            .O(N__17369),
            .I(N__17366));
    CascadeBuf I__3812 (
            .O(N__17366),
            .I(N__17363));
    CascadeMux I__3811 (
            .O(N__17363),
            .I(N__17360));
    CascadeBuf I__3810 (
            .O(N__17360),
            .I(N__17357));
    CascadeMux I__3809 (
            .O(N__17357),
            .I(N__17354));
    CascadeBuf I__3808 (
            .O(N__17354),
            .I(N__17351));
    CascadeMux I__3807 (
            .O(N__17351),
            .I(N__17348));
    CascadeBuf I__3806 (
            .O(N__17348),
            .I(N__17345));
    CascadeMux I__3805 (
            .O(N__17345),
            .I(N__17342));
    CascadeBuf I__3804 (
            .O(N__17342),
            .I(N__17339));
    CascadeMux I__3803 (
            .O(N__17339),
            .I(N__17336));
    CascadeBuf I__3802 (
            .O(N__17336),
            .I(N__17333));
    CascadeMux I__3801 (
            .O(N__17333),
            .I(N__17330));
    CascadeBuf I__3800 (
            .O(N__17330),
            .I(N__17327));
    CascadeMux I__3799 (
            .O(N__17327),
            .I(N__17324));
    InMux I__3798 (
            .O(N__17324),
            .I(N__17320));
    InMux I__3797 (
            .O(N__17323),
            .I(N__17317));
    LocalMux I__3796 (
            .O(N__17320),
            .I(N__17314));
    LocalMux I__3795 (
            .O(N__17317),
            .I(N__17310));
    Span4Mux_s2_v I__3794 (
            .O(N__17314),
            .I(N__17307));
    CascadeMux I__3793 (
            .O(N__17313),
            .I(N__17304));
    Span4Mux_h I__3792 (
            .O(N__17310),
            .I(N__17301));
    Span4Mux_h I__3791 (
            .O(N__17307),
            .I(N__17298));
    InMux I__3790 (
            .O(N__17304),
            .I(N__17295));
    Span4Mux_h I__3789 (
            .O(N__17301),
            .I(N__17290));
    Span4Mux_v I__3788 (
            .O(N__17298),
            .I(N__17290));
    LocalMux I__3787 (
            .O(N__17295),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv4 I__3786 (
            .O(N__17290),
            .I(M_this_sprites_address_qZ0Z_3));
    InMux I__3785 (
            .O(N__17285),
            .I(N__17282));
    LocalMux I__3784 (
            .O(N__17282),
            .I(N__17279));
    Span4Mux_v I__3783 (
            .O(N__17279),
            .I(N__17276));
    Span4Mux_h I__3782 (
            .O(N__17276),
            .I(N__17273));
    Sp12to4 I__3781 (
            .O(N__17273),
            .I(N__17270));
    Odrv12 I__3780 (
            .O(N__17270),
            .I(\this_sprites_ram.mem_out_bus5_3 ));
    InMux I__3779 (
            .O(N__17267),
            .I(N__17264));
    LocalMux I__3778 (
            .O(N__17264),
            .I(N__17261));
    Span4Mux_h I__3777 (
            .O(N__17261),
            .I(N__17258));
    Odrv4 I__3776 (
            .O(N__17258),
            .I(\this_sprites_ram.mem_out_bus1_3 ));
    InMux I__3775 (
            .O(N__17255),
            .I(N__17252));
    LocalMux I__3774 (
            .O(N__17252),
            .I(N__17249));
    Span4Mux_h I__3773 (
            .O(N__17249),
            .I(N__17246));
    Span4Mux_h I__3772 (
            .O(N__17246),
            .I(N__17243));
    Odrv4 I__3771 (
            .O(N__17243),
            .I(\this_sprites_ram.mem_out_bus3_3 ));
    CascadeMux I__3770 (
            .O(N__17240),
            .I(N__17237));
    InMux I__3769 (
            .O(N__17237),
            .I(N__17234));
    LocalMux I__3768 (
            .O(N__17234),
            .I(N__17231));
    Span12Mux_h I__3767 (
            .O(N__17231),
            .I(N__17228));
    Span12Mux_v I__3766 (
            .O(N__17228),
            .I(N__17225));
    Odrv12 I__3765 (
            .O(N__17225),
            .I(\this_sprites_ram.mem_out_bus7_3 ));
    InMux I__3764 (
            .O(N__17222),
            .I(N__17219));
    LocalMux I__3763 (
            .O(N__17219),
            .I(\this_sprites_ram.mem_DOUT_6_i_m2_ns_1_3 ));
    InMux I__3762 (
            .O(N__17216),
            .I(N__17213));
    LocalMux I__3761 (
            .O(N__17213),
            .I(this_sprites_ram_mem_N_102));
    InMux I__3760 (
            .O(N__17210),
            .I(N__17207));
    LocalMux I__3759 (
            .O(N__17207),
            .I(N__17204));
    Span4Mux_v I__3758 (
            .O(N__17204),
            .I(N__17201));
    Span4Mux_h I__3757 (
            .O(N__17201),
            .I(N__17198));
    Sp12to4 I__3756 (
            .O(N__17198),
            .I(N__17195));
    Odrv12 I__3755 (
            .O(N__17195),
            .I(M_this_ppu_vram_data_1));
    InMux I__3754 (
            .O(N__17192),
            .I(N__17189));
    LocalMux I__3753 (
            .O(N__17189),
            .I(N__17186));
    Span4Mux_v I__3752 (
            .O(N__17186),
            .I(N__17183));
    Span4Mux_h I__3751 (
            .O(N__17183),
            .I(N__17180));
    Odrv4 I__3750 (
            .O(N__17180),
            .I(\this_sprites_ram.mem_out_bus2_1 ));
    CascadeMux I__3749 (
            .O(N__17177),
            .I(N__17174));
    InMux I__3748 (
            .O(N__17174),
            .I(N__17171));
    LocalMux I__3747 (
            .O(N__17171),
            .I(N__17168));
    Span4Mux_v I__3746 (
            .O(N__17168),
            .I(N__17165));
    Span4Mux_v I__3745 (
            .O(N__17165),
            .I(N__17162));
    Span4Mux_h I__3744 (
            .O(N__17162),
            .I(N__17159));
    Odrv4 I__3743 (
            .O(N__17159),
            .I(\this_sprites_ram.mem_out_bus6_1 ));
    InMux I__3742 (
            .O(N__17156),
            .I(N__17153));
    LocalMux I__3741 (
            .O(N__17153),
            .I(this_sprites_ram_mem_N_91));
    InMux I__3740 (
            .O(N__17150),
            .I(N__17147));
    LocalMux I__3739 (
            .O(N__17147),
            .I(N__17144));
    Span4Mux_h I__3738 (
            .O(N__17144),
            .I(N__17141));
    Odrv4 I__3737 (
            .O(N__17141),
            .I(\this_sprites_ram.mem_out_bus4_1 ));
    InMux I__3736 (
            .O(N__17138),
            .I(N__17135));
    LocalMux I__3735 (
            .O(N__17135),
            .I(N__17132));
    Span4Mux_h I__3734 (
            .O(N__17132),
            .I(N__17129));
    Sp12to4 I__3733 (
            .O(N__17129),
            .I(N__17126));
    Span12Mux_v I__3732 (
            .O(N__17126),
            .I(N__17123));
    Odrv12 I__3731 (
            .O(N__17123),
            .I(\this_sprites_ram.mem_out_bus0_1 ));
    InMux I__3730 (
            .O(N__17120),
            .I(N__17117));
    LocalMux I__3729 (
            .O(N__17117),
            .I(\this_sprites_ram.mem_DOUT_3_i_m2_ns_1_1 ));
    CascadeMux I__3728 (
            .O(N__17114),
            .I(N__17111));
    InMux I__3727 (
            .O(N__17111),
            .I(N__17108));
    LocalMux I__3726 (
            .O(N__17108),
            .I(N__17104));
    CascadeMux I__3725 (
            .O(N__17107),
            .I(N__17101));
    Span4Mux_v I__3724 (
            .O(N__17104),
            .I(N__17096));
    InMux I__3723 (
            .O(N__17101),
            .I(N__17093));
    InMux I__3722 (
            .O(N__17100),
            .I(N__17090));
    CascadeMux I__3721 (
            .O(N__17099),
            .I(N__17087));
    Sp12to4 I__3720 (
            .O(N__17096),
            .I(N__17082));
    LocalMux I__3719 (
            .O(N__17093),
            .I(N__17076));
    LocalMux I__3718 (
            .O(N__17090),
            .I(N__17076));
    InMux I__3717 (
            .O(N__17087),
            .I(N__17073));
    InMux I__3716 (
            .O(N__17086),
            .I(N__17070));
    InMux I__3715 (
            .O(N__17085),
            .I(N__17067));
    Span12Mux_h I__3714 (
            .O(N__17082),
            .I(N__17064));
    InMux I__3713 (
            .O(N__17081),
            .I(N__17061));
    Span4Mux_h I__3712 (
            .O(N__17076),
            .I(N__17056));
    LocalMux I__3711 (
            .O(N__17073),
            .I(N__17056));
    LocalMux I__3710 (
            .O(N__17070),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__3709 (
            .O(N__17067),
            .I(M_this_ppu_vram_addr_1));
    Odrv12 I__3708 (
            .O(N__17064),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__3707 (
            .O(N__17061),
            .I(M_this_ppu_vram_addr_1));
    Odrv4 I__3706 (
            .O(N__17056),
            .I(M_this_ppu_vram_addr_1));
    CascadeMux I__3705 (
            .O(N__17045),
            .I(N__17042));
    InMux I__3704 (
            .O(N__17042),
            .I(N__17039));
    LocalMux I__3703 (
            .O(N__17039),
            .I(N__17036));
    Span4Mux_v I__3702 (
            .O(N__17036),
            .I(N__17032));
    CascadeMux I__3701 (
            .O(N__17035),
            .I(N__17028));
    Sp12to4 I__3700 (
            .O(N__17032),
            .I(N__17022));
    InMux I__3699 (
            .O(N__17031),
            .I(N__17018));
    InMux I__3698 (
            .O(N__17028),
            .I(N__17013));
    InMux I__3697 (
            .O(N__17027),
            .I(N__17013));
    InMux I__3696 (
            .O(N__17026),
            .I(N__17010));
    InMux I__3695 (
            .O(N__17025),
            .I(N__17007));
    Span12Mux_h I__3694 (
            .O(N__17022),
            .I(N__17004));
    InMux I__3693 (
            .O(N__17021),
            .I(N__17001));
    LocalMux I__3692 (
            .O(N__17018),
            .I(N__16998));
    LocalMux I__3691 (
            .O(N__17013),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__3690 (
            .O(N__17010),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__3689 (
            .O(N__17007),
            .I(M_this_ppu_vram_addr_2));
    Odrv12 I__3688 (
            .O(N__17004),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__3687 (
            .O(N__17001),
            .I(M_this_ppu_vram_addr_2));
    Odrv4 I__3686 (
            .O(N__16998),
            .I(M_this_ppu_vram_addr_2));
    CascadeMux I__3685 (
            .O(N__16985),
            .I(N__16982));
    CascadeBuf I__3684 (
            .O(N__16982),
            .I(N__16979));
    CascadeMux I__3683 (
            .O(N__16979),
            .I(N__16976));
    CascadeBuf I__3682 (
            .O(N__16976),
            .I(N__16973));
    CascadeMux I__3681 (
            .O(N__16973),
            .I(N__16970));
    CascadeBuf I__3680 (
            .O(N__16970),
            .I(N__16967));
    CascadeMux I__3679 (
            .O(N__16967),
            .I(N__16964));
    CascadeBuf I__3678 (
            .O(N__16964),
            .I(N__16961));
    CascadeMux I__3677 (
            .O(N__16961),
            .I(N__16958));
    CascadeBuf I__3676 (
            .O(N__16958),
            .I(N__16955));
    CascadeMux I__3675 (
            .O(N__16955),
            .I(N__16952));
    CascadeBuf I__3674 (
            .O(N__16952),
            .I(N__16949));
    CascadeMux I__3673 (
            .O(N__16949),
            .I(N__16946));
    CascadeBuf I__3672 (
            .O(N__16946),
            .I(N__16943));
    CascadeMux I__3671 (
            .O(N__16943),
            .I(N__16940));
    CascadeBuf I__3670 (
            .O(N__16940),
            .I(N__16937));
    CascadeMux I__3669 (
            .O(N__16937),
            .I(N__16934));
    CascadeBuf I__3668 (
            .O(N__16934),
            .I(N__16931));
    CascadeMux I__3667 (
            .O(N__16931),
            .I(N__16928));
    CascadeBuf I__3666 (
            .O(N__16928),
            .I(N__16925));
    CascadeMux I__3665 (
            .O(N__16925),
            .I(N__16922));
    CascadeBuf I__3664 (
            .O(N__16922),
            .I(N__16919));
    CascadeMux I__3663 (
            .O(N__16919),
            .I(N__16916));
    CascadeBuf I__3662 (
            .O(N__16916),
            .I(N__16913));
    CascadeMux I__3661 (
            .O(N__16913),
            .I(N__16910));
    CascadeBuf I__3660 (
            .O(N__16910),
            .I(N__16907));
    CascadeMux I__3659 (
            .O(N__16907),
            .I(N__16904));
    CascadeBuf I__3658 (
            .O(N__16904),
            .I(N__16901));
    CascadeMux I__3657 (
            .O(N__16901),
            .I(N__16898));
    CascadeBuf I__3656 (
            .O(N__16898),
            .I(N__16895));
    CascadeMux I__3655 (
            .O(N__16895),
            .I(N__16892));
    InMux I__3654 (
            .O(N__16892),
            .I(N__16889));
    LocalMux I__3653 (
            .O(N__16889),
            .I(N__16886));
    Span4Mux_v I__3652 (
            .O(N__16886),
            .I(N__16883));
    Span4Mux_h I__3651 (
            .O(N__16883),
            .I(N__16880));
    Sp12to4 I__3650 (
            .O(N__16880),
            .I(N__16877));
    Odrv12 I__3649 (
            .O(N__16877),
            .I(M_this_ppu_sprites_addr_2));
    InMux I__3648 (
            .O(N__16874),
            .I(N__16871));
    LocalMux I__3647 (
            .O(N__16871),
            .I(\this_ppu.un1_M_vaddress_q_c5 ));
    InMux I__3646 (
            .O(N__16868),
            .I(N__16856));
    InMux I__3645 (
            .O(N__16867),
            .I(N__16856));
    InMux I__3644 (
            .O(N__16866),
            .I(N__16856));
    InMux I__3643 (
            .O(N__16865),
            .I(N__16851));
    InMux I__3642 (
            .O(N__16864),
            .I(N__16851));
    InMux I__3641 (
            .O(N__16863),
            .I(N__16847));
    LocalMux I__3640 (
            .O(N__16856),
            .I(N__16842));
    LocalMux I__3639 (
            .O(N__16851),
            .I(N__16842));
    InMux I__3638 (
            .O(N__16850),
            .I(N__16839));
    LocalMux I__3637 (
            .O(N__16847),
            .I(N__16832));
    Span4Mux_h I__3636 (
            .O(N__16842),
            .I(N__16832));
    LocalMux I__3635 (
            .O(N__16839),
            .I(N__16832));
    Odrv4 I__3634 (
            .O(N__16832),
            .I(\this_ppu.N_258_1 ));
    CascadeMux I__3633 (
            .O(N__16829),
            .I(\this_ppu.un1_M_vaddress_q_c5_cascade_ ));
    InMux I__3632 (
            .O(N__16826),
            .I(N__16823));
    LocalMux I__3631 (
            .O(N__16823),
            .I(N__16820));
    Odrv4 I__3630 (
            .O(N__16820),
            .I(\this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_13 ));
    CascadeMux I__3629 (
            .O(N__16817),
            .I(N__16814));
    CascadeBuf I__3628 (
            .O(N__16814),
            .I(N__16811));
    CascadeMux I__3627 (
            .O(N__16811),
            .I(N__16808));
    CascadeBuf I__3626 (
            .O(N__16808),
            .I(N__16805));
    CascadeMux I__3625 (
            .O(N__16805),
            .I(N__16802));
    CascadeBuf I__3624 (
            .O(N__16802),
            .I(N__16799));
    CascadeMux I__3623 (
            .O(N__16799),
            .I(N__16796));
    CascadeBuf I__3622 (
            .O(N__16796),
            .I(N__16793));
    CascadeMux I__3621 (
            .O(N__16793),
            .I(N__16790));
    CascadeBuf I__3620 (
            .O(N__16790),
            .I(N__16787));
    CascadeMux I__3619 (
            .O(N__16787),
            .I(N__16784));
    CascadeBuf I__3618 (
            .O(N__16784),
            .I(N__16781));
    CascadeMux I__3617 (
            .O(N__16781),
            .I(N__16778));
    CascadeBuf I__3616 (
            .O(N__16778),
            .I(N__16775));
    CascadeMux I__3615 (
            .O(N__16775),
            .I(N__16772));
    CascadeBuf I__3614 (
            .O(N__16772),
            .I(N__16769));
    CascadeMux I__3613 (
            .O(N__16769),
            .I(N__16766));
    CascadeBuf I__3612 (
            .O(N__16766),
            .I(N__16763));
    CascadeMux I__3611 (
            .O(N__16763),
            .I(N__16760));
    CascadeBuf I__3610 (
            .O(N__16760),
            .I(N__16757));
    CascadeMux I__3609 (
            .O(N__16757),
            .I(N__16754));
    CascadeBuf I__3608 (
            .O(N__16754),
            .I(N__16751));
    CascadeMux I__3607 (
            .O(N__16751),
            .I(N__16748));
    CascadeBuf I__3606 (
            .O(N__16748),
            .I(N__16745));
    CascadeMux I__3605 (
            .O(N__16745),
            .I(N__16742));
    CascadeBuf I__3604 (
            .O(N__16742),
            .I(N__16739));
    CascadeMux I__3603 (
            .O(N__16739),
            .I(N__16736));
    CascadeBuf I__3602 (
            .O(N__16736),
            .I(N__16733));
    CascadeMux I__3601 (
            .O(N__16733),
            .I(N__16730));
    CascadeBuf I__3600 (
            .O(N__16730),
            .I(N__16727));
    CascadeMux I__3599 (
            .O(N__16727),
            .I(N__16723));
    InMux I__3598 (
            .O(N__16726),
            .I(N__16720));
    InMux I__3597 (
            .O(N__16723),
            .I(N__16717));
    LocalMux I__3596 (
            .O(N__16720),
            .I(N__16713));
    LocalMux I__3595 (
            .O(N__16717),
            .I(N__16710));
    InMux I__3594 (
            .O(N__16716),
            .I(N__16707));
    Span4Mux_h I__3593 (
            .O(N__16713),
            .I(N__16704));
    Span12Mux_h I__3592 (
            .O(N__16710),
            .I(N__16701));
    LocalMux I__3591 (
            .O(N__16707),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv4 I__3590 (
            .O(N__16704),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv12 I__3589 (
            .O(N__16701),
            .I(M_this_sprites_address_qZ0Z_2));
    CascadeMux I__3588 (
            .O(N__16694),
            .I(N__16691));
    InMux I__3587 (
            .O(N__16691),
            .I(N__16688));
    LocalMux I__3586 (
            .O(N__16688),
            .I(N__16685));
    Span4Mux_v I__3585 (
            .O(N__16685),
            .I(N__16682));
    Span4Mux_h I__3584 (
            .O(N__16682),
            .I(N__16679));
    Odrv4 I__3583 (
            .O(N__16679),
            .I(M_this_sprites_address_q_3_ns_1_2));
    InMux I__3582 (
            .O(N__16676),
            .I(N__16673));
    LocalMux I__3581 (
            .O(N__16673),
            .I(N__16670));
    Span12Mux_h I__3580 (
            .O(N__16670),
            .I(N__16667));
    Odrv12 I__3579 (
            .O(N__16667),
            .I(M_this_ppu_vram_data_3));
    CascadeMux I__3578 (
            .O(N__16664),
            .I(N__16661));
    CascadeBuf I__3577 (
            .O(N__16661),
            .I(N__16658));
    CascadeMux I__3576 (
            .O(N__16658),
            .I(N__16655));
    CascadeBuf I__3575 (
            .O(N__16655),
            .I(N__16652));
    CascadeMux I__3574 (
            .O(N__16652),
            .I(N__16649));
    CascadeBuf I__3573 (
            .O(N__16649),
            .I(N__16646));
    CascadeMux I__3572 (
            .O(N__16646),
            .I(N__16643));
    CascadeBuf I__3571 (
            .O(N__16643),
            .I(N__16640));
    CascadeMux I__3570 (
            .O(N__16640),
            .I(N__16637));
    CascadeBuf I__3569 (
            .O(N__16637),
            .I(N__16634));
    CascadeMux I__3568 (
            .O(N__16634),
            .I(N__16631));
    CascadeBuf I__3567 (
            .O(N__16631),
            .I(N__16628));
    CascadeMux I__3566 (
            .O(N__16628),
            .I(N__16625));
    CascadeBuf I__3565 (
            .O(N__16625),
            .I(N__16622));
    CascadeMux I__3564 (
            .O(N__16622),
            .I(N__16619));
    CascadeBuf I__3563 (
            .O(N__16619),
            .I(N__16616));
    CascadeMux I__3562 (
            .O(N__16616),
            .I(N__16613));
    CascadeBuf I__3561 (
            .O(N__16613),
            .I(N__16610));
    CascadeMux I__3560 (
            .O(N__16610),
            .I(N__16607));
    CascadeBuf I__3559 (
            .O(N__16607),
            .I(N__16604));
    CascadeMux I__3558 (
            .O(N__16604),
            .I(N__16601));
    CascadeBuf I__3557 (
            .O(N__16601),
            .I(N__16598));
    CascadeMux I__3556 (
            .O(N__16598),
            .I(N__16595));
    CascadeBuf I__3555 (
            .O(N__16595),
            .I(N__16592));
    CascadeMux I__3554 (
            .O(N__16592),
            .I(N__16589));
    CascadeBuf I__3553 (
            .O(N__16589),
            .I(N__16586));
    CascadeMux I__3552 (
            .O(N__16586),
            .I(N__16583));
    CascadeBuf I__3551 (
            .O(N__16583),
            .I(N__16580));
    CascadeMux I__3550 (
            .O(N__16580),
            .I(N__16577));
    CascadeBuf I__3549 (
            .O(N__16577),
            .I(N__16574));
    CascadeMux I__3548 (
            .O(N__16574),
            .I(N__16571));
    InMux I__3547 (
            .O(N__16571),
            .I(N__16568));
    LocalMux I__3546 (
            .O(N__16568),
            .I(N__16565));
    Span12Mux_s3_v I__3545 (
            .O(N__16565),
            .I(N__16562));
    Span12Mux_v I__3544 (
            .O(N__16562),
            .I(N__16559));
    Odrv12 I__3543 (
            .O(N__16559),
            .I(M_this_ppu_sprites_addr_1));
    InMux I__3542 (
            .O(N__16556),
            .I(N__16553));
    LocalMux I__3541 (
            .O(N__16553),
            .I(M_this_sprites_address_q_3_ns_1_10));
    InMux I__3540 (
            .O(N__16550),
            .I(N__16547));
    LocalMux I__3539 (
            .O(N__16547),
            .I(N__16544));
    Odrv12 I__3538 (
            .O(N__16544),
            .I(M_this_sprites_address_q_RNO_1Z0Z_10));
    CascadeMux I__3537 (
            .O(N__16541),
            .I(N__16538));
    CascadeBuf I__3536 (
            .O(N__16538),
            .I(N__16535));
    CascadeMux I__3535 (
            .O(N__16535),
            .I(N__16532));
    CascadeBuf I__3534 (
            .O(N__16532),
            .I(N__16529));
    CascadeMux I__3533 (
            .O(N__16529),
            .I(N__16526));
    CascadeBuf I__3532 (
            .O(N__16526),
            .I(N__16523));
    CascadeMux I__3531 (
            .O(N__16523),
            .I(N__16520));
    CascadeBuf I__3530 (
            .O(N__16520),
            .I(N__16517));
    CascadeMux I__3529 (
            .O(N__16517),
            .I(N__16514));
    CascadeBuf I__3528 (
            .O(N__16514),
            .I(N__16511));
    CascadeMux I__3527 (
            .O(N__16511),
            .I(N__16508));
    CascadeBuf I__3526 (
            .O(N__16508),
            .I(N__16505));
    CascadeMux I__3525 (
            .O(N__16505),
            .I(N__16502));
    CascadeBuf I__3524 (
            .O(N__16502),
            .I(N__16499));
    CascadeMux I__3523 (
            .O(N__16499),
            .I(N__16496));
    CascadeBuf I__3522 (
            .O(N__16496),
            .I(N__16493));
    CascadeMux I__3521 (
            .O(N__16493),
            .I(N__16490));
    CascadeBuf I__3520 (
            .O(N__16490),
            .I(N__16487));
    CascadeMux I__3519 (
            .O(N__16487),
            .I(N__16484));
    CascadeBuf I__3518 (
            .O(N__16484),
            .I(N__16481));
    CascadeMux I__3517 (
            .O(N__16481),
            .I(N__16478));
    CascadeBuf I__3516 (
            .O(N__16478),
            .I(N__16475));
    CascadeMux I__3515 (
            .O(N__16475),
            .I(N__16472));
    CascadeBuf I__3514 (
            .O(N__16472),
            .I(N__16469));
    CascadeMux I__3513 (
            .O(N__16469),
            .I(N__16466));
    CascadeBuf I__3512 (
            .O(N__16466),
            .I(N__16463));
    CascadeMux I__3511 (
            .O(N__16463),
            .I(N__16460));
    CascadeBuf I__3510 (
            .O(N__16460),
            .I(N__16457));
    CascadeMux I__3509 (
            .O(N__16457),
            .I(N__16454));
    CascadeBuf I__3508 (
            .O(N__16454),
            .I(N__16451));
    CascadeMux I__3507 (
            .O(N__16451),
            .I(N__16448));
    InMux I__3506 (
            .O(N__16448),
            .I(N__16445));
    LocalMux I__3505 (
            .O(N__16445),
            .I(N__16441));
    InMux I__3504 (
            .O(N__16444),
            .I(N__16438));
    Sp12to4 I__3503 (
            .O(N__16441),
            .I(N__16434));
    LocalMux I__3502 (
            .O(N__16438),
            .I(N__16431));
    InMux I__3501 (
            .O(N__16437),
            .I(N__16428));
    Span12Mux_h I__3500 (
            .O(N__16434),
            .I(N__16425));
    Odrv12 I__3499 (
            .O(N__16431),
            .I(M_this_sprites_address_qZ0Z_10));
    LocalMux I__3498 (
            .O(N__16428),
            .I(M_this_sprites_address_qZ0Z_10));
    Odrv12 I__3497 (
            .O(N__16425),
            .I(M_this_sprites_address_qZ0Z_10));
    InMux I__3496 (
            .O(N__16418),
            .I(N__16405));
    InMux I__3495 (
            .O(N__16417),
            .I(N__16405));
    InMux I__3494 (
            .O(N__16416),
            .I(N__16401));
    InMux I__3493 (
            .O(N__16415),
            .I(N__16397));
    InMux I__3492 (
            .O(N__16414),
            .I(N__16393));
    InMux I__3491 (
            .O(N__16413),
            .I(N__16390));
    InMux I__3490 (
            .O(N__16412),
            .I(N__16387));
    InMux I__3489 (
            .O(N__16411),
            .I(N__16382));
    InMux I__3488 (
            .O(N__16410),
            .I(N__16379));
    LocalMux I__3487 (
            .O(N__16405),
            .I(N__16376));
    CascadeMux I__3486 (
            .O(N__16404),
            .I(N__16372));
    LocalMux I__3485 (
            .O(N__16401),
            .I(N__16368));
    InMux I__3484 (
            .O(N__16400),
            .I(N__16365));
    LocalMux I__3483 (
            .O(N__16397),
            .I(N__16362));
    InMux I__3482 (
            .O(N__16396),
            .I(N__16359));
    LocalMux I__3481 (
            .O(N__16393),
            .I(N__16354));
    LocalMux I__3480 (
            .O(N__16390),
            .I(N__16354));
    LocalMux I__3479 (
            .O(N__16387),
            .I(N__16351));
    InMux I__3478 (
            .O(N__16386),
            .I(N__16348));
    InMux I__3477 (
            .O(N__16385),
            .I(N__16345));
    LocalMux I__3476 (
            .O(N__16382),
            .I(N__16338));
    LocalMux I__3475 (
            .O(N__16379),
            .I(N__16338));
    Span4Mux_v I__3474 (
            .O(N__16376),
            .I(N__16338));
    InMux I__3473 (
            .O(N__16375),
            .I(N__16335));
    InMux I__3472 (
            .O(N__16372),
            .I(N__16332));
    InMux I__3471 (
            .O(N__16371),
            .I(N__16329));
    Span4Mux_v I__3470 (
            .O(N__16368),
            .I(N__16324));
    LocalMux I__3469 (
            .O(N__16365),
            .I(N__16324));
    Span4Mux_v I__3468 (
            .O(N__16362),
            .I(N__16313));
    LocalMux I__3467 (
            .O(N__16359),
            .I(N__16313));
    Span4Mux_v I__3466 (
            .O(N__16354),
            .I(N__16313));
    Span4Mux_v I__3465 (
            .O(N__16351),
            .I(N__16313));
    LocalMux I__3464 (
            .O(N__16348),
            .I(N__16313));
    LocalMux I__3463 (
            .O(N__16345),
            .I(N__16310));
    Span4Mux_h I__3462 (
            .O(N__16338),
            .I(N__16305));
    LocalMux I__3461 (
            .O(N__16335),
            .I(N__16305));
    LocalMux I__3460 (
            .O(N__16332),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__3459 (
            .O(N__16329),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3458 (
            .O(N__16324),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3457 (
            .O(N__16313),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3456 (
            .O(N__16310),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3455 (
            .O(N__16305),
            .I(M_this_state_qZ0Z_5));
    InMux I__3454 (
            .O(N__16292),
            .I(N__16289));
    LocalMux I__3453 (
            .O(N__16289),
            .I(N_202));
    InMux I__3452 (
            .O(N__16286),
            .I(N__16280));
    InMux I__3451 (
            .O(N__16285),
            .I(N__16280));
    LocalMux I__3450 (
            .O(N__16280),
            .I(M_this_state_qZ0Z_6));
    InMux I__3449 (
            .O(N__16277),
            .I(N__16272));
    InMux I__3448 (
            .O(N__16276),
            .I(N__16269));
    InMux I__3447 (
            .O(N__16275),
            .I(N__16266));
    LocalMux I__3446 (
            .O(N__16272),
            .I(N__16263));
    LocalMux I__3445 (
            .O(N__16269),
            .I(N_233));
    LocalMux I__3444 (
            .O(N__16266),
            .I(N_233));
    Odrv4 I__3443 (
            .O(N__16263),
            .I(N_233));
    InMux I__3442 (
            .O(N__16256),
            .I(N__16253));
    LocalMux I__3441 (
            .O(N__16253),
            .I(N__16250));
    Span4Mux_h I__3440 (
            .O(N__16250),
            .I(N__16244));
    CascadeMux I__3439 (
            .O(N__16249),
            .I(N__16241));
    InMux I__3438 (
            .O(N__16248),
            .I(N__16236));
    InMux I__3437 (
            .O(N__16247),
            .I(N__16236));
    Span4Mux_h I__3436 (
            .O(N__16244),
            .I(N__16233));
    InMux I__3435 (
            .O(N__16241),
            .I(N__16230));
    LocalMux I__3434 (
            .O(N__16236),
            .I(N__16227));
    Odrv4 I__3433 (
            .O(N__16233),
            .I(M_this_start_address_delay_out_0));
    LocalMux I__3432 (
            .O(N__16230),
            .I(M_this_start_address_delay_out_0));
    Odrv4 I__3431 (
            .O(N__16227),
            .I(M_this_start_address_delay_out_0));
    CascadeMux I__3430 (
            .O(N__16220),
            .I(M_this_state_q_srsts_i_1_1_cascade_));
    InMux I__3429 (
            .O(N__16217),
            .I(N__16210));
    InMux I__3428 (
            .O(N__16216),
            .I(N__16205));
    InMux I__3427 (
            .O(N__16215),
            .I(N__16205));
    InMux I__3426 (
            .O(N__16214),
            .I(N__16201));
    InMux I__3425 (
            .O(N__16213),
            .I(N__16198));
    LocalMux I__3424 (
            .O(N__16210),
            .I(N__16193));
    LocalMux I__3423 (
            .O(N__16205),
            .I(N__16193));
    InMux I__3422 (
            .O(N__16204),
            .I(N__16190));
    LocalMux I__3421 (
            .O(N__16201),
            .I(N__16185));
    LocalMux I__3420 (
            .O(N__16198),
            .I(N__16185));
    Span4Mux_h I__3419 (
            .O(N__16193),
            .I(N__16182));
    LocalMux I__3418 (
            .O(N__16190),
            .I(M_this_state_qZ0Z_1));
    Odrv12 I__3417 (
            .O(N__16185),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__3416 (
            .O(N__16182),
            .I(M_this_state_qZ0Z_1));
    CascadeMux I__3415 (
            .O(N__16175),
            .I(N__16171));
    InMux I__3414 (
            .O(N__16174),
            .I(N__16167));
    InMux I__3413 (
            .O(N__16171),
            .I(N__16162));
    InMux I__3412 (
            .O(N__16170),
            .I(N__16162));
    LocalMux I__3411 (
            .O(N__16167),
            .I(N__16153));
    LocalMux I__3410 (
            .O(N__16162),
            .I(N__16153));
    InMux I__3409 (
            .O(N__16161),
            .I(N__16144));
    InMux I__3408 (
            .O(N__16160),
            .I(N__16144));
    InMux I__3407 (
            .O(N__16159),
            .I(N__16144));
    InMux I__3406 (
            .O(N__16158),
            .I(N__16144));
    Span4Mux_h I__3405 (
            .O(N__16153),
            .I(N__16141));
    LocalMux I__3404 (
            .O(N__16144),
            .I(N__16138));
    Odrv4 I__3403 (
            .O(N__16141),
            .I(\this_ppu.N_250_1 ));
    Odrv4 I__3402 (
            .O(N__16138),
            .I(\this_ppu.N_250_1 ));
    InMux I__3401 (
            .O(N__16133),
            .I(N__16124));
    InMux I__3400 (
            .O(N__16132),
            .I(N__16124));
    InMux I__3399 (
            .O(N__16131),
            .I(N__16124));
    LocalMux I__3398 (
            .O(N__16124),
            .I(N__16121));
    Span4Mux_h I__3397 (
            .O(N__16121),
            .I(N__16116));
    InMux I__3396 (
            .O(N__16120),
            .I(N__16113));
    InMux I__3395 (
            .O(N__16119),
            .I(N__16110));
    Odrv4 I__3394 (
            .O(N__16116),
            .I(\this_ppu.M_last_q_RNI5NOQ4 ));
    LocalMux I__3393 (
            .O(N__16113),
            .I(\this_ppu.M_last_q_RNI5NOQ4 ));
    LocalMux I__3392 (
            .O(N__16110),
            .I(\this_ppu.M_last_q_RNI5NOQ4 ));
    InMux I__3391 (
            .O(N__16103),
            .I(N__16098));
    InMux I__3390 (
            .O(N__16102),
            .I(N__16093));
    InMux I__3389 (
            .O(N__16101),
            .I(N__16093));
    LocalMux I__3388 (
            .O(N__16098),
            .I(\this_ppu.un1_M_vaddress_q_c3 ));
    LocalMux I__3387 (
            .O(N__16093),
            .I(\this_ppu.un1_M_vaddress_q_c3 ));
    InMux I__3386 (
            .O(N__16088),
            .I(N__16085));
    LocalMux I__3385 (
            .O(N__16085),
            .I(\this_ppu.un1_M_haddress_q_c5 ));
    InMux I__3384 (
            .O(N__16082),
            .I(N__16076));
    InMux I__3383 (
            .O(N__16081),
            .I(N__16076));
    LocalMux I__3382 (
            .O(N__16076),
            .I(\this_ppu.un1_M_haddress_q_c2 ));
    InMux I__3381 (
            .O(N__16073),
            .I(N__16068));
    InMux I__3380 (
            .O(N__16072),
            .I(N__16065));
    InMux I__3379 (
            .O(N__16071),
            .I(N__16062));
    LocalMux I__3378 (
            .O(N__16068),
            .I(\this_ppu.un1_M_vaddress_q_c1 ));
    LocalMux I__3377 (
            .O(N__16065),
            .I(\this_ppu.un1_M_vaddress_q_c1 ));
    LocalMux I__3376 (
            .O(N__16062),
            .I(\this_ppu.un1_M_vaddress_q_c1 ));
    InMux I__3375 (
            .O(N__16055),
            .I(N__16046));
    InMux I__3374 (
            .O(N__16054),
            .I(N__16046));
    InMux I__3373 (
            .O(N__16053),
            .I(N__16046));
    LocalMux I__3372 (
            .O(N__16046),
            .I(N__16042));
    InMux I__3371 (
            .O(N__16045),
            .I(N__16039));
    Span4Mux_v I__3370 (
            .O(N__16042),
            .I(N__16036));
    LocalMux I__3369 (
            .O(N__16039),
            .I(N__16033));
    Span4Mux_v I__3368 (
            .O(N__16036),
            .I(N__16030));
    Sp12to4 I__3367 (
            .O(N__16033),
            .I(N__16027));
    IoSpan4Mux I__3366 (
            .O(N__16030),
            .I(N__16024));
    Odrv12 I__3365 (
            .O(N__16027),
            .I(port_address_in_0));
    Odrv4 I__3364 (
            .O(N__16024),
            .I(port_address_in_0));
    InMux I__3363 (
            .O(N__16019),
            .I(N__16013));
    InMux I__3362 (
            .O(N__16018),
            .I(N__16006));
    InMux I__3361 (
            .O(N__16017),
            .I(N__16006));
    InMux I__3360 (
            .O(N__16016),
            .I(N__16006));
    LocalMux I__3359 (
            .O(N__16013),
            .I(N__16003));
    LocalMux I__3358 (
            .O(N__16006),
            .I(N__16000));
    Span4Mux_v I__3357 (
            .O(N__16003),
            .I(N__15997));
    Span4Mux_v I__3356 (
            .O(N__16000),
            .I(N__15994));
    Sp12to4 I__3355 (
            .O(N__15997),
            .I(N__15991));
    Sp12to4 I__3354 (
            .O(N__15994),
            .I(N__15988));
    Span12Mux_h I__3353 (
            .O(N__15991),
            .I(N__15985));
    Span12Mux_h I__3352 (
            .O(N__15988),
            .I(N__15982));
    Odrv12 I__3351 (
            .O(N__15985),
            .I(port_address_in_1));
    Odrv12 I__3350 (
            .O(N__15982),
            .I(port_address_in_1));
    InMux I__3349 (
            .O(N__15977),
            .I(N__15968));
    InMux I__3348 (
            .O(N__15976),
            .I(N__15968));
    InMux I__3347 (
            .O(N__15975),
            .I(N__15968));
    LocalMux I__3346 (
            .O(N__15968),
            .I(N__15965));
    Odrv4 I__3345 (
            .O(N__15965),
            .I(N_218));
    InMux I__3344 (
            .O(N__15962),
            .I(N__15959));
    LocalMux I__3343 (
            .O(N__15959),
            .I(N_204));
    CascadeMux I__3342 (
            .O(N__15956),
            .I(N__15952));
    CascadeMux I__3341 (
            .O(N__15955),
            .I(N__15949));
    InMux I__3340 (
            .O(N__15952),
            .I(N__15946));
    InMux I__3339 (
            .O(N__15949),
            .I(N__15943));
    LocalMux I__3338 (
            .O(N__15946),
            .I(N__15940));
    LocalMux I__3337 (
            .O(N__15943),
            .I(M_this_data_count_qZ0Z_12));
    Odrv4 I__3336 (
            .O(N__15940),
            .I(M_this_data_count_qZ0Z_12));
    InMux I__3335 (
            .O(N__15935),
            .I(un1_M_this_data_count_q_cry_11));
    SRMux I__3334 (
            .O(N__15932),
            .I(N__15929));
    LocalMux I__3333 (
            .O(N__15929),
            .I(N__15926));
    Span4Mux_v I__3332 (
            .O(N__15926),
            .I(N__15922));
    SRMux I__3331 (
            .O(N__15925),
            .I(N__15919));
    Span4Mux_h I__3330 (
            .O(N__15922),
            .I(N__15916));
    LocalMux I__3329 (
            .O(N__15919),
            .I(N__15913));
    Odrv4 I__3328 (
            .O(N__15916),
            .I(M_this_state_q_RNI20CEZ0Z_0));
    Odrv12 I__3327 (
            .O(N__15913),
            .I(M_this_state_q_RNI20CEZ0Z_0));
    SRMux I__3326 (
            .O(N__15908),
            .I(N__15899));
    SRMux I__3325 (
            .O(N__15907),
            .I(N__15896));
    SRMux I__3324 (
            .O(N__15906),
            .I(N__15893));
    SRMux I__3323 (
            .O(N__15905),
            .I(N__15890));
    SRMux I__3322 (
            .O(N__15904),
            .I(N__15884));
    SRMux I__3321 (
            .O(N__15903),
            .I(N__15877));
    SRMux I__3320 (
            .O(N__15902),
            .I(N__15872));
    LocalMux I__3319 (
            .O(N__15899),
            .I(N__15869));
    LocalMux I__3318 (
            .O(N__15896),
            .I(N__15866));
    LocalMux I__3317 (
            .O(N__15893),
            .I(N__15861));
    LocalMux I__3316 (
            .O(N__15890),
            .I(N__15861));
    SRMux I__3315 (
            .O(N__15889),
            .I(N__15858));
    SRMux I__3314 (
            .O(N__15888),
            .I(N__15855));
    SRMux I__3313 (
            .O(N__15887),
            .I(N__15850));
    LocalMux I__3312 (
            .O(N__15884),
            .I(N__15845));
    SRMux I__3311 (
            .O(N__15883),
            .I(N__15842));
    SRMux I__3310 (
            .O(N__15882),
            .I(N__15837));
    SRMux I__3309 (
            .O(N__15881),
            .I(N__15834));
    SRMux I__3308 (
            .O(N__15880),
            .I(N__15831));
    LocalMux I__3307 (
            .O(N__15877),
            .I(N__15826));
    SRMux I__3306 (
            .O(N__15876),
            .I(N__15823));
    SRMux I__3305 (
            .O(N__15875),
            .I(N__15820));
    LocalMux I__3304 (
            .O(N__15872),
            .I(N__15817));
    Span4Mux_s3_v I__3303 (
            .O(N__15869),
            .I(N__15806));
    Span4Mux_h I__3302 (
            .O(N__15866),
            .I(N__15806));
    Span4Mux_s3_v I__3301 (
            .O(N__15861),
            .I(N__15806));
    LocalMux I__3300 (
            .O(N__15858),
            .I(N__15806));
    LocalMux I__3299 (
            .O(N__15855),
            .I(N__15806));
    SRMux I__3298 (
            .O(N__15854),
            .I(N__15803));
    SRMux I__3297 (
            .O(N__15853),
            .I(N__15800));
    LocalMux I__3296 (
            .O(N__15850),
            .I(N__15794));
    SRMux I__3295 (
            .O(N__15849),
            .I(N__15791));
    SRMux I__3294 (
            .O(N__15848),
            .I(N__15787));
    Span4Mux_h I__3293 (
            .O(N__15845),
            .I(N__15781));
    LocalMux I__3292 (
            .O(N__15842),
            .I(N__15781));
    SRMux I__3291 (
            .O(N__15841),
            .I(N__15778));
    SRMux I__3290 (
            .O(N__15840),
            .I(N__15775));
    LocalMux I__3289 (
            .O(N__15837),
            .I(N__15769));
    LocalMux I__3288 (
            .O(N__15834),
            .I(N__15769));
    LocalMux I__3287 (
            .O(N__15831),
            .I(N__15766));
    SRMux I__3286 (
            .O(N__15830),
            .I(N__15763));
    SRMux I__3285 (
            .O(N__15829),
            .I(N__15760));
    Span4Mux_v I__3284 (
            .O(N__15826),
            .I(N__15753));
    LocalMux I__3283 (
            .O(N__15823),
            .I(N__15753));
    LocalMux I__3282 (
            .O(N__15820),
            .I(N__15750));
    Span4Mux_h I__3281 (
            .O(N__15817),
            .I(N__15741));
    Span4Mux_v I__3280 (
            .O(N__15806),
            .I(N__15741));
    LocalMux I__3279 (
            .O(N__15803),
            .I(N__15741));
    LocalMux I__3278 (
            .O(N__15800),
            .I(N__15741));
    SRMux I__3277 (
            .O(N__15799),
            .I(N__15738));
    SRMux I__3276 (
            .O(N__15798),
            .I(N__15735));
    IoInMux I__3275 (
            .O(N__15797),
            .I(N__15730));
    Span4Mux_v I__3274 (
            .O(N__15794),
            .I(N__15727));
    LocalMux I__3273 (
            .O(N__15791),
            .I(N__15724));
    SRMux I__3272 (
            .O(N__15790),
            .I(N__15721));
    LocalMux I__3271 (
            .O(N__15787),
            .I(N__15718));
    SRMux I__3270 (
            .O(N__15786),
            .I(N__15715));
    Span4Mux_v I__3269 (
            .O(N__15781),
            .I(N__15710));
    LocalMux I__3268 (
            .O(N__15778),
            .I(N__15710));
    LocalMux I__3267 (
            .O(N__15775),
            .I(N__15707));
    SRMux I__3266 (
            .O(N__15774),
            .I(N__15704));
    Span4Mux_v I__3265 (
            .O(N__15769),
            .I(N__15695));
    Span4Mux_h I__3264 (
            .O(N__15766),
            .I(N__15695));
    LocalMux I__3263 (
            .O(N__15763),
            .I(N__15695));
    LocalMux I__3262 (
            .O(N__15760),
            .I(N__15695));
    SRMux I__3261 (
            .O(N__15759),
            .I(N__15692));
    SRMux I__3260 (
            .O(N__15758),
            .I(N__15689));
    Span4Mux_v I__3259 (
            .O(N__15753),
            .I(N__15677));
    Span4Mux_h I__3258 (
            .O(N__15750),
            .I(N__15677));
    Span4Mux_v I__3257 (
            .O(N__15741),
            .I(N__15677));
    LocalMux I__3256 (
            .O(N__15738),
            .I(N__15677));
    LocalMux I__3255 (
            .O(N__15735),
            .I(N__15677));
    SRMux I__3254 (
            .O(N__15734),
            .I(N__15674));
    SRMux I__3253 (
            .O(N__15733),
            .I(N__15671));
    LocalMux I__3252 (
            .O(N__15730),
            .I(N__15665));
    Span4Mux_h I__3251 (
            .O(N__15727),
            .I(N__15660));
    Span4Mux_v I__3250 (
            .O(N__15724),
            .I(N__15660));
    LocalMux I__3249 (
            .O(N__15721),
            .I(N__15657));
    Span4Mux_v I__3248 (
            .O(N__15718),
            .I(N__15652));
    LocalMux I__3247 (
            .O(N__15715),
            .I(N__15652));
    Span4Mux_v I__3246 (
            .O(N__15710),
            .I(N__15645));
    Span4Mux_h I__3245 (
            .O(N__15707),
            .I(N__15645));
    LocalMux I__3244 (
            .O(N__15704),
            .I(N__15645));
    Span4Mux_v I__3243 (
            .O(N__15695),
            .I(N__15638));
    LocalMux I__3242 (
            .O(N__15692),
            .I(N__15638));
    LocalMux I__3241 (
            .O(N__15689),
            .I(N__15638));
    SRMux I__3240 (
            .O(N__15688),
            .I(N__15635));
    Span4Mux_v I__3239 (
            .O(N__15677),
            .I(N__15628));
    LocalMux I__3238 (
            .O(N__15674),
            .I(N__15628));
    LocalMux I__3237 (
            .O(N__15671),
            .I(N__15628));
    InMux I__3236 (
            .O(N__15670),
            .I(N__15625));
    InMux I__3235 (
            .O(N__15669),
            .I(N__15620));
    InMux I__3234 (
            .O(N__15668),
            .I(N__15620));
    Span4Mux_s1_h I__3233 (
            .O(N__15665),
            .I(N__15617));
    Sp12to4 I__3232 (
            .O(N__15660),
            .I(N__15614));
    Span4Mux_h I__3231 (
            .O(N__15657),
            .I(N__15611));
    Span4Mux_v I__3230 (
            .O(N__15652),
            .I(N__15606));
    Span4Mux_v I__3229 (
            .O(N__15645),
            .I(N__15606));
    Span4Mux_v I__3228 (
            .O(N__15638),
            .I(N__15599));
    LocalMux I__3227 (
            .O(N__15635),
            .I(N__15599));
    Span4Mux_v I__3226 (
            .O(N__15628),
            .I(N__15599));
    LocalMux I__3225 (
            .O(N__15625),
            .I(N__15594));
    LocalMux I__3224 (
            .O(N__15620),
            .I(N__15594));
    Sp12to4 I__3223 (
            .O(N__15617),
            .I(N__15591));
    Span12Mux_s9_h I__3222 (
            .O(N__15614),
            .I(N__15588));
    Span4Mux_v I__3221 (
            .O(N__15611),
            .I(N__15581));
    Span4Mux_h I__3220 (
            .O(N__15606),
            .I(N__15581));
    Span4Mux_h I__3219 (
            .O(N__15599),
            .I(N__15581));
    Span4Mux_h I__3218 (
            .O(N__15594),
            .I(N__15578));
    Span12Mux_v I__3217 (
            .O(N__15591),
            .I(N__15575));
    Span12Mux_v I__3216 (
            .O(N__15588),
            .I(N__15570));
    Sp12to4 I__3215 (
            .O(N__15581),
            .I(N__15570));
    Span4Mux_v I__3214 (
            .O(N__15578),
            .I(N__15567));
    Odrv12 I__3213 (
            .O(N__15575),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3212 (
            .O(N__15570),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3211 (
            .O(N__15567),
            .I(CONSTANT_ONE_NET));
    InMux I__3210 (
            .O(N__15560),
            .I(bfn_17_25_0_));
    InMux I__3209 (
            .O(N__15557),
            .I(N__15553));
    InMux I__3208 (
            .O(N__15556),
            .I(N__15550));
    LocalMux I__3207 (
            .O(N__15553),
            .I(N__15547));
    LocalMux I__3206 (
            .O(N__15550),
            .I(M_this_data_count_qZ0Z_13));
    Odrv4 I__3205 (
            .O(N__15547),
            .I(M_this_data_count_qZ0Z_13));
    CascadeMux I__3204 (
            .O(N__15542),
            .I(\this_ppu.un1_M_haddress_q_c2_cascade_ ));
    CascadeMux I__3203 (
            .O(N__15539),
            .I(\this_ppu.un1_M_haddress_q_c5_cascade_ ));
    CascadeMux I__3202 (
            .O(N__15536),
            .I(N__15532));
    CascadeMux I__3201 (
            .O(N__15535),
            .I(N__15529));
    InMux I__3200 (
            .O(N__15532),
            .I(N__15526));
    InMux I__3199 (
            .O(N__15529),
            .I(N__15523));
    LocalMux I__3198 (
            .O(N__15526),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__3197 (
            .O(N__15523),
            .I(M_this_data_count_qZ0Z_4));
    InMux I__3196 (
            .O(N__15518),
            .I(un1_M_this_data_count_q_cry_3));
    CascadeMux I__3195 (
            .O(N__15515),
            .I(N__15512));
    InMux I__3194 (
            .O(N__15512),
            .I(N__15508));
    InMux I__3193 (
            .O(N__15511),
            .I(N__15505));
    LocalMux I__3192 (
            .O(N__15508),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__3191 (
            .O(N__15505),
            .I(M_this_data_count_qZ0Z_5));
    InMux I__3190 (
            .O(N__15500),
            .I(un1_M_this_data_count_q_cry_4));
    CascadeMux I__3189 (
            .O(N__15497),
            .I(N__15494));
    InMux I__3188 (
            .O(N__15494),
            .I(N__15490));
    InMux I__3187 (
            .O(N__15493),
            .I(N__15487));
    LocalMux I__3186 (
            .O(N__15490),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__3185 (
            .O(N__15487),
            .I(M_this_data_count_qZ0Z_6));
    InMux I__3184 (
            .O(N__15482),
            .I(un1_M_this_data_count_q_cry_5));
    CascadeMux I__3183 (
            .O(N__15479),
            .I(N__15476));
    InMux I__3182 (
            .O(N__15476),
            .I(N__15472));
    InMux I__3181 (
            .O(N__15475),
            .I(N__15469));
    LocalMux I__3180 (
            .O(N__15472),
            .I(M_this_data_count_qZ0Z_7));
    LocalMux I__3179 (
            .O(N__15469),
            .I(M_this_data_count_qZ0Z_7));
    InMux I__3178 (
            .O(N__15464),
            .I(un1_M_this_data_count_q_cry_6));
    CascadeMux I__3177 (
            .O(N__15461),
            .I(N__15457));
    InMux I__3176 (
            .O(N__15460),
            .I(N__15454));
    InMux I__3175 (
            .O(N__15457),
            .I(N__15451));
    LocalMux I__3174 (
            .O(N__15454),
            .I(N__15448));
    LocalMux I__3173 (
            .O(N__15451),
            .I(M_this_data_count_qZ0Z_8));
    Odrv4 I__3172 (
            .O(N__15448),
            .I(M_this_data_count_qZ0Z_8));
    InMux I__3171 (
            .O(N__15443),
            .I(bfn_17_24_0_));
    CascadeMux I__3170 (
            .O(N__15440),
            .I(N__15436));
    InMux I__3169 (
            .O(N__15439),
            .I(N__15433));
    InMux I__3168 (
            .O(N__15436),
            .I(N__15430));
    LocalMux I__3167 (
            .O(N__15433),
            .I(N__15427));
    LocalMux I__3166 (
            .O(N__15430),
            .I(M_this_data_count_qZ0Z_9));
    Odrv4 I__3165 (
            .O(N__15427),
            .I(M_this_data_count_qZ0Z_9));
    InMux I__3164 (
            .O(N__15422),
            .I(un1_M_this_data_count_q_cry_8));
    CascadeMux I__3163 (
            .O(N__15419),
            .I(N__15415));
    CascadeMux I__3162 (
            .O(N__15418),
            .I(N__15412));
    InMux I__3161 (
            .O(N__15415),
            .I(N__15409));
    InMux I__3160 (
            .O(N__15412),
            .I(N__15406));
    LocalMux I__3159 (
            .O(N__15409),
            .I(N__15403));
    LocalMux I__3158 (
            .O(N__15406),
            .I(M_this_data_count_qZ0Z_10));
    Odrv4 I__3157 (
            .O(N__15403),
            .I(M_this_data_count_qZ0Z_10));
    InMux I__3156 (
            .O(N__15398),
            .I(un1_M_this_data_count_q_cry_9));
    CascadeMux I__3155 (
            .O(N__15395),
            .I(N__15391));
    InMux I__3154 (
            .O(N__15394),
            .I(N__15388));
    InMux I__3153 (
            .O(N__15391),
            .I(N__15385));
    LocalMux I__3152 (
            .O(N__15388),
            .I(N__15382));
    LocalMux I__3151 (
            .O(N__15385),
            .I(M_this_data_count_qZ0Z_11));
    Odrv4 I__3150 (
            .O(N__15382),
            .I(M_this_data_count_qZ0Z_11));
    InMux I__3149 (
            .O(N__15377),
            .I(un1_M_this_data_count_q_cry_10));
    CascadeMux I__3148 (
            .O(N__15374),
            .I(N__15371));
    CascadeBuf I__3147 (
            .O(N__15371),
            .I(N__15368));
    CascadeMux I__3146 (
            .O(N__15368),
            .I(N__15365));
    CascadeBuf I__3145 (
            .O(N__15365),
            .I(N__15362));
    CascadeMux I__3144 (
            .O(N__15362),
            .I(N__15359));
    CascadeBuf I__3143 (
            .O(N__15359),
            .I(N__15356));
    CascadeMux I__3142 (
            .O(N__15356),
            .I(N__15353));
    CascadeBuf I__3141 (
            .O(N__15353),
            .I(N__15350));
    CascadeMux I__3140 (
            .O(N__15350),
            .I(N__15347));
    CascadeBuf I__3139 (
            .O(N__15347),
            .I(N__15344));
    CascadeMux I__3138 (
            .O(N__15344),
            .I(N__15341));
    CascadeBuf I__3137 (
            .O(N__15341),
            .I(N__15338));
    CascadeMux I__3136 (
            .O(N__15338),
            .I(N__15335));
    CascadeBuf I__3135 (
            .O(N__15335),
            .I(N__15332));
    CascadeMux I__3134 (
            .O(N__15332),
            .I(N__15329));
    CascadeBuf I__3133 (
            .O(N__15329),
            .I(N__15326));
    CascadeMux I__3132 (
            .O(N__15326),
            .I(N__15323));
    CascadeBuf I__3131 (
            .O(N__15323),
            .I(N__15320));
    CascadeMux I__3130 (
            .O(N__15320),
            .I(N__15317));
    CascadeBuf I__3129 (
            .O(N__15317),
            .I(N__15314));
    CascadeMux I__3128 (
            .O(N__15314),
            .I(N__15311));
    CascadeBuf I__3127 (
            .O(N__15311),
            .I(N__15308));
    CascadeMux I__3126 (
            .O(N__15308),
            .I(N__15305));
    CascadeBuf I__3125 (
            .O(N__15305),
            .I(N__15302));
    CascadeMux I__3124 (
            .O(N__15302),
            .I(N__15299));
    CascadeBuf I__3123 (
            .O(N__15299),
            .I(N__15296));
    CascadeMux I__3122 (
            .O(N__15296),
            .I(N__15293));
    CascadeBuf I__3121 (
            .O(N__15293),
            .I(N__15290));
    CascadeMux I__3120 (
            .O(N__15290),
            .I(N__15287));
    CascadeBuf I__3119 (
            .O(N__15287),
            .I(N__15284));
    CascadeMux I__3118 (
            .O(N__15284),
            .I(N__15280));
    InMux I__3117 (
            .O(N__15283),
            .I(N__15277));
    InMux I__3116 (
            .O(N__15280),
            .I(N__15274));
    LocalMux I__3115 (
            .O(N__15277),
            .I(N__15271));
    LocalMux I__3114 (
            .O(N__15274),
            .I(N__15267));
    Span4Mux_h I__3113 (
            .O(N__15271),
            .I(N__15264));
    InMux I__3112 (
            .O(N__15270),
            .I(N__15261));
    Span12Mux_s11_v I__3111 (
            .O(N__15267),
            .I(N__15258));
    Odrv4 I__3110 (
            .O(N__15264),
            .I(M_this_sprites_address_qZ0Z_0));
    LocalMux I__3109 (
            .O(N__15261),
            .I(M_this_sprites_address_qZ0Z_0));
    Odrv12 I__3108 (
            .O(N__15258),
            .I(M_this_sprites_address_qZ0Z_0));
    InMux I__3107 (
            .O(N__15251),
            .I(N__15248));
    LocalMux I__3106 (
            .O(N__15248),
            .I(M_this_sprites_address_q_3_ns_1_0));
    InMux I__3105 (
            .O(N__15245),
            .I(N__15242));
    LocalMux I__3104 (
            .O(N__15242),
            .I(M_this_state_q_srsts_i_a2_1_8_1));
    CascadeMux I__3103 (
            .O(N__15239),
            .I(M_this_state_q_srsts_i_a2_1_7_1_cascade_));
    InMux I__3102 (
            .O(N__15236),
            .I(N__15233));
    LocalMux I__3101 (
            .O(N__15233),
            .I(M_this_state_q_srsts_i_a2_1_9_1));
    InMux I__3100 (
            .O(N__15230),
            .I(N__15227));
    LocalMux I__3099 (
            .O(N__15227),
            .I(M_this_state_q_srsts_i_a2_1_6_1));
    CascadeMux I__3098 (
            .O(N__15224),
            .I(N__15221));
    InMux I__3097 (
            .O(N__15221),
            .I(N__15217));
    InMux I__3096 (
            .O(N__15220),
            .I(N__15214));
    LocalMux I__3095 (
            .O(N__15217),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__3094 (
            .O(N__15214),
            .I(M_this_data_count_qZ0Z_0));
    CascadeMux I__3093 (
            .O(N__15209),
            .I(N__15206));
    InMux I__3092 (
            .O(N__15206),
            .I(N__15202));
    InMux I__3091 (
            .O(N__15205),
            .I(N__15199));
    LocalMux I__3090 (
            .O(N__15202),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__3089 (
            .O(N__15199),
            .I(M_this_data_count_qZ0Z_1));
    InMux I__3088 (
            .O(N__15194),
            .I(un1_M_this_data_count_q_cry_0));
    CascadeMux I__3087 (
            .O(N__15191),
            .I(N__15188));
    InMux I__3086 (
            .O(N__15188),
            .I(N__15184));
    InMux I__3085 (
            .O(N__15187),
            .I(N__15181));
    LocalMux I__3084 (
            .O(N__15184),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__3083 (
            .O(N__15181),
            .I(M_this_data_count_qZ0Z_2));
    InMux I__3082 (
            .O(N__15176),
            .I(un1_M_this_data_count_q_cry_1));
    CascadeMux I__3081 (
            .O(N__15173),
            .I(N__15170));
    InMux I__3080 (
            .O(N__15170),
            .I(N__15166));
    InMux I__3079 (
            .O(N__15169),
            .I(N__15163));
    LocalMux I__3078 (
            .O(N__15166),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__3077 (
            .O(N__15163),
            .I(M_this_data_count_qZ0Z_3));
    InMux I__3076 (
            .O(N__15158),
            .I(un1_M_this_data_count_q_cry_2));
    InMux I__3075 (
            .O(N__15155),
            .I(N__15152));
    LocalMux I__3074 (
            .O(N__15152),
            .I(\this_ppu.M_haddress_d8lto6_4 ));
    InMux I__3073 (
            .O(N__15149),
            .I(N__15146));
    LocalMux I__3072 (
            .O(N__15146),
            .I(\this_ppu.un1_M_line_clk_out_ns_1_0 ));
    InMux I__3071 (
            .O(N__15143),
            .I(N__15140));
    LocalMux I__3070 (
            .O(N__15140),
            .I(N__15134));
    InMux I__3069 (
            .O(N__15139),
            .I(N__15129));
    InMux I__3068 (
            .O(N__15138),
            .I(N__15129));
    InMux I__3067 (
            .O(N__15137),
            .I(N__15126));
    Span4Mux_v I__3066 (
            .O(N__15134),
            .I(N__15121));
    LocalMux I__3065 (
            .O(N__15129),
            .I(N__15121));
    LocalMux I__3064 (
            .O(N__15126),
            .I(M_this_vga_signals_line_clk_0));
    Odrv4 I__3063 (
            .O(N__15121),
            .I(M_this_vga_signals_line_clk_0));
    CascadeMux I__3062 (
            .O(N__15116),
            .I(N__15111));
    CascadeMux I__3061 (
            .O(N__15115),
            .I(N__15108));
    CascadeMux I__3060 (
            .O(N__15114),
            .I(N__15105));
    InMux I__3059 (
            .O(N__15111),
            .I(N__15102));
    InMux I__3058 (
            .O(N__15108),
            .I(N__15096));
    InMux I__3057 (
            .O(N__15105),
            .I(N__15096));
    LocalMux I__3056 (
            .O(N__15102),
            .I(N__15093));
    InMux I__3055 (
            .O(N__15101),
            .I(N__15090));
    LocalMux I__3054 (
            .O(N__15096),
            .I(N__15087));
    Span4Mux_h I__3053 (
            .O(N__15093),
            .I(N__15084));
    LocalMux I__3052 (
            .O(N__15090),
            .I(\this_ppu.line_clk.M_last_qZ0 ));
    Odrv12 I__3051 (
            .O(N__15087),
            .I(\this_ppu.line_clk.M_last_qZ0 ));
    Odrv4 I__3050 (
            .O(N__15084),
            .I(\this_ppu.line_clk.M_last_qZ0 ));
    InMux I__3049 (
            .O(N__15077),
            .I(N__15074));
    LocalMux I__3048 (
            .O(N__15074),
            .I(N__15070));
    InMux I__3047 (
            .O(N__15073),
            .I(N__15067));
    Span4Mux_h I__3046 (
            .O(N__15070),
            .I(N__15064));
    LocalMux I__3045 (
            .O(N__15067),
            .I(N__15061));
    Odrv4 I__3044 (
            .O(N__15064),
            .I(\this_vga_signals.M_vcounter_d8 ));
    Odrv12 I__3043 (
            .O(N__15061),
            .I(\this_vga_signals.M_vcounter_d8 ));
    SRMux I__3042 (
            .O(N__15056),
            .I(N__15052));
    SRMux I__3041 (
            .O(N__15055),
            .I(N__15049));
    LocalMux I__3040 (
            .O(N__15052),
            .I(N__15044));
    LocalMux I__3039 (
            .O(N__15049),
            .I(N__15041));
    SRMux I__3038 (
            .O(N__15048),
            .I(N__15038));
    InMux I__3037 (
            .O(N__15047),
            .I(N__15034));
    Span4Mux_v I__3036 (
            .O(N__15044),
            .I(N__15029));
    Span4Mux_v I__3035 (
            .O(N__15041),
            .I(N__15029));
    LocalMux I__3034 (
            .O(N__15038),
            .I(N__15026));
    SRMux I__3033 (
            .O(N__15037),
            .I(N__15023));
    LocalMux I__3032 (
            .O(N__15034),
            .I(N__15020));
    Span4Mux_h I__3031 (
            .O(N__15029),
            .I(N__15016));
    Span12Mux_s11_v I__3030 (
            .O(N__15026),
            .I(N__15011));
    LocalMux I__3029 (
            .O(N__15023),
            .I(N__15011));
    Span4Mux_h I__3028 (
            .O(N__15020),
            .I(N__15008));
    InMux I__3027 (
            .O(N__15019),
            .I(N__15005));
    Odrv4 I__3026 (
            .O(N__15016),
            .I(\this_vga_signals.M_vcounter_q_249_0 ));
    Odrv12 I__3025 (
            .O(N__15011),
            .I(\this_vga_signals.M_vcounter_q_249_0 ));
    Odrv4 I__3024 (
            .O(N__15008),
            .I(\this_vga_signals.M_vcounter_q_249_0 ));
    LocalMux I__3023 (
            .O(N__15005),
            .I(\this_vga_signals.M_vcounter_q_249_0 ));
    IoInMux I__3022 (
            .O(N__14996),
            .I(N__14993));
    LocalMux I__3021 (
            .O(N__14993),
            .I(N__14990));
    IoSpan4Mux I__3020 (
            .O(N__14990),
            .I(N__14987));
    Span4Mux_s2_h I__3019 (
            .O(N__14987),
            .I(N__14984));
    Sp12to4 I__3018 (
            .O(N__14984),
            .I(N__14981));
    Odrv12 I__3017 (
            .O(N__14981),
            .I(\this_vga_signals.M_vcounter_q_esr_RNIRO2H5Z0Z_9 ));
    InMux I__3016 (
            .O(N__14978),
            .I(N__14975));
    LocalMux I__3015 (
            .O(N__14975),
            .I(N__14972));
    Span4Mux_v I__3014 (
            .O(N__14972),
            .I(N__14969));
    Odrv4 I__3013 (
            .O(N__14969),
            .I(M_this_sprites_address_q_RNO_1Z0Z_0));
    InMux I__3012 (
            .O(N__14966),
            .I(N__14961));
    InMux I__3011 (
            .O(N__14965),
            .I(N__14956));
    InMux I__3010 (
            .O(N__14964),
            .I(N__14956));
    LocalMux I__3009 (
            .O(N__14961),
            .I(\this_pixel_clk.M_counter_qZ0Z_0 ));
    LocalMux I__3008 (
            .O(N__14956),
            .I(\this_pixel_clk.M_counter_qZ0Z_0 ));
    InMux I__3007 (
            .O(N__14951),
            .I(N__14948));
    LocalMux I__3006 (
            .O(N__14948),
            .I(M_this_sprites_address_q_RNO_1Z0Z_9));
    InMux I__3005 (
            .O(N__14945),
            .I(N__14942));
    LocalMux I__3004 (
            .O(N__14942),
            .I(un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0));
    InMux I__3003 (
            .O(N__14939),
            .I(N__14936));
    LocalMux I__3002 (
            .O(N__14936),
            .I(M_this_sprites_address_q_3_ns_1_6));
    InMux I__3001 (
            .O(N__14933),
            .I(N__14930));
    LocalMux I__3000 (
            .O(N__14930),
            .I(M_this_sprites_address_q_RNO_1Z0Z_6));
    CascadeMux I__2999 (
            .O(N__14927),
            .I(N__14924));
    CascadeBuf I__2998 (
            .O(N__14924),
            .I(N__14921));
    CascadeMux I__2997 (
            .O(N__14921),
            .I(N__14918));
    CascadeBuf I__2996 (
            .O(N__14918),
            .I(N__14915));
    CascadeMux I__2995 (
            .O(N__14915),
            .I(N__14912));
    CascadeBuf I__2994 (
            .O(N__14912),
            .I(N__14909));
    CascadeMux I__2993 (
            .O(N__14909),
            .I(N__14906));
    CascadeBuf I__2992 (
            .O(N__14906),
            .I(N__14903));
    CascadeMux I__2991 (
            .O(N__14903),
            .I(N__14900));
    CascadeBuf I__2990 (
            .O(N__14900),
            .I(N__14897));
    CascadeMux I__2989 (
            .O(N__14897),
            .I(N__14894));
    CascadeBuf I__2988 (
            .O(N__14894),
            .I(N__14891));
    CascadeMux I__2987 (
            .O(N__14891),
            .I(N__14888));
    CascadeBuf I__2986 (
            .O(N__14888),
            .I(N__14885));
    CascadeMux I__2985 (
            .O(N__14885),
            .I(N__14882));
    CascadeBuf I__2984 (
            .O(N__14882),
            .I(N__14879));
    CascadeMux I__2983 (
            .O(N__14879),
            .I(N__14876));
    CascadeBuf I__2982 (
            .O(N__14876),
            .I(N__14873));
    CascadeMux I__2981 (
            .O(N__14873),
            .I(N__14870));
    CascadeBuf I__2980 (
            .O(N__14870),
            .I(N__14867));
    CascadeMux I__2979 (
            .O(N__14867),
            .I(N__14864));
    CascadeBuf I__2978 (
            .O(N__14864),
            .I(N__14861));
    CascadeMux I__2977 (
            .O(N__14861),
            .I(N__14858));
    CascadeBuf I__2976 (
            .O(N__14858),
            .I(N__14855));
    CascadeMux I__2975 (
            .O(N__14855),
            .I(N__14852));
    CascadeBuf I__2974 (
            .O(N__14852),
            .I(N__14849));
    CascadeMux I__2973 (
            .O(N__14849),
            .I(N__14846));
    CascadeBuf I__2972 (
            .O(N__14846),
            .I(N__14843));
    CascadeMux I__2971 (
            .O(N__14843),
            .I(N__14840));
    CascadeBuf I__2970 (
            .O(N__14840),
            .I(N__14837));
    CascadeMux I__2969 (
            .O(N__14837),
            .I(N__14834));
    InMux I__2968 (
            .O(N__14834),
            .I(N__14831));
    LocalMux I__2967 (
            .O(N__14831),
            .I(N__14826));
    InMux I__2966 (
            .O(N__14830),
            .I(N__14823));
    InMux I__2965 (
            .O(N__14829),
            .I(N__14820));
    Span12Mux_s9_v I__2964 (
            .O(N__14826),
            .I(N__14817));
    LocalMux I__2963 (
            .O(N__14823),
            .I(M_this_sprites_address_qZ0Z_6));
    LocalMux I__2962 (
            .O(N__14820),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv12 I__2961 (
            .O(N__14817),
            .I(M_this_sprites_address_qZ0Z_6));
    CascadeMux I__2960 (
            .O(N__14810),
            .I(N__14807));
    CascadeBuf I__2959 (
            .O(N__14807),
            .I(N__14804));
    CascadeMux I__2958 (
            .O(N__14804),
            .I(N__14801));
    CascadeBuf I__2957 (
            .O(N__14801),
            .I(N__14798));
    CascadeMux I__2956 (
            .O(N__14798),
            .I(N__14795));
    CascadeBuf I__2955 (
            .O(N__14795),
            .I(N__14792));
    CascadeMux I__2954 (
            .O(N__14792),
            .I(N__14789));
    CascadeBuf I__2953 (
            .O(N__14789),
            .I(N__14786));
    CascadeMux I__2952 (
            .O(N__14786),
            .I(N__14783));
    CascadeBuf I__2951 (
            .O(N__14783),
            .I(N__14780));
    CascadeMux I__2950 (
            .O(N__14780),
            .I(N__14777));
    CascadeBuf I__2949 (
            .O(N__14777),
            .I(N__14774));
    CascadeMux I__2948 (
            .O(N__14774),
            .I(N__14771));
    CascadeBuf I__2947 (
            .O(N__14771),
            .I(N__14768));
    CascadeMux I__2946 (
            .O(N__14768),
            .I(N__14765));
    CascadeBuf I__2945 (
            .O(N__14765),
            .I(N__14762));
    CascadeMux I__2944 (
            .O(N__14762),
            .I(N__14759));
    CascadeBuf I__2943 (
            .O(N__14759),
            .I(N__14756));
    CascadeMux I__2942 (
            .O(N__14756),
            .I(N__14753));
    CascadeBuf I__2941 (
            .O(N__14753),
            .I(N__14750));
    CascadeMux I__2940 (
            .O(N__14750),
            .I(N__14747));
    CascadeBuf I__2939 (
            .O(N__14747),
            .I(N__14744));
    CascadeMux I__2938 (
            .O(N__14744),
            .I(N__14741));
    CascadeBuf I__2937 (
            .O(N__14741),
            .I(N__14738));
    CascadeMux I__2936 (
            .O(N__14738),
            .I(N__14735));
    CascadeBuf I__2935 (
            .O(N__14735),
            .I(N__14732));
    CascadeMux I__2934 (
            .O(N__14732),
            .I(N__14729));
    CascadeBuf I__2933 (
            .O(N__14729),
            .I(N__14726));
    CascadeMux I__2932 (
            .O(N__14726),
            .I(N__14723));
    CascadeBuf I__2931 (
            .O(N__14723),
            .I(N__14720));
    CascadeMux I__2930 (
            .O(N__14720),
            .I(N__14717));
    InMux I__2929 (
            .O(N__14717),
            .I(N__14714));
    LocalMux I__2928 (
            .O(N__14714),
            .I(N__14711));
    Span4Mux_s2_v I__2927 (
            .O(N__14711),
            .I(N__14708));
    Span4Mux_h I__2926 (
            .O(N__14708),
            .I(N__14705));
    Span4Mux_h I__2925 (
            .O(N__14705),
            .I(N__14700));
    InMux I__2924 (
            .O(N__14704),
            .I(N__14697));
    InMux I__2923 (
            .O(N__14703),
            .I(N__14694));
    Span4Mux_v I__2922 (
            .O(N__14700),
            .I(N__14691));
    LocalMux I__2921 (
            .O(N__14697),
            .I(M_this_sprites_address_qZ0Z_9));
    LocalMux I__2920 (
            .O(N__14694),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv4 I__2919 (
            .O(N__14691),
            .I(M_this_sprites_address_qZ0Z_9));
    CascadeMux I__2918 (
            .O(N__14684),
            .I(N__14681));
    InMux I__2917 (
            .O(N__14681),
            .I(N__14678));
    LocalMux I__2916 (
            .O(N__14678),
            .I(N__14675));
    Odrv4 I__2915 (
            .O(N__14675),
            .I(M_this_sprites_address_q_3_ns_1_9));
    CascadeMux I__2914 (
            .O(N__14672),
            .I(N__14669));
    CascadeBuf I__2913 (
            .O(N__14669),
            .I(N__14666));
    CascadeMux I__2912 (
            .O(N__14666),
            .I(N__14663));
    CascadeBuf I__2911 (
            .O(N__14663),
            .I(N__14660));
    CascadeMux I__2910 (
            .O(N__14660),
            .I(N__14657));
    CascadeBuf I__2909 (
            .O(N__14657),
            .I(N__14654));
    CascadeMux I__2908 (
            .O(N__14654),
            .I(N__14651));
    CascadeBuf I__2907 (
            .O(N__14651),
            .I(N__14648));
    CascadeMux I__2906 (
            .O(N__14648),
            .I(N__14645));
    CascadeBuf I__2905 (
            .O(N__14645),
            .I(N__14642));
    CascadeMux I__2904 (
            .O(N__14642),
            .I(N__14639));
    CascadeBuf I__2903 (
            .O(N__14639),
            .I(N__14636));
    CascadeMux I__2902 (
            .O(N__14636),
            .I(N__14633));
    CascadeBuf I__2901 (
            .O(N__14633),
            .I(N__14630));
    CascadeMux I__2900 (
            .O(N__14630),
            .I(N__14627));
    CascadeBuf I__2899 (
            .O(N__14627),
            .I(N__14624));
    CascadeMux I__2898 (
            .O(N__14624),
            .I(N__14621));
    CascadeBuf I__2897 (
            .O(N__14621),
            .I(N__14618));
    CascadeMux I__2896 (
            .O(N__14618),
            .I(N__14615));
    CascadeBuf I__2895 (
            .O(N__14615),
            .I(N__14612));
    CascadeMux I__2894 (
            .O(N__14612),
            .I(N__14609));
    CascadeBuf I__2893 (
            .O(N__14609),
            .I(N__14606));
    CascadeMux I__2892 (
            .O(N__14606),
            .I(N__14603));
    CascadeBuf I__2891 (
            .O(N__14603),
            .I(N__14600));
    CascadeMux I__2890 (
            .O(N__14600),
            .I(N__14597));
    CascadeBuf I__2889 (
            .O(N__14597),
            .I(N__14594));
    CascadeMux I__2888 (
            .O(N__14594),
            .I(N__14591));
    CascadeBuf I__2887 (
            .O(N__14591),
            .I(N__14588));
    CascadeMux I__2886 (
            .O(N__14588),
            .I(N__14585));
    CascadeBuf I__2885 (
            .O(N__14585),
            .I(N__14582));
    CascadeMux I__2884 (
            .O(N__14582),
            .I(N__14579));
    InMux I__2883 (
            .O(N__14579),
            .I(N__14576));
    LocalMux I__2882 (
            .O(N__14576),
            .I(N__14573));
    Span4Mux_h I__2881 (
            .O(N__14573),
            .I(N__14570));
    Span4Mux_h I__2880 (
            .O(N__14570),
            .I(N__14566));
    InMux I__2879 (
            .O(N__14569),
            .I(N__14563));
    Span4Mux_h I__2878 (
            .O(N__14566),
            .I(N__14559));
    LocalMux I__2877 (
            .O(N__14563),
            .I(N__14556));
    InMux I__2876 (
            .O(N__14562),
            .I(N__14553));
    Span4Mux_v I__2875 (
            .O(N__14559),
            .I(N__14550));
    Odrv4 I__2874 (
            .O(N__14556),
            .I(M_this_sprites_address_qZ0Z_1));
    LocalMux I__2873 (
            .O(N__14553),
            .I(M_this_sprites_address_qZ0Z_1));
    Odrv4 I__2872 (
            .O(N__14550),
            .I(M_this_sprites_address_qZ0Z_1));
    InMux I__2871 (
            .O(N__14543),
            .I(N__14540));
    LocalMux I__2870 (
            .O(N__14540),
            .I(M_this_sprites_address_q_3_ns_1_1));
    CascadeMux I__2869 (
            .O(N__14537),
            .I(\this_ppu.un1_M_haddress_q_c3_cascade_ ));
    InMux I__2868 (
            .O(N__14534),
            .I(N__14528));
    InMux I__2867 (
            .O(N__14533),
            .I(N__14528));
    LocalMux I__2866 (
            .O(N__14528),
            .I(N__14525));
    Span4Mux_v I__2865 (
            .O(N__14525),
            .I(N__14516));
    InMux I__2864 (
            .O(N__14524),
            .I(N__14505));
    InMux I__2863 (
            .O(N__14523),
            .I(N__14505));
    InMux I__2862 (
            .O(N__14522),
            .I(N__14505));
    InMux I__2861 (
            .O(N__14521),
            .I(N__14505));
    InMux I__2860 (
            .O(N__14520),
            .I(N__14505));
    IoInMux I__2859 (
            .O(N__14519),
            .I(N__14502));
    Span4Mux_h I__2858 (
            .O(N__14516),
            .I(N__14498));
    LocalMux I__2857 (
            .O(N__14505),
            .I(N__14495));
    LocalMux I__2856 (
            .O(N__14502),
            .I(N__14492));
    InMux I__2855 (
            .O(N__14501),
            .I(N__14489));
    Sp12to4 I__2854 (
            .O(N__14498),
            .I(N__14484));
    Span12Mux_s8_h I__2853 (
            .O(N__14495),
            .I(N__14484));
    Span12Mux_s1_v I__2852 (
            .O(N__14492),
            .I(N__14481));
    LocalMux I__2851 (
            .O(N__14489),
            .I(M_this_state_q_nss_0));
    Odrv12 I__2850 (
            .O(N__14484),
            .I(M_this_state_q_nss_0));
    Odrv12 I__2849 (
            .O(N__14481),
            .I(M_this_state_q_nss_0));
    InMux I__2848 (
            .O(N__14474),
            .I(N__14468));
    InMux I__2847 (
            .O(N__14473),
            .I(N__14468));
    LocalMux I__2846 (
            .O(N__14468),
            .I(\this_pixel_clk.M_counter_q_i_1 ));
    CascadeMux I__2845 (
            .O(N__14465),
            .I(N__14462));
    InMux I__2844 (
            .O(N__14462),
            .I(N__14459));
    LocalMux I__2843 (
            .O(N__14459),
            .I(N__14456));
    Span4Mux_h I__2842 (
            .O(N__14456),
            .I(N__14453));
    Odrv4 I__2841 (
            .O(N__14453),
            .I(M_this_state_q_srsts_i_1_2));
    CascadeMux I__2840 (
            .O(N__14450),
            .I(N__14447));
    InMux I__2839 (
            .O(N__14447),
            .I(N__14441));
    InMux I__2838 (
            .O(N__14446),
            .I(N__14441));
    LocalMux I__2837 (
            .O(N__14441),
            .I(N__14438));
    Span4Mux_v I__2836 (
            .O(N__14438),
            .I(N__14435));
    Sp12to4 I__2835 (
            .O(N__14435),
            .I(N__14432));
    Span12Mux_h I__2834 (
            .O(N__14432),
            .I(N__14428));
    InMux I__2833 (
            .O(N__14431),
            .I(N__14425));
    Odrv12 I__2832 (
            .O(N__14428),
            .I(port_rw_in));
    LocalMux I__2831 (
            .O(N__14425),
            .I(port_rw_in));
    CascadeMux I__2830 (
            .O(N__14420),
            .I(N_171_0_cascade_));
    InMux I__2829 (
            .O(N__14417),
            .I(N__14414));
    LocalMux I__2828 (
            .O(N__14414),
            .I(N__14411));
    Odrv4 I__2827 (
            .O(N__14411),
            .I(N_176_0));
    CascadeMux I__2826 (
            .O(N__14408),
            .I(N__14403));
    InMux I__2825 (
            .O(N__14407),
            .I(N__14400));
    InMux I__2824 (
            .O(N__14406),
            .I(N__14395));
    InMux I__2823 (
            .O(N__14403),
            .I(N__14395));
    LocalMux I__2822 (
            .O(N__14400),
            .I(N__14390));
    LocalMux I__2821 (
            .O(N__14395),
            .I(N__14390));
    Odrv4 I__2820 (
            .O(N__14390),
            .I(M_this_state_qZ0Z_4));
    CascadeMux I__2819 (
            .O(N__14387),
            .I(N__14383));
    InMux I__2818 (
            .O(N__14386),
            .I(N__14380));
    InMux I__2817 (
            .O(N__14383),
            .I(N__14377));
    LocalMux I__2816 (
            .O(N__14380),
            .I(N_153_0));
    LocalMux I__2815 (
            .O(N__14377),
            .I(N_153_0));
    InMux I__2814 (
            .O(N__14372),
            .I(N__14369));
    LocalMux I__2813 (
            .O(N__14369),
            .I(M_this_sprites_address_q_RNO_1Z0Z_2));
    InMux I__2812 (
            .O(N__14366),
            .I(N__14361));
    InMux I__2811 (
            .O(N__14365),
            .I(N__14358));
    InMux I__2810 (
            .O(N__14364),
            .I(N__14355));
    LocalMux I__2809 (
            .O(N__14361),
            .I(N__14352));
    LocalMux I__2808 (
            .O(N__14358),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    LocalMux I__2807 (
            .O(N__14355),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    Odrv4 I__2806 (
            .O(N__14352),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    InMux I__2805 (
            .O(N__14345),
            .I(N__14342));
    LocalMux I__2804 (
            .O(N__14342),
            .I(\this_vga_signals.un1_M_hcounter_d7_1_0 ));
    CascadeMux I__2803 (
            .O(N__14339),
            .I(\this_vga_signals.CO0_cascade_ ));
    InMux I__2802 (
            .O(N__14336),
            .I(N__14331));
    InMux I__2801 (
            .O(N__14335),
            .I(N__14326));
    InMux I__2800 (
            .O(N__14334),
            .I(N__14326));
    LocalMux I__2799 (
            .O(N__14331),
            .I(N__14323));
    LocalMux I__2798 (
            .O(N__14326),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    Odrv4 I__2797 (
            .O(N__14323),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    InMux I__2796 (
            .O(N__14318),
            .I(N__14315));
    LocalMux I__2795 (
            .O(N__14315),
            .I(\this_ppu.M_line_clk_out_0 ));
    InMux I__2794 (
            .O(N__14312),
            .I(N__14309));
    LocalMux I__2793 (
            .O(N__14309),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__2792 (
            .O(N__14306),
            .I(N__14294));
    InMux I__2791 (
            .O(N__14305),
            .I(N__14294));
    InMux I__2790 (
            .O(N__14304),
            .I(N__14294));
    InMux I__2789 (
            .O(N__14303),
            .I(N__14294));
    LocalMux I__2788 (
            .O(N__14294),
            .I(N__14291));
    Sp12to4 I__2787 (
            .O(N__14291),
            .I(N__14288));
    Span12Mux_v I__2786 (
            .O(N__14288),
            .I(N__14285));
    Odrv12 I__2785 (
            .O(N__14285),
            .I(rst_n_c));
    InMux I__2784 (
            .O(N__14282),
            .I(N__14279));
    LocalMux I__2783 (
            .O(N__14279),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__2782 (
            .O(N__14276),
            .I(N__14273));
    LocalMux I__2781 (
            .O(N__14273),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    InMux I__2780 (
            .O(N__14270),
            .I(N__14247));
    InMux I__2779 (
            .O(N__14269),
            .I(N__14247));
    InMux I__2778 (
            .O(N__14268),
            .I(N__14247));
    InMux I__2777 (
            .O(N__14267),
            .I(N__14247));
    InMux I__2776 (
            .O(N__14266),
            .I(N__14240));
    InMux I__2775 (
            .O(N__14265),
            .I(N__14240));
    InMux I__2774 (
            .O(N__14264),
            .I(N__14240));
    InMux I__2773 (
            .O(N__14263),
            .I(N__14236));
    CEMux I__2772 (
            .O(N__14262),
            .I(N__14232));
    InMux I__2771 (
            .O(N__14261),
            .I(N__14228));
    InMux I__2770 (
            .O(N__14260),
            .I(N__14225));
    InMux I__2769 (
            .O(N__14259),
            .I(N__14220));
    InMux I__2768 (
            .O(N__14258),
            .I(N__14220));
    InMux I__2767 (
            .O(N__14257),
            .I(N__14215));
    InMux I__2766 (
            .O(N__14256),
            .I(N__14215));
    LocalMux I__2765 (
            .O(N__14247),
            .I(N__14212));
    LocalMux I__2764 (
            .O(N__14240),
            .I(N__14209));
    InMux I__2763 (
            .O(N__14239),
            .I(N__14206));
    LocalMux I__2762 (
            .O(N__14236),
            .I(N__14201));
    InMux I__2761 (
            .O(N__14235),
            .I(N__14198));
    LocalMux I__2760 (
            .O(N__14232),
            .I(N__14195));
    InMux I__2759 (
            .O(N__14231),
            .I(N__14192));
    LocalMux I__2758 (
            .O(N__14228),
            .I(N__14187));
    LocalMux I__2757 (
            .O(N__14225),
            .I(N__14187));
    LocalMux I__2756 (
            .O(N__14220),
            .I(N__14184));
    LocalMux I__2755 (
            .O(N__14215),
            .I(N__14181));
    Span4Mux_v I__2754 (
            .O(N__14212),
            .I(N__14178));
    Span4Mux_v I__2753 (
            .O(N__14209),
            .I(N__14173));
    LocalMux I__2752 (
            .O(N__14206),
            .I(N__14173));
    InMux I__2751 (
            .O(N__14205),
            .I(N__14168));
    InMux I__2750 (
            .O(N__14204),
            .I(N__14168));
    Span12Mux_s3_h I__2749 (
            .O(N__14201),
            .I(N__14165));
    LocalMux I__2748 (
            .O(N__14198),
            .I(N__14162));
    Span4Mux_v I__2747 (
            .O(N__14195),
            .I(N__14159));
    LocalMux I__2746 (
            .O(N__14192),
            .I(N__14154));
    Span4Mux_v I__2745 (
            .O(N__14187),
            .I(N__14154));
    Span4Mux_h I__2744 (
            .O(N__14184),
            .I(N__14149));
    Span4Mux_h I__2743 (
            .O(N__14181),
            .I(N__14149));
    Span4Mux_h I__2742 (
            .O(N__14178),
            .I(N__14144));
    Span4Mux_h I__2741 (
            .O(N__14173),
            .I(N__14144));
    LocalMux I__2740 (
            .O(N__14168),
            .I(N__14139));
    Span12Mux_h I__2739 (
            .O(N__14165),
            .I(N__14139));
    Span4Mux_v I__2738 (
            .O(N__14162),
            .I(N__14132));
    Span4Mux_h I__2737 (
            .O(N__14159),
            .I(N__14132));
    Span4Mux_h I__2736 (
            .O(N__14154),
            .I(N__14132));
    Odrv4 I__2735 (
            .O(N__14149),
            .I(M_counter_q_RNIFKS8_1));
    Odrv4 I__2734 (
            .O(N__14144),
            .I(M_counter_q_RNIFKS8_1));
    Odrv12 I__2733 (
            .O(N__14139),
            .I(M_counter_q_RNIFKS8_1));
    Odrv4 I__2732 (
            .O(N__14132),
            .I(M_counter_q_RNIFKS8_1));
    CascadeMux I__2731 (
            .O(N__14123),
            .I(M_counter_q_RNIFKS8_1_cascade_));
    CascadeMux I__2730 (
            .O(N__14120),
            .I(N__14111));
    InMux I__2729 (
            .O(N__14119),
            .I(N__14102));
    InMux I__2728 (
            .O(N__14118),
            .I(N__14102));
    InMux I__2727 (
            .O(N__14117),
            .I(N__14102));
    InMux I__2726 (
            .O(N__14116),
            .I(N__14096));
    InMux I__2725 (
            .O(N__14115),
            .I(N__14096));
    InMux I__2724 (
            .O(N__14114),
            .I(N__14093));
    InMux I__2723 (
            .O(N__14111),
            .I(N__14090));
    InMux I__2722 (
            .O(N__14110),
            .I(N__14085));
    InMux I__2721 (
            .O(N__14109),
            .I(N__14085));
    LocalMux I__2720 (
            .O(N__14102),
            .I(N__14082));
    InMux I__2719 (
            .O(N__14101),
            .I(N__14079));
    LocalMux I__2718 (
            .O(N__14096),
            .I(N__14076));
    LocalMux I__2717 (
            .O(N__14093),
            .I(N__14071));
    LocalMux I__2716 (
            .O(N__14090),
            .I(N__14071));
    LocalMux I__2715 (
            .O(N__14085),
            .I(N__14068));
    Span4Mux_v I__2714 (
            .O(N__14082),
            .I(N__14063));
    LocalMux I__2713 (
            .O(N__14079),
            .I(N__14063));
    Span4Mux_v I__2712 (
            .O(N__14076),
            .I(N__14060));
    Span4Mux_v I__2711 (
            .O(N__14071),
            .I(N__14057));
    Span4Mux_h I__2710 (
            .O(N__14068),
            .I(N__14054));
    Span4Mux_h I__2709 (
            .O(N__14063),
            .I(N__14051));
    Odrv4 I__2708 (
            .O(N__14060),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__2707 (
            .O(N__14057),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__2706 (
            .O(N__14054),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__2705 (
            .O(N__14051),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    InMux I__2704 (
            .O(N__14042),
            .I(un1_M_this_sprites_address_q_cry_12));
    InMux I__2703 (
            .O(N__14039),
            .I(N__14036));
    LocalMux I__2702 (
            .O(N__14036),
            .I(M_this_sprites_address_q_RNO_1Z0Z_8));
    CascadeMux I__2701 (
            .O(N__14033),
            .I(M_this_sprites_address_q_3_ns_1_8_cascade_));
    CascadeMux I__2700 (
            .O(N__14030),
            .I(N__14027));
    CascadeBuf I__2699 (
            .O(N__14027),
            .I(N__14024));
    CascadeMux I__2698 (
            .O(N__14024),
            .I(N__14021));
    CascadeBuf I__2697 (
            .O(N__14021),
            .I(N__14018));
    CascadeMux I__2696 (
            .O(N__14018),
            .I(N__14015));
    CascadeBuf I__2695 (
            .O(N__14015),
            .I(N__14012));
    CascadeMux I__2694 (
            .O(N__14012),
            .I(N__14009));
    CascadeBuf I__2693 (
            .O(N__14009),
            .I(N__14006));
    CascadeMux I__2692 (
            .O(N__14006),
            .I(N__14003));
    CascadeBuf I__2691 (
            .O(N__14003),
            .I(N__14000));
    CascadeMux I__2690 (
            .O(N__14000),
            .I(N__13997));
    CascadeBuf I__2689 (
            .O(N__13997),
            .I(N__13994));
    CascadeMux I__2688 (
            .O(N__13994),
            .I(N__13991));
    CascadeBuf I__2687 (
            .O(N__13991),
            .I(N__13988));
    CascadeMux I__2686 (
            .O(N__13988),
            .I(N__13985));
    CascadeBuf I__2685 (
            .O(N__13985),
            .I(N__13982));
    CascadeMux I__2684 (
            .O(N__13982),
            .I(N__13979));
    CascadeBuf I__2683 (
            .O(N__13979),
            .I(N__13976));
    CascadeMux I__2682 (
            .O(N__13976),
            .I(N__13973));
    CascadeBuf I__2681 (
            .O(N__13973),
            .I(N__13970));
    CascadeMux I__2680 (
            .O(N__13970),
            .I(N__13967));
    CascadeBuf I__2679 (
            .O(N__13967),
            .I(N__13964));
    CascadeMux I__2678 (
            .O(N__13964),
            .I(N__13961));
    CascadeBuf I__2677 (
            .O(N__13961),
            .I(N__13958));
    CascadeMux I__2676 (
            .O(N__13958),
            .I(N__13955));
    CascadeBuf I__2675 (
            .O(N__13955),
            .I(N__13952));
    CascadeMux I__2674 (
            .O(N__13952),
            .I(N__13949));
    CascadeBuf I__2673 (
            .O(N__13949),
            .I(N__13946));
    CascadeMux I__2672 (
            .O(N__13946),
            .I(N__13943));
    CascadeBuf I__2671 (
            .O(N__13943),
            .I(N__13940));
    CascadeMux I__2670 (
            .O(N__13940),
            .I(N__13937));
    InMux I__2669 (
            .O(N__13937),
            .I(N__13934));
    LocalMux I__2668 (
            .O(N__13934),
            .I(N__13931));
    Span4Mux_h I__2667 (
            .O(N__13931),
            .I(N__13928));
    Span4Mux_h I__2666 (
            .O(N__13928),
            .I(N__13925));
    Span4Mux_v I__2665 (
            .O(N__13925),
            .I(N__13920));
    InMux I__2664 (
            .O(N__13924),
            .I(N__13917));
    InMux I__2663 (
            .O(N__13923),
            .I(N__13914));
    Span4Mux_v I__2662 (
            .O(N__13920),
            .I(N__13911));
    LocalMux I__2661 (
            .O(N__13917),
            .I(M_this_sprites_address_qZ0Z_8));
    LocalMux I__2660 (
            .O(N__13914),
            .I(M_this_sprites_address_qZ0Z_8));
    Odrv4 I__2659 (
            .O(N__13911),
            .I(M_this_sprites_address_qZ0Z_8));
    InMux I__2658 (
            .O(N__13904),
            .I(N__13901));
    LocalMux I__2657 (
            .O(N__13901),
            .I(\this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_11 ));
    InMux I__2656 (
            .O(N__13898),
            .I(N__13895));
    LocalMux I__2655 (
            .O(N__13895),
            .I(un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0));
    InMux I__2654 (
            .O(N__13892),
            .I(N__13889));
    LocalMux I__2653 (
            .O(N__13889),
            .I(\this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_12 ));
    InMux I__2652 (
            .O(N__13886),
            .I(N__13883));
    LocalMux I__2651 (
            .O(N__13883),
            .I(un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0));
    InMux I__2650 (
            .O(N__13880),
            .I(N__13877));
    LocalMux I__2649 (
            .O(N__13877),
            .I(N__13874));
    Odrv12 I__2648 (
            .O(N__13874),
            .I(M_this_sprites_address_q_RNO_1Z0Z_1));
    CascadeMux I__2647 (
            .O(N__13871),
            .I(\this_vga_signals.un1_M_hcounter_d7_1_0_cascade_ ));
    CascadeMux I__2646 (
            .O(N__13868),
            .I(N__13865));
    CascadeBuf I__2645 (
            .O(N__13865),
            .I(N__13862));
    CascadeMux I__2644 (
            .O(N__13862),
            .I(N__13859));
    CascadeBuf I__2643 (
            .O(N__13859),
            .I(N__13856));
    CascadeMux I__2642 (
            .O(N__13856),
            .I(N__13853));
    CascadeBuf I__2641 (
            .O(N__13853),
            .I(N__13850));
    CascadeMux I__2640 (
            .O(N__13850),
            .I(N__13847));
    CascadeBuf I__2639 (
            .O(N__13847),
            .I(N__13844));
    CascadeMux I__2638 (
            .O(N__13844),
            .I(N__13841));
    CascadeBuf I__2637 (
            .O(N__13841),
            .I(N__13838));
    CascadeMux I__2636 (
            .O(N__13838),
            .I(N__13835));
    CascadeBuf I__2635 (
            .O(N__13835),
            .I(N__13832));
    CascadeMux I__2634 (
            .O(N__13832),
            .I(N__13829));
    CascadeBuf I__2633 (
            .O(N__13829),
            .I(N__13826));
    CascadeMux I__2632 (
            .O(N__13826),
            .I(N__13823));
    CascadeBuf I__2631 (
            .O(N__13823),
            .I(N__13820));
    CascadeMux I__2630 (
            .O(N__13820),
            .I(N__13817));
    CascadeBuf I__2629 (
            .O(N__13817),
            .I(N__13814));
    CascadeMux I__2628 (
            .O(N__13814),
            .I(N__13811));
    CascadeBuf I__2627 (
            .O(N__13811),
            .I(N__13808));
    CascadeMux I__2626 (
            .O(N__13808),
            .I(N__13805));
    CascadeBuf I__2625 (
            .O(N__13805),
            .I(N__13802));
    CascadeMux I__2624 (
            .O(N__13802),
            .I(N__13799));
    CascadeBuf I__2623 (
            .O(N__13799),
            .I(N__13796));
    CascadeMux I__2622 (
            .O(N__13796),
            .I(N__13793));
    CascadeBuf I__2621 (
            .O(N__13793),
            .I(N__13790));
    CascadeMux I__2620 (
            .O(N__13790),
            .I(N__13787));
    CascadeBuf I__2619 (
            .O(N__13787),
            .I(N__13784));
    CascadeMux I__2618 (
            .O(N__13784),
            .I(N__13781));
    CascadeBuf I__2617 (
            .O(N__13781),
            .I(N__13778));
    CascadeMux I__2616 (
            .O(N__13778),
            .I(N__13775));
    InMux I__2615 (
            .O(N__13775),
            .I(N__13772));
    LocalMux I__2614 (
            .O(N__13772),
            .I(N__13767));
    InMux I__2613 (
            .O(N__13771),
            .I(N__13764));
    InMux I__2612 (
            .O(N__13770),
            .I(N__13761));
    Span12Mux_h I__2611 (
            .O(N__13767),
            .I(N__13758));
    LocalMux I__2610 (
            .O(N__13764),
            .I(M_this_sprites_address_qZ0Z_4));
    LocalMux I__2609 (
            .O(N__13761),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv12 I__2608 (
            .O(N__13758),
            .I(M_this_sprites_address_qZ0Z_4));
    InMux I__2607 (
            .O(N__13751),
            .I(N__13748));
    LocalMux I__2606 (
            .O(N__13748),
            .I(M_this_sprites_address_q_RNO_1Z0Z_4));
    InMux I__2605 (
            .O(N__13745),
            .I(un1_M_this_sprites_address_q_cry_3));
    CascadeMux I__2604 (
            .O(N__13742),
            .I(N__13739));
    CascadeBuf I__2603 (
            .O(N__13739),
            .I(N__13736));
    CascadeMux I__2602 (
            .O(N__13736),
            .I(N__13733));
    CascadeBuf I__2601 (
            .O(N__13733),
            .I(N__13730));
    CascadeMux I__2600 (
            .O(N__13730),
            .I(N__13727));
    CascadeBuf I__2599 (
            .O(N__13727),
            .I(N__13724));
    CascadeMux I__2598 (
            .O(N__13724),
            .I(N__13721));
    CascadeBuf I__2597 (
            .O(N__13721),
            .I(N__13718));
    CascadeMux I__2596 (
            .O(N__13718),
            .I(N__13715));
    CascadeBuf I__2595 (
            .O(N__13715),
            .I(N__13712));
    CascadeMux I__2594 (
            .O(N__13712),
            .I(N__13709));
    CascadeBuf I__2593 (
            .O(N__13709),
            .I(N__13706));
    CascadeMux I__2592 (
            .O(N__13706),
            .I(N__13703));
    CascadeBuf I__2591 (
            .O(N__13703),
            .I(N__13700));
    CascadeMux I__2590 (
            .O(N__13700),
            .I(N__13697));
    CascadeBuf I__2589 (
            .O(N__13697),
            .I(N__13694));
    CascadeMux I__2588 (
            .O(N__13694),
            .I(N__13691));
    CascadeBuf I__2587 (
            .O(N__13691),
            .I(N__13688));
    CascadeMux I__2586 (
            .O(N__13688),
            .I(N__13685));
    CascadeBuf I__2585 (
            .O(N__13685),
            .I(N__13682));
    CascadeMux I__2584 (
            .O(N__13682),
            .I(N__13679));
    CascadeBuf I__2583 (
            .O(N__13679),
            .I(N__13676));
    CascadeMux I__2582 (
            .O(N__13676),
            .I(N__13673));
    CascadeBuf I__2581 (
            .O(N__13673),
            .I(N__13670));
    CascadeMux I__2580 (
            .O(N__13670),
            .I(N__13667));
    CascadeBuf I__2579 (
            .O(N__13667),
            .I(N__13664));
    CascadeMux I__2578 (
            .O(N__13664),
            .I(N__13661));
    CascadeBuf I__2577 (
            .O(N__13661),
            .I(N__13658));
    CascadeMux I__2576 (
            .O(N__13658),
            .I(N__13655));
    CascadeBuf I__2575 (
            .O(N__13655),
            .I(N__13652));
    CascadeMux I__2574 (
            .O(N__13652),
            .I(N__13649));
    InMux I__2573 (
            .O(N__13649),
            .I(N__13646));
    LocalMux I__2572 (
            .O(N__13646),
            .I(N__13643));
    Span4Mux_s1_v I__2571 (
            .O(N__13643),
            .I(N__13640));
    Span4Mux_h I__2570 (
            .O(N__13640),
            .I(N__13637));
    Sp12to4 I__2569 (
            .O(N__13637),
            .I(N__13632));
    InMux I__2568 (
            .O(N__13636),
            .I(N__13629));
    InMux I__2567 (
            .O(N__13635),
            .I(N__13626));
    Span12Mux_s11_v I__2566 (
            .O(N__13632),
            .I(N__13623));
    LocalMux I__2565 (
            .O(N__13629),
            .I(M_this_sprites_address_qZ0Z_5));
    LocalMux I__2564 (
            .O(N__13626),
            .I(M_this_sprites_address_qZ0Z_5));
    Odrv12 I__2563 (
            .O(N__13623),
            .I(M_this_sprites_address_qZ0Z_5));
    InMux I__2562 (
            .O(N__13616),
            .I(N__13613));
    LocalMux I__2561 (
            .O(N__13613),
            .I(M_this_sprites_address_q_RNO_1Z0Z_5));
    InMux I__2560 (
            .O(N__13610),
            .I(un1_M_this_sprites_address_q_cry_4));
    InMux I__2559 (
            .O(N__13607),
            .I(un1_M_this_sprites_address_q_cry_5));
    CascadeMux I__2558 (
            .O(N__13604),
            .I(N__13601));
    CascadeBuf I__2557 (
            .O(N__13601),
            .I(N__13598));
    CascadeMux I__2556 (
            .O(N__13598),
            .I(N__13595));
    CascadeBuf I__2555 (
            .O(N__13595),
            .I(N__13592));
    CascadeMux I__2554 (
            .O(N__13592),
            .I(N__13589));
    CascadeBuf I__2553 (
            .O(N__13589),
            .I(N__13586));
    CascadeMux I__2552 (
            .O(N__13586),
            .I(N__13583));
    CascadeBuf I__2551 (
            .O(N__13583),
            .I(N__13580));
    CascadeMux I__2550 (
            .O(N__13580),
            .I(N__13577));
    CascadeBuf I__2549 (
            .O(N__13577),
            .I(N__13574));
    CascadeMux I__2548 (
            .O(N__13574),
            .I(N__13571));
    CascadeBuf I__2547 (
            .O(N__13571),
            .I(N__13568));
    CascadeMux I__2546 (
            .O(N__13568),
            .I(N__13565));
    CascadeBuf I__2545 (
            .O(N__13565),
            .I(N__13562));
    CascadeMux I__2544 (
            .O(N__13562),
            .I(N__13559));
    CascadeBuf I__2543 (
            .O(N__13559),
            .I(N__13556));
    CascadeMux I__2542 (
            .O(N__13556),
            .I(N__13553));
    CascadeBuf I__2541 (
            .O(N__13553),
            .I(N__13550));
    CascadeMux I__2540 (
            .O(N__13550),
            .I(N__13547));
    CascadeBuf I__2539 (
            .O(N__13547),
            .I(N__13544));
    CascadeMux I__2538 (
            .O(N__13544),
            .I(N__13541));
    CascadeBuf I__2537 (
            .O(N__13541),
            .I(N__13538));
    CascadeMux I__2536 (
            .O(N__13538),
            .I(N__13535));
    CascadeBuf I__2535 (
            .O(N__13535),
            .I(N__13532));
    CascadeMux I__2534 (
            .O(N__13532),
            .I(N__13529));
    CascadeBuf I__2533 (
            .O(N__13529),
            .I(N__13526));
    CascadeMux I__2532 (
            .O(N__13526),
            .I(N__13523));
    CascadeBuf I__2531 (
            .O(N__13523),
            .I(N__13520));
    CascadeMux I__2530 (
            .O(N__13520),
            .I(N__13517));
    CascadeBuf I__2529 (
            .O(N__13517),
            .I(N__13514));
    CascadeMux I__2528 (
            .O(N__13514),
            .I(N__13511));
    InMux I__2527 (
            .O(N__13511),
            .I(N__13508));
    LocalMux I__2526 (
            .O(N__13508),
            .I(N__13505));
    Sp12to4 I__2525 (
            .O(N__13505),
            .I(N__13500));
    InMux I__2524 (
            .O(N__13504),
            .I(N__13497));
    InMux I__2523 (
            .O(N__13503),
            .I(N__13494));
    Span12Mux_s11_v I__2522 (
            .O(N__13500),
            .I(N__13491));
    LocalMux I__2521 (
            .O(N__13497),
            .I(M_this_sprites_address_qZ0Z_7));
    LocalMux I__2520 (
            .O(N__13494),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv12 I__2519 (
            .O(N__13491),
            .I(M_this_sprites_address_qZ0Z_7));
    InMux I__2518 (
            .O(N__13484),
            .I(N__13481));
    LocalMux I__2517 (
            .O(N__13481),
            .I(M_this_sprites_address_q_RNO_1Z0Z_7));
    InMux I__2516 (
            .O(N__13478),
            .I(un1_M_this_sprites_address_q_cry_6));
    InMux I__2515 (
            .O(N__13475),
            .I(bfn_15_23_0_));
    InMux I__2514 (
            .O(N__13472),
            .I(un1_M_this_sprites_address_q_cry_8));
    InMux I__2513 (
            .O(N__13469),
            .I(un1_M_this_sprites_address_q_cry_9));
    InMux I__2512 (
            .O(N__13466),
            .I(un1_M_this_sprites_address_q_cry_10));
    InMux I__2511 (
            .O(N__13463),
            .I(un1_M_this_sprites_address_q_cry_11));
    InMux I__2510 (
            .O(N__13460),
            .I(N__13457));
    LocalMux I__2509 (
            .O(N__13457),
            .I(M_this_ppu_vga_is_drawing_0));
    CascadeMux I__2508 (
            .O(N__13454),
            .I(\this_ppu.M_line_clk_out_0_cascade_ ));
    InMux I__2507 (
            .O(N__13451),
            .I(N__13448));
    LocalMux I__2506 (
            .O(N__13448),
            .I(M_this_sprites_address_q_3_ns_1_5));
    InMux I__2505 (
            .O(N__13445),
            .I(N__13442));
    LocalMux I__2504 (
            .O(N__13442),
            .I(M_this_sprites_address_q_3_ns_1_4));
    CascadeMux I__2503 (
            .O(N__13439),
            .I(M_this_sprites_address_q_3_ns_1_7_cascade_));
    InMux I__2502 (
            .O(N__13436),
            .I(un1_M_this_sprites_address_q_cry_0));
    InMux I__2501 (
            .O(N__13433),
            .I(un1_M_this_sprites_address_q_cry_1));
    InMux I__2500 (
            .O(N__13430),
            .I(un1_M_this_sprites_address_q_cry_2));
    CascadeMux I__2499 (
            .O(N__13427),
            .I(N__13420));
    CascadeMux I__2498 (
            .O(N__13426),
            .I(N__13414));
    InMux I__2497 (
            .O(N__13425),
            .I(N__13411));
    InMux I__2496 (
            .O(N__13424),
            .I(N__13408));
    InMux I__2495 (
            .O(N__13423),
            .I(N__13405));
    InMux I__2494 (
            .O(N__13420),
            .I(N__13397));
    InMux I__2493 (
            .O(N__13419),
            .I(N__13394));
    InMux I__2492 (
            .O(N__13418),
            .I(N__13389));
    InMux I__2491 (
            .O(N__13417),
            .I(N__13389));
    InMux I__2490 (
            .O(N__13414),
            .I(N__13386));
    LocalMux I__2489 (
            .O(N__13411),
            .I(N__13381));
    LocalMux I__2488 (
            .O(N__13408),
            .I(N__13381));
    LocalMux I__2487 (
            .O(N__13405),
            .I(N__13378));
    InMux I__2486 (
            .O(N__13404),
            .I(N__13371));
    InMux I__2485 (
            .O(N__13403),
            .I(N__13371));
    InMux I__2484 (
            .O(N__13402),
            .I(N__13371));
    InMux I__2483 (
            .O(N__13401),
            .I(N__13368));
    InMux I__2482 (
            .O(N__13400),
            .I(N__13365));
    LocalMux I__2481 (
            .O(N__13397),
            .I(N__13358));
    LocalMux I__2480 (
            .O(N__13394),
            .I(N__13358));
    LocalMux I__2479 (
            .O(N__13389),
            .I(N__13353));
    LocalMux I__2478 (
            .O(N__13386),
            .I(N__13353));
    Span4Mux_v I__2477 (
            .O(N__13381),
            .I(N__13346));
    Span4Mux_h I__2476 (
            .O(N__13378),
            .I(N__13346));
    LocalMux I__2475 (
            .O(N__13371),
            .I(N__13346));
    LocalMux I__2474 (
            .O(N__13368),
            .I(N__13343));
    LocalMux I__2473 (
            .O(N__13365),
            .I(N__13340));
    CascadeMux I__2472 (
            .O(N__13364),
            .I(N__13336));
    InMux I__2471 (
            .O(N__13363),
            .I(N__13333));
    Span4Mux_v I__2470 (
            .O(N__13358),
            .I(N__13328));
    Span4Mux_v I__2469 (
            .O(N__13353),
            .I(N__13328));
    Span4Mux_v I__2468 (
            .O(N__13346),
            .I(N__13325));
    Span4Mux_h I__2467 (
            .O(N__13343),
            .I(N__13320));
    Span4Mux_v I__2466 (
            .O(N__13340),
            .I(N__13320));
    InMux I__2465 (
            .O(N__13339),
            .I(N__13315));
    InMux I__2464 (
            .O(N__13336),
            .I(N__13315));
    LocalMux I__2463 (
            .O(N__13333),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2462 (
            .O(N__13328),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2461 (
            .O(N__13325),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2460 (
            .O(N__13320),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__2459 (
            .O(N__13315),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    InMux I__2458 (
            .O(N__13304),
            .I(N__13297));
    InMux I__2457 (
            .O(N__13303),
            .I(N__13292));
    InMux I__2456 (
            .O(N__13302),
            .I(N__13292));
    InMux I__2455 (
            .O(N__13301),
            .I(N__13289));
    InMux I__2454 (
            .O(N__13300),
            .I(N__13286));
    LocalMux I__2453 (
            .O(N__13297),
            .I(N__13282));
    LocalMux I__2452 (
            .O(N__13292),
            .I(N__13279));
    LocalMux I__2451 (
            .O(N__13289),
            .I(N__13276));
    LocalMux I__2450 (
            .O(N__13286),
            .I(N__13273));
    InMux I__2449 (
            .O(N__13285),
            .I(N__13269));
    Span4Mux_v I__2448 (
            .O(N__13282),
            .I(N__13264));
    Span4Mux_h I__2447 (
            .O(N__13279),
            .I(N__13264));
    Span4Mux_v I__2446 (
            .O(N__13276),
            .I(N__13259));
    Span4Mux_v I__2445 (
            .O(N__13273),
            .I(N__13259));
    InMux I__2444 (
            .O(N__13272),
            .I(N__13256));
    LocalMux I__2443 (
            .O(N__13269),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__2442 (
            .O(N__13264),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__2441 (
            .O(N__13259),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2440 (
            .O(N__13256),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    CascadeMux I__2439 (
            .O(N__13247),
            .I(N__13244));
    InMux I__2438 (
            .O(N__13244),
            .I(N__13241));
    LocalMux I__2437 (
            .O(N__13241),
            .I(N__13238));
    Span4Mux_h I__2436 (
            .O(N__13238),
            .I(N__13235));
    Odrv4 I__2435 (
            .O(N__13235),
            .I(\this_vga_signals.g0_0 ));
    CascadeMux I__2434 (
            .O(N__13232),
            .I(N_206_cascade_));
    InMux I__2433 (
            .O(N__13229),
            .I(N__13226));
    LocalMux I__2432 (
            .O(N__13226),
            .I(N_207));
    InMux I__2431 (
            .O(N__13223),
            .I(N__13220));
    LocalMux I__2430 (
            .O(N__13220),
            .I(M_this_state_q_srsts_0_a2_1_4));
    IoInMux I__2429 (
            .O(N__13217),
            .I(N__13214));
    LocalMux I__2428 (
            .O(N__13214),
            .I(N__13210));
    InMux I__2427 (
            .O(N__13213),
            .I(N__13205));
    IoSpan4Mux I__2426 (
            .O(N__13210),
            .I(N__13202));
    InMux I__2425 (
            .O(N__13209),
            .I(N__13199));
    CascadeMux I__2424 (
            .O(N__13208),
            .I(N__13196));
    LocalMux I__2423 (
            .O(N__13205),
            .I(N__13193));
    Sp12to4 I__2422 (
            .O(N__13202),
            .I(N__13190));
    LocalMux I__2421 (
            .O(N__13199),
            .I(N__13187));
    InMux I__2420 (
            .O(N__13196),
            .I(N__13184));
    Sp12to4 I__2419 (
            .O(N__13193),
            .I(N__13181));
    Span12Mux_h I__2418 (
            .O(N__13190),
            .I(N__13178));
    Span12Mux_v I__2417 (
            .O(N__13187),
            .I(N__13175));
    LocalMux I__2416 (
            .O(N__13184),
            .I(N__13170));
    Span12Mux_v I__2415 (
            .O(N__13181),
            .I(N__13167));
    Span12Mux_v I__2414 (
            .O(N__13178),
            .I(N__13162));
    Span12Mux_h I__2413 (
            .O(N__13175),
            .I(N__13162));
    InMux I__2412 (
            .O(N__13174),
            .I(N__13159));
    InMux I__2411 (
            .O(N__13173),
            .I(N__13156));
    Span4Mux_v I__2410 (
            .O(N__13170),
            .I(N__13153));
    Odrv12 I__2409 (
            .O(N__13167),
            .I(port_dmab_c));
    Odrv12 I__2408 (
            .O(N__13162),
            .I(port_dmab_c));
    LocalMux I__2407 (
            .O(N__13159),
            .I(port_dmab_c));
    LocalMux I__2406 (
            .O(N__13156),
            .I(port_dmab_c));
    Odrv4 I__2405 (
            .O(N__13153),
            .I(port_dmab_c));
    IoInMux I__2404 (
            .O(N__13142),
            .I(N__13138));
    IoInMux I__2403 (
            .O(N__13141),
            .I(N__13135));
    LocalMux I__2402 (
            .O(N__13138),
            .I(N__13130));
    LocalMux I__2401 (
            .O(N__13135),
            .I(N__13130));
    IoSpan4Mux I__2400 (
            .O(N__13130),
            .I(N__13126));
    IoInMux I__2399 (
            .O(N__13129),
            .I(N__13121));
    IoSpan4Mux I__2398 (
            .O(N__13126),
            .I(N__13117));
    IoInMux I__2397 (
            .O(N__13125),
            .I(N__13114));
    IoInMux I__2396 (
            .O(N__13124),
            .I(N__13111));
    LocalMux I__2395 (
            .O(N__13121),
            .I(N__13106));
    IoInMux I__2394 (
            .O(N__13120),
            .I(N__13103));
    IoSpan4Mux I__2393 (
            .O(N__13117),
            .I(N__13092));
    LocalMux I__2392 (
            .O(N__13114),
            .I(N__13092));
    LocalMux I__2391 (
            .O(N__13111),
            .I(N__13092));
    IoInMux I__2390 (
            .O(N__13110),
            .I(N__13089));
    IoInMux I__2389 (
            .O(N__13109),
            .I(N__13086));
    IoSpan4Mux I__2388 (
            .O(N__13106),
            .I(N__13081));
    LocalMux I__2387 (
            .O(N__13103),
            .I(N__13081));
    IoInMux I__2386 (
            .O(N__13102),
            .I(N__13078));
    IoInMux I__2385 (
            .O(N__13101),
            .I(N__13075));
    IoInMux I__2384 (
            .O(N__13100),
            .I(N__13072));
    IoInMux I__2383 (
            .O(N__13099),
            .I(N__13069));
    IoSpan4Mux I__2382 (
            .O(N__13092),
            .I(N__13061));
    LocalMux I__2381 (
            .O(N__13089),
            .I(N__13061));
    LocalMux I__2380 (
            .O(N__13086),
            .I(N__13061));
    IoSpan4Mux I__2379 (
            .O(N__13081),
            .I(N__13056));
    LocalMux I__2378 (
            .O(N__13078),
            .I(N__13056));
    LocalMux I__2377 (
            .O(N__13075),
            .I(N__13053));
    LocalMux I__2376 (
            .O(N__13072),
            .I(N__13049));
    LocalMux I__2375 (
            .O(N__13069),
            .I(N__13046));
    IoInMux I__2374 (
            .O(N__13068),
            .I(N__13043));
    IoSpan4Mux I__2373 (
            .O(N__13061),
            .I(N__13036));
    IoSpan4Mux I__2372 (
            .O(N__13056),
            .I(N__13036));
    Span4Mux_s2_h I__2371 (
            .O(N__13053),
            .I(N__13032));
    IoInMux I__2370 (
            .O(N__13052),
            .I(N__13029));
    IoSpan4Mux I__2369 (
            .O(N__13049),
            .I(N__13022));
    IoSpan4Mux I__2368 (
            .O(N__13046),
            .I(N__13022));
    LocalMux I__2367 (
            .O(N__13043),
            .I(N__13022));
    IoInMux I__2366 (
            .O(N__13042),
            .I(N__13019));
    IoInMux I__2365 (
            .O(N__13041),
            .I(N__13016));
    Span4Mux_s3_h I__2364 (
            .O(N__13036),
            .I(N__13013));
    IoInMux I__2363 (
            .O(N__13035),
            .I(N__13010));
    Span4Mux_h I__2362 (
            .O(N__13032),
            .I(N__13007));
    LocalMux I__2361 (
            .O(N__13029),
            .I(N__13004));
    IoSpan4Mux I__2360 (
            .O(N__13022),
            .I(N__12997));
    LocalMux I__2359 (
            .O(N__13019),
            .I(N__12997));
    LocalMux I__2358 (
            .O(N__13016),
            .I(N__12997));
    Sp12to4 I__2357 (
            .O(N__13013),
            .I(N__12992));
    LocalMux I__2356 (
            .O(N__13010),
            .I(N__12992));
    Span4Mux_h I__2355 (
            .O(N__13007),
            .I(N__12989));
    Span12Mux_s0_v I__2354 (
            .O(N__13004),
            .I(N__12986));
    IoSpan4Mux I__2353 (
            .O(N__12997),
            .I(N__12983));
    Span12Mux_s11_h I__2352 (
            .O(N__12992),
            .I(N__12980));
    Span4Mux_h I__2351 (
            .O(N__12989),
            .I(N__12977));
    Span12Mux_h I__2350 (
            .O(N__12986),
            .I(N__12972));
    Sp12to4 I__2349 (
            .O(N__12983),
            .I(N__12972));
    Odrv12 I__2348 (
            .O(N__12980),
            .I(port_dmab_c_i));
    Odrv4 I__2347 (
            .O(N__12977),
            .I(port_dmab_c_i));
    Odrv12 I__2346 (
            .O(N__12972),
            .I(port_dmab_c_i));
    InMux I__2345 (
            .O(N__12965),
            .I(N__12959));
    CascadeMux I__2344 (
            .O(N__12964),
            .I(N__12954));
    InMux I__2343 (
            .O(N__12963),
            .I(N__12945));
    CascadeMux I__2342 (
            .O(N__12962),
            .I(N__12942));
    LocalMux I__2341 (
            .O(N__12959),
            .I(N__12939));
    InMux I__2340 (
            .O(N__12958),
            .I(N__12936));
    InMux I__2339 (
            .O(N__12957),
            .I(N__12931));
    InMux I__2338 (
            .O(N__12954),
            .I(N__12931));
    InMux I__2337 (
            .O(N__12953),
            .I(N__12926));
    InMux I__2336 (
            .O(N__12952),
            .I(N__12926));
    InMux I__2335 (
            .O(N__12951),
            .I(N__12923));
    InMux I__2334 (
            .O(N__12950),
            .I(N__12920));
    InMux I__2333 (
            .O(N__12949),
            .I(N__12917));
    InMux I__2332 (
            .O(N__12948),
            .I(N__12914));
    LocalMux I__2331 (
            .O(N__12945),
            .I(N__12911));
    InMux I__2330 (
            .O(N__12942),
            .I(N__12908));
    Span4Mux_v I__2329 (
            .O(N__12939),
            .I(N__12901));
    LocalMux I__2328 (
            .O(N__12936),
            .I(N__12901));
    LocalMux I__2327 (
            .O(N__12931),
            .I(N__12901));
    LocalMux I__2326 (
            .O(N__12926),
            .I(N__12898));
    LocalMux I__2325 (
            .O(N__12923),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2324 (
            .O(N__12920),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2323 (
            .O(N__12917),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2322 (
            .O(N__12914),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__2321 (
            .O(N__12911),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2320 (
            .O(N__12908),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__2319 (
            .O(N__12901),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv12 I__2318 (
            .O(N__12898),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    CascadeMux I__2317 (
            .O(N__12881),
            .I(N__12878));
    InMux I__2316 (
            .O(N__12878),
            .I(N__12875));
    LocalMux I__2315 (
            .O(N__12875),
            .I(N__12872));
    Span4Mux_v I__2314 (
            .O(N__12872),
            .I(N__12869));
    Odrv4 I__2313 (
            .O(N__12869),
            .I(\this_vga_signals.g1_0 ));
    InMux I__2312 (
            .O(N__12866),
            .I(N__12863));
    LocalMux I__2311 (
            .O(N__12863),
            .I(N__12859));
    InMux I__2310 (
            .O(N__12862),
            .I(N__12856));
    Span4Mux_v I__2309 (
            .O(N__12859),
            .I(N__12853));
    LocalMux I__2308 (
            .O(N__12856),
            .I(N__12847));
    Span4Mux_h I__2307 (
            .O(N__12853),
            .I(N__12847));
    InMux I__2306 (
            .O(N__12852),
            .I(N__12844));
    Odrv4 I__2305 (
            .O(N__12847),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__2304 (
            .O(N__12844),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    CascadeMux I__2303 (
            .O(N__12839),
            .I(N__12833));
    CascadeMux I__2302 (
            .O(N__12838),
            .I(N__12829));
    CascadeMux I__2301 (
            .O(N__12837),
            .I(N__12823));
    InMux I__2300 (
            .O(N__12836),
            .I(N__12820));
    InMux I__2299 (
            .O(N__12833),
            .I(N__12813));
    InMux I__2298 (
            .O(N__12832),
            .I(N__12803));
    InMux I__2297 (
            .O(N__12829),
            .I(N__12794));
    InMux I__2296 (
            .O(N__12828),
            .I(N__12794));
    InMux I__2295 (
            .O(N__12827),
            .I(N__12794));
    InMux I__2294 (
            .O(N__12826),
            .I(N__12794));
    InMux I__2293 (
            .O(N__12823),
            .I(N__12790));
    LocalMux I__2292 (
            .O(N__12820),
            .I(N__12787));
    InMux I__2291 (
            .O(N__12819),
            .I(N__12784));
    InMux I__2290 (
            .O(N__12818),
            .I(N__12781));
    InMux I__2289 (
            .O(N__12817),
            .I(N__12778));
    CascadeMux I__2288 (
            .O(N__12816),
            .I(N__12770));
    LocalMux I__2287 (
            .O(N__12813),
            .I(N__12766));
    InMux I__2286 (
            .O(N__12812),
            .I(N__12763));
    InMux I__2285 (
            .O(N__12811),
            .I(N__12760));
    InMux I__2284 (
            .O(N__12810),
            .I(N__12749));
    InMux I__2283 (
            .O(N__12809),
            .I(N__12749));
    InMux I__2282 (
            .O(N__12808),
            .I(N__12749));
    InMux I__2281 (
            .O(N__12807),
            .I(N__12749));
    InMux I__2280 (
            .O(N__12806),
            .I(N__12749));
    LocalMux I__2279 (
            .O(N__12803),
            .I(N__12746));
    LocalMux I__2278 (
            .O(N__12794),
            .I(N__12743));
    InMux I__2277 (
            .O(N__12793),
            .I(N__12740));
    LocalMux I__2276 (
            .O(N__12790),
            .I(N__12729));
    Span4Mux_v I__2275 (
            .O(N__12787),
            .I(N__12729));
    LocalMux I__2274 (
            .O(N__12784),
            .I(N__12729));
    LocalMux I__2273 (
            .O(N__12781),
            .I(N__12729));
    LocalMux I__2272 (
            .O(N__12778),
            .I(N__12729));
    InMux I__2271 (
            .O(N__12777),
            .I(N__12725));
    InMux I__2270 (
            .O(N__12776),
            .I(N__12720));
    InMux I__2269 (
            .O(N__12775),
            .I(N__12720));
    InMux I__2268 (
            .O(N__12774),
            .I(N__12711));
    InMux I__2267 (
            .O(N__12773),
            .I(N__12711));
    InMux I__2266 (
            .O(N__12770),
            .I(N__12711));
    InMux I__2265 (
            .O(N__12769),
            .I(N__12711));
    Span4Mux_v I__2264 (
            .O(N__12766),
            .I(N__12701));
    LocalMux I__2263 (
            .O(N__12763),
            .I(N__12701));
    LocalMux I__2262 (
            .O(N__12760),
            .I(N__12701));
    LocalMux I__2261 (
            .O(N__12749),
            .I(N__12701));
    Span4Mux_v I__2260 (
            .O(N__12746),
            .I(N__12692));
    Span4Mux_v I__2259 (
            .O(N__12743),
            .I(N__12692));
    LocalMux I__2258 (
            .O(N__12740),
            .I(N__12692));
    Span4Mux_v I__2257 (
            .O(N__12729),
            .I(N__12692));
    InMux I__2256 (
            .O(N__12728),
            .I(N__12689));
    LocalMux I__2255 (
            .O(N__12725),
            .I(N__12682));
    LocalMux I__2254 (
            .O(N__12720),
            .I(N__12682));
    LocalMux I__2253 (
            .O(N__12711),
            .I(N__12682));
    InMux I__2252 (
            .O(N__12710),
            .I(N__12677));
    Span4Mux_v I__2251 (
            .O(N__12701),
            .I(N__12674));
    Span4Mux_h I__2250 (
            .O(N__12692),
            .I(N__12671));
    LocalMux I__2249 (
            .O(N__12689),
            .I(N__12666));
    Span4Mux_h I__2248 (
            .O(N__12682),
            .I(N__12666));
    InMux I__2247 (
            .O(N__12681),
            .I(N__12661));
    InMux I__2246 (
            .O(N__12680),
            .I(N__12661));
    LocalMux I__2245 (
            .O(N__12677),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2244 (
            .O(N__12674),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2243 (
            .O(N__12671),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2242 (
            .O(N__12666),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2241 (
            .O(N__12661),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    InMux I__2240 (
            .O(N__12650),
            .I(N__12636));
    CascadeMux I__2239 (
            .O(N__12649),
            .I(N__12632));
    InMux I__2238 (
            .O(N__12648),
            .I(N__12629));
    InMux I__2237 (
            .O(N__12647),
            .I(N__12626));
    CascadeMux I__2236 (
            .O(N__12646),
            .I(N__12620));
    InMux I__2235 (
            .O(N__12645),
            .I(N__12614));
    CascadeMux I__2234 (
            .O(N__12644),
            .I(N__12611));
    CascadeMux I__2233 (
            .O(N__12643),
            .I(N__12606));
    CascadeMux I__2232 (
            .O(N__12642),
            .I(N__12603));
    CascadeMux I__2231 (
            .O(N__12641),
            .I(N__12597));
    CascadeMux I__2230 (
            .O(N__12640),
            .I(N__12592));
    InMux I__2229 (
            .O(N__12639),
            .I(N__12587));
    LocalMux I__2228 (
            .O(N__12636),
            .I(N__12584));
    InMux I__2227 (
            .O(N__12635),
            .I(N__12579));
    InMux I__2226 (
            .O(N__12632),
            .I(N__12579));
    LocalMux I__2225 (
            .O(N__12629),
            .I(N__12576));
    LocalMux I__2224 (
            .O(N__12626),
            .I(N__12573));
    InMux I__2223 (
            .O(N__12625),
            .I(N__12570));
    InMux I__2222 (
            .O(N__12624),
            .I(N__12567));
    InMux I__2221 (
            .O(N__12623),
            .I(N__12564));
    InMux I__2220 (
            .O(N__12620),
            .I(N__12559));
    InMux I__2219 (
            .O(N__12619),
            .I(N__12559));
    InMux I__2218 (
            .O(N__12618),
            .I(N__12554));
    InMux I__2217 (
            .O(N__12617),
            .I(N__12554));
    LocalMux I__2216 (
            .O(N__12614),
            .I(N__12551));
    InMux I__2215 (
            .O(N__12611),
            .I(N__12546));
    InMux I__2214 (
            .O(N__12610),
            .I(N__12546));
    CascadeMux I__2213 (
            .O(N__12609),
            .I(N__12542));
    InMux I__2212 (
            .O(N__12606),
            .I(N__12535));
    InMux I__2211 (
            .O(N__12603),
            .I(N__12535));
    InMux I__2210 (
            .O(N__12602),
            .I(N__12535));
    InMux I__2209 (
            .O(N__12601),
            .I(N__12532));
    InMux I__2208 (
            .O(N__12600),
            .I(N__12528));
    InMux I__2207 (
            .O(N__12597),
            .I(N__12525));
    InMux I__2206 (
            .O(N__12596),
            .I(N__12516));
    InMux I__2205 (
            .O(N__12595),
            .I(N__12516));
    InMux I__2204 (
            .O(N__12592),
            .I(N__12516));
    InMux I__2203 (
            .O(N__12591),
            .I(N__12516));
    InMux I__2202 (
            .O(N__12590),
            .I(N__12513));
    LocalMux I__2201 (
            .O(N__12587),
            .I(N__12510));
    Span4Mux_v I__2200 (
            .O(N__12584),
            .I(N__12505));
    LocalMux I__2199 (
            .O(N__12579),
            .I(N__12505));
    Span4Mux_v I__2198 (
            .O(N__12576),
            .I(N__12498));
    Span4Mux_v I__2197 (
            .O(N__12573),
            .I(N__12498));
    LocalMux I__2196 (
            .O(N__12570),
            .I(N__12483));
    LocalMux I__2195 (
            .O(N__12567),
            .I(N__12483));
    LocalMux I__2194 (
            .O(N__12564),
            .I(N__12483));
    LocalMux I__2193 (
            .O(N__12559),
            .I(N__12483));
    LocalMux I__2192 (
            .O(N__12554),
            .I(N__12483));
    Span4Mux_v I__2191 (
            .O(N__12551),
            .I(N__12483));
    LocalMux I__2190 (
            .O(N__12546),
            .I(N__12483));
    InMux I__2189 (
            .O(N__12545),
            .I(N__12480));
    InMux I__2188 (
            .O(N__12542),
            .I(N__12477));
    LocalMux I__2187 (
            .O(N__12535),
            .I(N__12472));
    LocalMux I__2186 (
            .O(N__12532),
            .I(N__12472));
    InMux I__2185 (
            .O(N__12531),
            .I(N__12469));
    LocalMux I__2184 (
            .O(N__12528),
            .I(N__12460));
    LocalMux I__2183 (
            .O(N__12525),
            .I(N__12460));
    LocalMux I__2182 (
            .O(N__12516),
            .I(N__12460));
    LocalMux I__2181 (
            .O(N__12513),
            .I(N__12460));
    Span4Mux_h I__2180 (
            .O(N__12510),
            .I(N__12455));
    Span4Mux_v I__2179 (
            .O(N__12505),
            .I(N__12455));
    InMux I__2178 (
            .O(N__12504),
            .I(N__12450));
    InMux I__2177 (
            .O(N__12503),
            .I(N__12450));
    Span4Mux_h I__2176 (
            .O(N__12498),
            .I(N__12445));
    Span4Mux_v I__2175 (
            .O(N__12483),
            .I(N__12445));
    LocalMux I__2174 (
            .O(N__12480),
            .I(N__12438));
    LocalMux I__2173 (
            .O(N__12477),
            .I(N__12438));
    Span4Mux_v I__2172 (
            .O(N__12472),
            .I(N__12438));
    LocalMux I__2171 (
            .O(N__12469),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv12 I__2170 (
            .O(N__12460),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2169 (
            .O(N__12455),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2168 (
            .O(N__12450),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2167 (
            .O(N__12445),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2166 (
            .O(N__12438),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    CascadeMux I__2165 (
            .O(N__12425),
            .I(N__12422));
    InMux I__2164 (
            .O(N__12422),
            .I(N__12415));
    CascadeMux I__2163 (
            .O(N__12421),
            .I(N__12410));
    InMux I__2162 (
            .O(N__12420),
            .I(N__12405));
    InMux I__2161 (
            .O(N__12419),
            .I(N__12402));
    InMux I__2160 (
            .O(N__12418),
            .I(N__12396));
    LocalMux I__2159 (
            .O(N__12415),
            .I(N__12393));
    InMux I__2158 (
            .O(N__12414),
            .I(N__12390));
    InMux I__2157 (
            .O(N__12413),
            .I(N__12387));
    InMux I__2156 (
            .O(N__12410),
            .I(N__12380));
    InMux I__2155 (
            .O(N__12409),
            .I(N__12380));
    CascadeMux I__2154 (
            .O(N__12408),
            .I(N__12376));
    LocalMux I__2153 (
            .O(N__12405),
            .I(N__12373));
    LocalMux I__2152 (
            .O(N__12402),
            .I(N__12370));
    InMux I__2151 (
            .O(N__12401),
            .I(N__12363));
    InMux I__2150 (
            .O(N__12400),
            .I(N__12363));
    InMux I__2149 (
            .O(N__12399),
            .I(N__12363));
    LocalMux I__2148 (
            .O(N__12396),
            .I(N__12358));
    Span4Mux_v I__2147 (
            .O(N__12393),
            .I(N__12351));
    LocalMux I__2146 (
            .O(N__12390),
            .I(N__12351));
    LocalMux I__2145 (
            .O(N__12387),
            .I(N__12351));
    InMux I__2144 (
            .O(N__12386),
            .I(N__12346));
    InMux I__2143 (
            .O(N__12385),
            .I(N__12346));
    LocalMux I__2142 (
            .O(N__12380),
            .I(N__12343));
    CascadeMux I__2141 (
            .O(N__12379),
            .I(N__12335));
    InMux I__2140 (
            .O(N__12376),
            .I(N__12331));
    Span4Mux_v I__2139 (
            .O(N__12373),
            .I(N__12326));
    Span4Mux_v I__2138 (
            .O(N__12370),
            .I(N__12326));
    LocalMux I__2137 (
            .O(N__12363),
            .I(N__12323));
    InMux I__2136 (
            .O(N__12362),
            .I(N__12318));
    InMux I__2135 (
            .O(N__12361),
            .I(N__12318));
    Span4Mux_h I__2134 (
            .O(N__12358),
            .I(N__12309));
    Span4Mux_h I__2133 (
            .O(N__12351),
            .I(N__12309));
    LocalMux I__2132 (
            .O(N__12346),
            .I(N__12309));
    Span4Mux_h I__2131 (
            .O(N__12343),
            .I(N__12309));
    InMux I__2130 (
            .O(N__12342),
            .I(N__12298));
    InMux I__2129 (
            .O(N__12341),
            .I(N__12298));
    InMux I__2128 (
            .O(N__12340),
            .I(N__12298));
    InMux I__2127 (
            .O(N__12339),
            .I(N__12298));
    InMux I__2126 (
            .O(N__12338),
            .I(N__12298));
    InMux I__2125 (
            .O(N__12335),
            .I(N__12293));
    InMux I__2124 (
            .O(N__12334),
            .I(N__12293));
    LocalMux I__2123 (
            .O(N__12331),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2122 (
            .O(N__12326),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv12 I__2121 (
            .O(N__12323),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2120 (
            .O(N__12318),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2119 (
            .O(N__12309),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2118 (
            .O(N__12298),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2117 (
            .O(N__12293),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    InMux I__2116 (
            .O(N__12278),
            .I(N__12274));
    CascadeMux I__2115 (
            .O(N__12277),
            .I(N__12271));
    LocalMux I__2114 (
            .O(N__12274),
            .I(N__12268));
    InMux I__2113 (
            .O(N__12271),
            .I(N__12265));
    Span4Mux_h I__2112 (
            .O(N__12268),
            .I(N__12262));
    LocalMux I__2111 (
            .O(N__12265),
            .I(\this_vga_signals.M_vcounter_d7lt8_0 ));
    Odrv4 I__2110 (
            .O(N__12262),
            .I(\this_vga_signals.M_vcounter_d7lt8_0 ));
    CascadeMux I__2109 (
            .O(N__12257),
            .I(N__12250));
    CascadeMux I__2108 (
            .O(N__12256),
            .I(N__12243));
    CascadeMux I__2107 (
            .O(N__12255),
            .I(N__12239));
    InMux I__2106 (
            .O(N__12254),
            .I(N__12236));
    InMux I__2105 (
            .O(N__12253),
            .I(N__12231));
    InMux I__2104 (
            .O(N__12250),
            .I(N__12231));
    CascadeMux I__2103 (
            .O(N__12249),
            .I(N__12228));
    InMux I__2102 (
            .O(N__12248),
            .I(N__12225));
    InMux I__2101 (
            .O(N__12247),
            .I(N__12220));
    InMux I__2100 (
            .O(N__12246),
            .I(N__12220));
    InMux I__2099 (
            .O(N__12243),
            .I(N__12215));
    InMux I__2098 (
            .O(N__12242),
            .I(N__12212));
    InMux I__2097 (
            .O(N__12239),
            .I(N__12206));
    LocalMux I__2096 (
            .O(N__12236),
            .I(N__12203));
    LocalMux I__2095 (
            .O(N__12231),
            .I(N__12200));
    InMux I__2094 (
            .O(N__12228),
            .I(N__12197));
    LocalMux I__2093 (
            .O(N__12225),
            .I(N__12192));
    LocalMux I__2092 (
            .O(N__12220),
            .I(N__12192));
    InMux I__2091 (
            .O(N__12219),
            .I(N__12187));
    InMux I__2090 (
            .O(N__12218),
            .I(N__12187));
    LocalMux I__2089 (
            .O(N__12215),
            .I(N__12180));
    LocalMux I__2088 (
            .O(N__12212),
            .I(N__12177));
    InMux I__2087 (
            .O(N__12211),
            .I(N__12174));
    InMux I__2086 (
            .O(N__12210),
            .I(N__12169));
    InMux I__2085 (
            .O(N__12209),
            .I(N__12169));
    LocalMux I__2084 (
            .O(N__12206),
            .I(N__12164));
    Span4Mux_v I__2083 (
            .O(N__12203),
            .I(N__12164));
    Span4Mux_v I__2082 (
            .O(N__12200),
            .I(N__12157));
    LocalMux I__2081 (
            .O(N__12197),
            .I(N__12157));
    Span4Mux_v I__2080 (
            .O(N__12192),
            .I(N__12157));
    LocalMux I__2079 (
            .O(N__12187),
            .I(N__12154));
    InMux I__2078 (
            .O(N__12186),
            .I(N__12149));
    InMux I__2077 (
            .O(N__12185),
            .I(N__12149));
    InMux I__2076 (
            .O(N__12184),
            .I(N__12144));
    InMux I__2075 (
            .O(N__12183),
            .I(N__12144));
    Odrv4 I__2074 (
            .O(N__12180),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2073 (
            .O(N__12177),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2072 (
            .O(N__12174),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2071 (
            .O(N__12169),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2070 (
            .O(N__12164),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2069 (
            .O(N__12157),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2068 (
            .O(N__12154),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2067 (
            .O(N__12149),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2066 (
            .O(N__12144),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    CascadeMux I__2065 (
            .O(N__12125),
            .I(\this_vga_signals.un4_lvisibility_1_cascade_ ));
    InMux I__2064 (
            .O(N__12122),
            .I(N__12119));
    LocalMux I__2063 (
            .O(N__12119),
            .I(N__12113));
    InMux I__2062 (
            .O(N__12118),
            .I(N__12107));
    CascadeMux I__2061 (
            .O(N__12117),
            .I(N__12104));
    CascadeMux I__2060 (
            .O(N__12116),
            .I(N__12101));
    Span4Mux_v I__2059 (
            .O(N__12113),
            .I(N__12098));
    InMux I__2058 (
            .O(N__12112),
            .I(N__12095));
    InMux I__2057 (
            .O(N__12111),
            .I(N__12090));
    InMux I__2056 (
            .O(N__12110),
            .I(N__12090));
    LocalMux I__2055 (
            .O(N__12107),
            .I(N__12087));
    InMux I__2054 (
            .O(N__12104),
            .I(N__12084));
    InMux I__2053 (
            .O(N__12101),
            .I(N__12081));
    Odrv4 I__2052 (
            .O(N__12098),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2051 (
            .O(N__12095),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2050 (
            .O(N__12090),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2049 (
            .O(N__12087),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2048 (
            .O(N__12084),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2047 (
            .O(N__12081),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    InMux I__2046 (
            .O(N__12068),
            .I(N__12062));
    InMux I__2045 (
            .O(N__12067),
            .I(N__12062));
    LocalMux I__2044 (
            .O(N__12062),
            .I(\this_vga_signals.line_clk_1 ));
    CascadeMux I__2043 (
            .O(N__12059),
            .I(N__12056));
    InMux I__2042 (
            .O(N__12056),
            .I(N__12053));
    LocalMux I__2041 (
            .O(N__12053),
            .I(\this_vga_signals.un4_lvisibility_1 ));
    InMux I__2040 (
            .O(N__12050),
            .I(N__12043));
    InMux I__2039 (
            .O(N__12049),
            .I(N__12040));
    InMux I__2038 (
            .O(N__12048),
            .I(N__12035));
    InMux I__2037 (
            .O(N__12047),
            .I(N__12032));
    InMux I__2036 (
            .O(N__12046),
            .I(N__12029));
    LocalMux I__2035 (
            .O(N__12043),
            .I(N__12024));
    LocalMux I__2034 (
            .O(N__12040),
            .I(N__12024));
    InMux I__2033 (
            .O(N__12039),
            .I(N__12020));
    CascadeMux I__2032 (
            .O(N__12038),
            .I(N__12016));
    LocalMux I__2031 (
            .O(N__12035),
            .I(N__12013));
    LocalMux I__2030 (
            .O(N__12032),
            .I(N__12010));
    LocalMux I__2029 (
            .O(N__12029),
            .I(N__12005));
    Span4Mux_v I__2028 (
            .O(N__12024),
            .I(N__12005));
    InMux I__2027 (
            .O(N__12023),
            .I(N__12002));
    LocalMux I__2026 (
            .O(N__12020),
            .I(N__11999));
    InMux I__2025 (
            .O(N__12019),
            .I(N__11994));
    InMux I__2024 (
            .O(N__12016),
            .I(N__11994));
    Span4Mux_h I__2023 (
            .O(N__12013),
            .I(N__11991));
    Odrv12 I__2022 (
            .O(N__12010),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2021 (
            .O(N__12005),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2020 (
            .O(N__12002),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2019 (
            .O(N__11999),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2018 (
            .O(N__11994),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2017 (
            .O(N__11991),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    CascadeMux I__2016 (
            .O(N__11978),
            .I(N__11974));
    InMux I__2015 (
            .O(N__11977),
            .I(N__11971));
    InMux I__2014 (
            .O(N__11974),
            .I(N__11968));
    LocalMux I__2013 (
            .O(N__11971),
            .I(N__11965));
    LocalMux I__2012 (
            .O(N__11968),
            .I(N__11960));
    Span4Mux_h I__2011 (
            .O(N__11965),
            .I(N__11957));
    InMux I__2010 (
            .O(N__11964),
            .I(N__11954));
    InMux I__2009 (
            .O(N__11963),
            .I(N__11951));
    Span4Mux_h I__2008 (
            .O(N__11960),
            .I(N__11946));
    Span4Mux_h I__2007 (
            .O(N__11957),
            .I(N__11946));
    LocalMux I__2006 (
            .O(N__11954),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__2005 (
            .O(N__11951),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    Odrv4 I__2004 (
            .O(N__11946),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    CascadeMux I__2003 (
            .O(N__11939),
            .I(N__11932));
    InMux I__2002 (
            .O(N__11938),
            .I(N__11927));
    InMux I__2001 (
            .O(N__11937),
            .I(N__11924));
    InMux I__2000 (
            .O(N__11936),
            .I(N__11919));
    InMux I__1999 (
            .O(N__11935),
            .I(N__11919));
    InMux I__1998 (
            .O(N__11932),
            .I(N__11914));
    InMux I__1997 (
            .O(N__11931),
            .I(N__11914));
    InMux I__1996 (
            .O(N__11930),
            .I(N__11911));
    LocalMux I__1995 (
            .O(N__11927),
            .I(N__11906));
    LocalMux I__1994 (
            .O(N__11924),
            .I(N__11906));
    LocalMux I__1993 (
            .O(N__11919),
            .I(N__11901));
    LocalMux I__1992 (
            .O(N__11914),
            .I(N__11901));
    LocalMux I__1991 (
            .O(N__11911),
            .I(N__11897));
    Span4Mux_v I__1990 (
            .O(N__11906),
            .I(N__11894));
    Span4Mux_v I__1989 (
            .O(N__11901),
            .I(N__11891));
    InMux I__1988 (
            .O(N__11900),
            .I(N__11888));
    Span4Mux_v I__1987 (
            .O(N__11897),
            .I(N__11881));
    Span4Mux_h I__1986 (
            .O(N__11894),
            .I(N__11881));
    Span4Mux_h I__1985 (
            .O(N__11891),
            .I(N__11881));
    LocalMux I__1984 (
            .O(N__11888),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__1983 (
            .O(N__11881),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    InMux I__1982 (
            .O(N__11876),
            .I(N__11873));
    LocalMux I__1981 (
            .O(N__11873),
            .I(N__11870));
    Span4Mux_h I__1980 (
            .O(N__11870),
            .I(N__11867));
    Span4Mux_h I__1979 (
            .O(N__11867),
            .I(N__11864));
    Odrv4 I__1978 (
            .O(N__11864),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    InMux I__1977 (
            .O(N__11861),
            .I(N__11858));
    LocalMux I__1976 (
            .O(N__11858),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    InMux I__1975 (
            .O(N__11855),
            .I(N__11846));
    InMux I__1974 (
            .O(N__11854),
            .I(N__11846));
    InMux I__1973 (
            .O(N__11853),
            .I(N__11846));
    LocalMux I__1972 (
            .O(N__11846),
            .I(M_this_delay_clk_out_0));
    InMux I__1971 (
            .O(N__11843),
            .I(N__11834));
    InMux I__1970 (
            .O(N__11842),
            .I(N__11834));
    InMux I__1969 (
            .O(N__11841),
            .I(N__11834));
    LocalMux I__1968 (
            .O(N__11834),
            .I(N__11831));
    Sp12to4 I__1967 (
            .O(N__11831),
            .I(N__11828));
    Span12Mux_v I__1966 (
            .O(N__11828),
            .I(N__11825));
    Span12Mux_h I__1965 (
            .O(N__11825),
            .I(N__11822));
    Odrv12 I__1964 (
            .O(N__11822),
            .I(port_enb_c));
    CascadeMux I__1963 (
            .O(N__11819),
            .I(N__11816));
    InMux I__1962 (
            .O(N__11816),
            .I(N__11810));
    InMux I__1961 (
            .O(N__11815),
            .I(N__11810));
    LocalMux I__1960 (
            .O(N__11810),
            .I(this_start_data_delay_M_last_q));
    InMux I__1959 (
            .O(N__11807),
            .I(N__11803));
    InMux I__1958 (
            .O(N__11806),
            .I(N__11800));
    LocalMux I__1957 (
            .O(N__11803),
            .I(N__11797));
    LocalMux I__1956 (
            .O(N__11800),
            .I(N__11794));
    Odrv4 I__1955 (
            .O(N__11797),
            .I(\this_vga_signals.vaddress_ac0_9_0_a0_0 ));
    Odrv4 I__1954 (
            .O(N__11794),
            .I(\this_vga_signals.vaddress_ac0_9_0_a0_0 ));
    InMux I__1953 (
            .O(N__11789),
            .I(N__11786));
    LocalMux I__1952 (
            .O(N__11786),
            .I(N__11783));
    Odrv4 I__1951 (
            .O(N__11783),
            .I(\this_vga_signals.un6_vvisibilitylt9_0 ));
    InMux I__1950 (
            .O(N__11780),
            .I(N__11777));
    LocalMux I__1949 (
            .O(N__11777),
            .I(N__11773));
    InMux I__1948 (
            .O(N__11776),
            .I(N__11770));
    Span4Mux_h I__1947 (
            .O(N__11773),
            .I(N__11764));
    LocalMux I__1946 (
            .O(N__11770),
            .I(N__11764));
    InMux I__1945 (
            .O(N__11769),
            .I(N__11761));
    Odrv4 I__1944 (
            .O(N__11764),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__1943 (
            .O(N__11761),
            .I(\this_vga_signals.vaddress_c2 ));
    InMux I__1942 (
            .O(N__11756),
            .I(N__11753));
    LocalMux I__1941 (
            .O(N__11753),
            .I(N__11749));
    InMux I__1940 (
            .O(N__11752),
            .I(N__11745));
    Span4Mux_h I__1939 (
            .O(N__11749),
            .I(N__11742));
    InMux I__1938 (
            .O(N__11748),
            .I(N__11739));
    LocalMux I__1937 (
            .O(N__11745),
            .I(N__11736));
    Odrv4 I__1936 (
            .O(N__11742),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    LocalMux I__1935 (
            .O(N__11739),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    Odrv12 I__1934 (
            .O(N__11736),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    InMux I__1933 (
            .O(N__11729),
            .I(N__11724));
    InMux I__1932 (
            .O(N__11728),
            .I(N__11721));
    InMux I__1931 (
            .O(N__11727),
            .I(N__11718));
    LocalMux I__1930 (
            .O(N__11724),
            .I(N__11715));
    LocalMux I__1929 (
            .O(N__11721),
            .I(N__11712));
    LocalMux I__1928 (
            .O(N__11718),
            .I(N__11709));
    Span4Mux_h I__1927 (
            .O(N__11715),
            .I(N__11706));
    Span4Mux_h I__1926 (
            .O(N__11712),
            .I(N__11703));
    Span4Mux_h I__1925 (
            .O(N__11709),
            .I(N__11700));
    Odrv4 I__1924 (
            .O(N__11706),
            .I(\this_vga_signals.vaddress_5_6 ));
    Odrv4 I__1923 (
            .O(N__11703),
            .I(\this_vga_signals.vaddress_5_6 ));
    Odrv4 I__1922 (
            .O(N__11700),
            .I(\this_vga_signals.vaddress_5_6 ));
    InMux I__1921 (
            .O(N__11693),
            .I(N__11690));
    LocalMux I__1920 (
            .O(N__11690),
            .I(N__11685));
    InMux I__1919 (
            .O(N__11689),
            .I(N__11682));
    InMux I__1918 (
            .O(N__11688),
            .I(N__11678));
    Span4Mux_v I__1917 (
            .O(N__11685),
            .I(N__11675));
    LocalMux I__1916 (
            .O(N__11682),
            .I(N__11672));
    InMux I__1915 (
            .O(N__11681),
            .I(N__11669));
    LocalMux I__1914 (
            .O(N__11678),
            .I(N__11666));
    Odrv4 I__1913 (
            .O(N__11675),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    Odrv12 I__1912 (
            .O(N__11672),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    LocalMux I__1911 (
            .O(N__11669),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    Odrv4 I__1910 (
            .O(N__11666),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    CascadeMux I__1909 (
            .O(N__11657),
            .I(N__11653));
    InMux I__1908 (
            .O(N__11656),
            .I(N__11650));
    InMux I__1907 (
            .O(N__11653),
            .I(N__11647));
    LocalMux I__1906 (
            .O(N__11650),
            .I(N__11644));
    LocalMux I__1905 (
            .O(N__11647),
            .I(N__11641));
    Span4Mux_h I__1904 (
            .O(N__11644),
            .I(N__11638));
    Span4Mux_h I__1903 (
            .O(N__11641),
            .I(N__11635));
    Odrv4 I__1902 (
            .O(N__11638),
            .I(\this_vga_signals.vaddress_3_5 ));
    Odrv4 I__1901 (
            .O(N__11635),
            .I(\this_vga_signals.vaddress_3_5 ));
    InMux I__1900 (
            .O(N__11630),
            .I(N__11627));
    LocalMux I__1899 (
            .O(N__11627),
            .I(N__11623));
    InMux I__1898 (
            .O(N__11626),
            .I(N__11620));
    Span4Mux_h I__1897 (
            .O(N__11623),
            .I(N__11615));
    LocalMux I__1896 (
            .O(N__11620),
            .I(N__11615));
    Span4Mux_v I__1895 (
            .O(N__11615),
            .I(N__11611));
    InMux I__1894 (
            .O(N__11614),
            .I(N__11608));
    Span4Mux_h I__1893 (
            .O(N__11611),
            .I(N__11605));
    LocalMux I__1892 (
            .O(N__11608),
            .I(N__11602));
    Odrv4 I__1891 (
            .O(N__11605),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    Odrv4 I__1890 (
            .O(N__11602),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    CEMux I__1889 (
            .O(N__11597),
            .I(N__11573));
    CEMux I__1888 (
            .O(N__11596),
            .I(N__11573));
    CEMux I__1887 (
            .O(N__11595),
            .I(N__11573));
    CEMux I__1886 (
            .O(N__11594),
            .I(N__11573));
    CEMux I__1885 (
            .O(N__11593),
            .I(N__11573));
    CEMux I__1884 (
            .O(N__11592),
            .I(N__11573));
    CEMux I__1883 (
            .O(N__11591),
            .I(N__11573));
    CEMux I__1882 (
            .O(N__11590),
            .I(N__11573));
    GlobalMux I__1881 (
            .O(N__11573),
            .I(N__11570));
    gio2CtrlBuf I__1880 (
            .O(N__11570),
            .I(\this_vga_signals.N_340_0_g ));
    InMux I__1879 (
            .O(N__11567),
            .I(N__11564));
    LocalMux I__1878 (
            .O(N__11564),
            .I(N__11552));
    SRMux I__1877 (
            .O(N__11563),
            .I(N__11531));
    SRMux I__1876 (
            .O(N__11562),
            .I(N__11531));
    SRMux I__1875 (
            .O(N__11561),
            .I(N__11531));
    SRMux I__1874 (
            .O(N__11560),
            .I(N__11531));
    SRMux I__1873 (
            .O(N__11559),
            .I(N__11531));
    SRMux I__1872 (
            .O(N__11558),
            .I(N__11531));
    SRMux I__1871 (
            .O(N__11557),
            .I(N__11531));
    SRMux I__1870 (
            .O(N__11556),
            .I(N__11531));
    SRMux I__1869 (
            .O(N__11555),
            .I(N__11531));
    Glb2LocalMux I__1868 (
            .O(N__11552),
            .I(N__11531));
    GlobalMux I__1867 (
            .O(N__11531),
            .I(N__11528));
    gio2CtrlBuf I__1866 (
            .O(N__11528),
            .I(\this_vga_signals.N_515_g ));
    CascadeMux I__1865 (
            .O(N__11525),
            .I(N__11522));
    InMux I__1864 (
            .O(N__11522),
            .I(N__11516));
    InMux I__1863 (
            .O(N__11521),
            .I(N__11513));
    CascadeMux I__1862 (
            .O(N__11520),
            .I(N__11509));
    InMux I__1861 (
            .O(N__11519),
            .I(N__11505));
    LocalMux I__1860 (
            .O(N__11516),
            .I(N__11500));
    LocalMux I__1859 (
            .O(N__11513),
            .I(N__11500));
    InMux I__1858 (
            .O(N__11512),
            .I(N__11497));
    InMux I__1857 (
            .O(N__11509),
            .I(N__11492));
    InMux I__1856 (
            .O(N__11508),
            .I(N__11492));
    LocalMux I__1855 (
            .O(N__11505),
            .I(N__11481));
    Span4Mux_h I__1854 (
            .O(N__11500),
            .I(N__11481));
    LocalMux I__1853 (
            .O(N__11497),
            .I(N__11476));
    LocalMux I__1852 (
            .O(N__11492),
            .I(N__11476));
    InMux I__1851 (
            .O(N__11491),
            .I(N__11469));
    InMux I__1850 (
            .O(N__11490),
            .I(N__11469));
    InMux I__1849 (
            .O(N__11489),
            .I(N__11469));
    InMux I__1848 (
            .O(N__11488),
            .I(N__11462));
    InMux I__1847 (
            .O(N__11487),
            .I(N__11462));
    InMux I__1846 (
            .O(N__11486),
            .I(N__11462));
    Odrv4 I__1845 (
            .O(N__11481),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv12 I__1844 (
            .O(N__11476),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__1843 (
            .O(N__11469),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__1842 (
            .O(N__11462),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    InMux I__1841 (
            .O(N__11453),
            .I(N__11445));
    InMux I__1840 (
            .O(N__11452),
            .I(N__11442));
    InMux I__1839 (
            .O(N__11451),
            .I(N__11433));
    InMux I__1838 (
            .O(N__11450),
            .I(N__11433));
    InMux I__1837 (
            .O(N__11449),
            .I(N__11433));
    InMux I__1836 (
            .O(N__11448),
            .I(N__11433));
    LocalMux I__1835 (
            .O(N__11445),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__1834 (
            .O(N__11442),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__1833 (
            .O(N__11433),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    InMux I__1832 (
            .O(N__11426),
            .I(N__11419));
    InMux I__1831 (
            .O(N__11425),
            .I(N__11416));
    InMux I__1830 (
            .O(N__11424),
            .I(N__11409));
    InMux I__1829 (
            .O(N__11423),
            .I(N__11409));
    InMux I__1828 (
            .O(N__11422),
            .I(N__11409));
    LocalMux I__1827 (
            .O(N__11419),
            .I(N__11406));
    LocalMux I__1826 (
            .O(N__11416),
            .I(N__11401));
    LocalMux I__1825 (
            .O(N__11409),
            .I(N__11401));
    Span4Mux_h I__1824 (
            .O(N__11406),
            .I(N__11398));
    Odrv4 I__1823 (
            .O(N__11401),
            .I(\this_vga_signals.vaddress_5 ));
    Odrv4 I__1822 (
            .O(N__11398),
            .I(\this_vga_signals.vaddress_5 ));
    CascadeMux I__1821 (
            .O(N__11393),
            .I(N__11384));
    InMux I__1820 (
            .O(N__11392),
            .I(N__11381));
    InMux I__1819 (
            .O(N__11391),
            .I(N__11372));
    InMux I__1818 (
            .O(N__11390),
            .I(N__11372));
    InMux I__1817 (
            .O(N__11389),
            .I(N__11372));
    InMux I__1816 (
            .O(N__11388),
            .I(N__11367));
    InMux I__1815 (
            .O(N__11387),
            .I(N__11367));
    InMux I__1814 (
            .O(N__11384),
            .I(N__11364));
    LocalMux I__1813 (
            .O(N__11381),
            .I(N__11361));
    InMux I__1812 (
            .O(N__11380),
            .I(N__11353));
    InMux I__1811 (
            .O(N__11379),
            .I(N__11350));
    LocalMux I__1810 (
            .O(N__11372),
            .I(N__11343));
    LocalMux I__1809 (
            .O(N__11367),
            .I(N__11343));
    LocalMux I__1808 (
            .O(N__11364),
            .I(N__11343));
    Span4Mux_v I__1807 (
            .O(N__11361),
            .I(N__11335));
    InMux I__1806 (
            .O(N__11360),
            .I(N__11332));
    InMux I__1805 (
            .O(N__11359),
            .I(N__11323));
    InMux I__1804 (
            .O(N__11358),
            .I(N__11323));
    InMux I__1803 (
            .O(N__11357),
            .I(N__11323));
    InMux I__1802 (
            .O(N__11356),
            .I(N__11323));
    LocalMux I__1801 (
            .O(N__11353),
            .I(N__11320));
    LocalMux I__1800 (
            .O(N__11350),
            .I(N__11315));
    Span4Mux_v I__1799 (
            .O(N__11343),
            .I(N__11315));
    InMux I__1798 (
            .O(N__11342),
            .I(N__11310));
    InMux I__1797 (
            .O(N__11341),
            .I(N__11310));
    InMux I__1796 (
            .O(N__11340),
            .I(N__11303));
    InMux I__1795 (
            .O(N__11339),
            .I(N__11303));
    InMux I__1794 (
            .O(N__11338),
            .I(N__11303));
    Odrv4 I__1793 (
            .O(N__11335),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    LocalMux I__1792 (
            .O(N__11332),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    LocalMux I__1791 (
            .O(N__11323),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    Odrv4 I__1790 (
            .O(N__11320),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    Odrv4 I__1789 (
            .O(N__11315),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    LocalMux I__1788 (
            .O(N__11310),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    LocalMux I__1787 (
            .O(N__11303),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ));
    InMux I__1786 (
            .O(N__11288),
            .I(N__11285));
    LocalMux I__1785 (
            .O(N__11285),
            .I(\this_vga_signals.vaddress_4_6 ));
    CascadeMux I__1784 (
            .O(N__11282),
            .I(\this_vga_signals.M_vcounter_d7lto8_1_cascade_ ));
    InMux I__1783 (
            .O(N__11279),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__1782 (
            .O(N__11276),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__1781 (
            .O(N__11273),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__1780 (
            .O(N__11270),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__1779 (
            .O(N__11267),
            .I(N__11261));
    InMux I__1778 (
            .O(N__11266),
            .I(N__11261));
    LocalMux I__1777 (
            .O(N__11261),
            .I(N__11257));
    InMux I__1776 (
            .O(N__11260),
            .I(N__11254));
    Span4Mux_h I__1775 (
            .O(N__11257),
            .I(N__11251));
    LocalMux I__1774 (
            .O(N__11254),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    Odrv4 I__1773 (
            .O(N__11251),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    InMux I__1772 (
            .O(N__11246),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    InMux I__1771 (
            .O(N__11243),
            .I(bfn_13_18_0_));
    InMux I__1770 (
            .O(N__11240),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    InMux I__1769 (
            .O(N__11237),
            .I(N__11234));
    LocalMux I__1768 (
            .O(N__11234),
            .I(N__11229));
    InMux I__1767 (
            .O(N__11233),
            .I(N__11226));
    InMux I__1766 (
            .O(N__11232),
            .I(N__11223));
    Odrv12 I__1765 (
            .O(N__11229),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    LocalMux I__1764 (
            .O(N__11226),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    LocalMux I__1763 (
            .O(N__11223),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    InMux I__1762 (
            .O(N__11216),
            .I(N__11213));
    LocalMux I__1761 (
            .O(N__11213),
            .I(\this_vga_signals.vsync_1_3 ));
    IoInMux I__1760 (
            .O(N__11210),
            .I(N__11207));
    LocalMux I__1759 (
            .O(N__11207),
            .I(N__11204));
    Span4Mux_s2_v I__1758 (
            .O(N__11204),
            .I(N__11201));
    Sp12to4 I__1757 (
            .O(N__11201),
            .I(N__11198));
    Span12Mux_s11_h I__1756 (
            .O(N__11198),
            .I(N__11195));
    Odrv12 I__1755 (
            .O(N__11195),
            .I(this_vga_signals_vsync_1_i));
    CascadeMux I__1754 (
            .O(N__11192),
            .I(N__11188));
    InMux I__1753 (
            .O(N__11191),
            .I(N__11183));
    InMux I__1752 (
            .O(N__11188),
            .I(N__11179));
    InMux I__1751 (
            .O(N__11187),
            .I(N__11176));
    CascadeMux I__1750 (
            .O(N__11186),
            .I(N__11170));
    LocalMux I__1749 (
            .O(N__11183),
            .I(N__11166));
    InMux I__1748 (
            .O(N__11182),
            .I(N__11163));
    LocalMux I__1747 (
            .O(N__11179),
            .I(N__11158));
    LocalMux I__1746 (
            .O(N__11176),
            .I(N__11158));
    InMux I__1745 (
            .O(N__11175),
            .I(N__11155));
    InMux I__1744 (
            .O(N__11174),
            .I(N__11152));
    InMux I__1743 (
            .O(N__11173),
            .I(N__11145));
    InMux I__1742 (
            .O(N__11170),
            .I(N__11145));
    InMux I__1741 (
            .O(N__11169),
            .I(N__11145));
    Odrv4 I__1740 (
            .O(N__11166),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1739 (
            .O(N__11163),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv12 I__1738 (
            .O(N__11158),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1737 (
            .O(N__11155),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1736 (
            .O(N__11152),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1735 (
            .O(N__11145),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    CascadeMux I__1734 (
            .O(N__11132),
            .I(N__11124));
    InMux I__1733 (
            .O(N__11131),
            .I(N__11115));
    InMux I__1732 (
            .O(N__11130),
            .I(N__11115));
    InMux I__1731 (
            .O(N__11129),
            .I(N__11112));
    CascadeMux I__1730 (
            .O(N__11128),
            .I(N__11108));
    InMux I__1729 (
            .O(N__11127),
            .I(N__11103));
    InMux I__1728 (
            .O(N__11124),
            .I(N__11100));
    InMux I__1727 (
            .O(N__11123),
            .I(N__11095));
    InMux I__1726 (
            .O(N__11122),
            .I(N__11095));
    InMux I__1725 (
            .O(N__11121),
            .I(N__11092));
    InMux I__1724 (
            .O(N__11120),
            .I(N__11089));
    LocalMux I__1723 (
            .O(N__11115),
            .I(N__11084));
    LocalMux I__1722 (
            .O(N__11112),
            .I(N__11084));
    InMux I__1721 (
            .O(N__11111),
            .I(N__11075));
    InMux I__1720 (
            .O(N__11108),
            .I(N__11075));
    InMux I__1719 (
            .O(N__11107),
            .I(N__11075));
    InMux I__1718 (
            .O(N__11106),
            .I(N__11075));
    LocalMux I__1717 (
            .O(N__11103),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1716 (
            .O(N__11100),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1715 (
            .O(N__11095),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1714 (
            .O(N__11092),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1713 (
            .O(N__11089),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1712 (
            .O(N__11084),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1711 (
            .O(N__11075),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    InMux I__1710 (
            .O(N__11060),
            .I(N__11052));
    CascadeMux I__1709 (
            .O(N__11059),
            .I(N__11049));
    CascadeMux I__1708 (
            .O(N__11058),
            .I(N__11044));
    CascadeMux I__1707 (
            .O(N__11057),
            .I(N__11041));
    InMux I__1706 (
            .O(N__11056),
            .I(N__11038));
    InMux I__1705 (
            .O(N__11055),
            .I(N__11035));
    LocalMux I__1704 (
            .O(N__11052),
            .I(N__11032));
    InMux I__1703 (
            .O(N__11049),
            .I(N__11029));
    InMux I__1702 (
            .O(N__11048),
            .I(N__11023));
    InMux I__1701 (
            .O(N__11047),
            .I(N__11020));
    InMux I__1700 (
            .O(N__11044),
            .I(N__11015));
    InMux I__1699 (
            .O(N__11041),
            .I(N__11015));
    LocalMux I__1698 (
            .O(N__11038),
            .I(N__11006));
    LocalMux I__1697 (
            .O(N__11035),
            .I(N__11006));
    Span4Mux_h I__1696 (
            .O(N__11032),
            .I(N__11006));
    LocalMux I__1695 (
            .O(N__11029),
            .I(N__11006));
    InMux I__1694 (
            .O(N__11028),
            .I(N__10999));
    InMux I__1693 (
            .O(N__11027),
            .I(N__10999));
    InMux I__1692 (
            .O(N__11026),
            .I(N__10999));
    LocalMux I__1691 (
            .O(N__11023),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1690 (
            .O(N__11020),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1689 (
            .O(N__11015),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__1688 (
            .O(N__11006),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1687 (
            .O(N__10999),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    InMux I__1686 (
            .O(N__10988),
            .I(N__10984));
    InMux I__1685 (
            .O(N__10987),
            .I(N__10978));
    LocalMux I__1684 (
            .O(N__10984),
            .I(N__10975));
    CascadeMux I__1683 (
            .O(N__10983),
            .I(N__10968));
    InMux I__1682 (
            .O(N__10982),
            .I(N__10965));
    InMux I__1681 (
            .O(N__10981),
            .I(N__10962));
    LocalMux I__1680 (
            .O(N__10978),
            .I(N__10957));
    Span4Mux_v I__1679 (
            .O(N__10975),
            .I(N__10957));
    InMux I__1678 (
            .O(N__10974),
            .I(N__10954));
    InMux I__1677 (
            .O(N__10973),
            .I(N__10951));
    InMux I__1676 (
            .O(N__10972),
            .I(N__10944));
    InMux I__1675 (
            .O(N__10971),
            .I(N__10944));
    InMux I__1674 (
            .O(N__10968),
            .I(N__10944));
    LocalMux I__1673 (
            .O(N__10965),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1672 (
            .O(N__10962),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__1671 (
            .O(N__10957),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1670 (
            .O(N__10954),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1669 (
            .O(N__10951),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1668 (
            .O(N__10944),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    CascadeMux I__1667 (
            .O(N__10931),
            .I(\this_vga_signals.M_hcounter_d7lto7_0_cascade_ ));
    CascadeMux I__1666 (
            .O(N__10928),
            .I(N__10924));
    InMux I__1665 (
            .O(N__10927),
            .I(N__10920));
    InMux I__1664 (
            .O(N__10924),
            .I(N__10916));
    InMux I__1663 (
            .O(N__10923),
            .I(N__10913));
    LocalMux I__1662 (
            .O(N__10920),
            .I(N__10910));
    InMux I__1661 (
            .O(N__10919),
            .I(N__10902));
    LocalMux I__1660 (
            .O(N__10916),
            .I(N__10895));
    LocalMux I__1659 (
            .O(N__10913),
            .I(N__10895));
    Span4Mux_v I__1658 (
            .O(N__10910),
            .I(N__10895));
    InMux I__1657 (
            .O(N__10909),
            .I(N__10892));
    InMux I__1656 (
            .O(N__10908),
            .I(N__10889));
    InMux I__1655 (
            .O(N__10907),
            .I(N__10882));
    InMux I__1654 (
            .O(N__10906),
            .I(N__10882));
    InMux I__1653 (
            .O(N__10905),
            .I(N__10882));
    LocalMux I__1652 (
            .O(N__10902),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__1651 (
            .O(N__10895),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1650 (
            .O(N__10892),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1649 (
            .O(N__10889),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1648 (
            .O(N__10882),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    InMux I__1647 (
            .O(N__10871),
            .I(N__10868));
    LocalMux I__1646 (
            .O(N__10868),
            .I(\this_vga_signals.un2_vsynclt8 ));
    CEMux I__1645 (
            .O(N__10865),
            .I(N__10862));
    LocalMux I__1644 (
            .O(N__10862),
            .I(\this_vga_signals.N_340_1 ));
    InMux I__1643 (
            .O(N__10859),
            .I(N__10856));
    LocalMux I__1642 (
            .O(N__10856),
            .I(\this_vga_signals.vsync_1_2 ));
    InMux I__1641 (
            .O(N__10853),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    InMux I__1640 (
            .O(N__10850),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__1639 (
            .O(N__10847),
            .I(N__10844));
    LocalMux I__1638 (
            .O(N__10844),
            .I(\this_vga_signals.g2_1 ));
    InMux I__1637 (
            .O(N__10841),
            .I(N__10838));
    LocalMux I__1636 (
            .O(N__10838),
            .I(N__10834));
    InMux I__1635 (
            .O(N__10837),
            .I(N__10831));
    Odrv4 I__1634 (
            .O(N__10834),
            .I(\this_vga_signals.if_N_5 ));
    LocalMux I__1633 (
            .O(N__10831),
            .I(\this_vga_signals.if_N_5 ));
    CascadeMux I__1632 (
            .O(N__10826),
            .I(N__10823));
    InMux I__1631 (
            .O(N__10823),
            .I(N__10820));
    LocalMux I__1630 (
            .O(N__10820),
            .I(\this_vga_signals.vaddress_4_5 ));
    InMux I__1629 (
            .O(N__10817),
            .I(N__10814));
    LocalMux I__1628 (
            .O(N__10814),
            .I(\this_vga_signals.vaddress_3_6 ));
    CascadeMux I__1627 (
            .O(N__10811),
            .I(N__10802));
    InMux I__1626 (
            .O(N__10810),
            .I(N__10796));
    InMux I__1625 (
            .O(N__10809),
            .I(N__10796));
    InMux I__1624 (
            .O(N__10808),
            .I(N__10793));
    InMux I__1623 (
            .O(N__10807),
            .I(N__10784));
    InMux I__1622 (
            .O(N__10806),
            .I(N__10784));
    InMux I__1621 (
            .O(N__10805),
            .I(N__10780));
    InMux I__1620 (
            .O(N__10802),
            .I(N__10774));
    InMux I__1619 (
            .O(N__10801),
            .I(N__10774));
    LocalMux I__1618 (
            .O(N__10796),
            .I(N__10768));
    LocalMux I__1617 (
            .O(N__10793),
            .I(N__10768));
    CascadeMux I__1616 (
            .O(N__10792),
            .I(N__10761));
    CascadeMux I__1615 (
            .O(N__10791),
            .I(N__10757));
    CascadeMux I__1614 (
            .O(N__10790),
            .I(N__10752));
    CascadeMux I__1613 (
            .O(N__10789),
            .I(N__10749));
    LocalMux I__1612 (
            .O(N__10784),
            .I(N__10746));
    InMux I__1611 (
            .O(N__10783),
            .I(N__10743));
    LocalMux I__1610 (
            .O(N__10780),
            .I(N__10740));
    InMux I__1609 (
            .O(N__10779),
            .I(N__10737));
    LocalMux I__1608 (
            .O(N__10774),
            .I(N__10734));
    InMux I__1607 (
            .O(N__10773),
            .I(N__10731));
    Span4Mux_v I__1606 (
            .O(N__10768),
            .I(N__10728));
    InMux I__1605 (
            .O(N__10767),
            .I(N__10715));
    InMux I__1604 (
            .O(N__10766),
            .I(N__10715));
    InMux I__1603 (
            .O(N__10765),
            .I(N__10715));
    InMux I__1602 (
            .O(N__10764),
            .I(N__10715));
    InMux I__1601 (
            .O(N__10761),
            .I(N__10715));
    InMux I__1600 (
            .O(N__10760),
            .I(N__10715));
    InMux I__1599 (
            .O(N__10757),
            .I(N__10704));
    InMux I__1598 (
            .O(N__10756),
            .I(N__10704));
    InMux I__1597 (
            .O(N__10755),
            .I(N__10704));
    InMux I__1596 (
            .O(N__10752),
            .I(N__10704));
    InMux I__1595 (
            .O(N__10749),
            .I(N__10704));
    Odrv4 I__1594 (
            .O(N__10746),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1593 (
            .O(N__10743),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__1592 (
            .O(N__10740),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1591 (
            .O(N__10737),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__1590 (
            .O(N__10734),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1589 (
            .O(N__10731),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__1588 (
            .O(N__10728),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1587 (
            .O(N__10715),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1586 (
            .O(N__10704),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    CascadeMux I__1585 (
            .O(N__10685),
            .I(\this_vga_signals.vaddress_0_5_cascade_ ));
    InMux I__1584 (
            .O(N__10682),
            .I(N__10677));
    InMux I__1583 (
            .O(N__10681),
            .I(N__10674));
    InMux I__1582 (
            .O(N__10680),
            .I(N__10666));
    LocalMux I__1581 (
            .O(N__10677),
            .I(N__10663));
    LocalMux I__1580 (
            .O(N__10674),
            .I(N__10660));
    InMux I__1579 (
            .O(N__10673),
            .I(N__10655));
    InMux I__1578 (
            .O(N__10672),
            .I(N__10655));
    InMux I__1577 (
            .O(N__10671),
            .I(N__10652));
    InMux I__1576 (
            .O(N__10670),
            .I(N__10649));
    InMux I__1575 (
            .O(N__10669),
            .I(N__10635));
    LocalMux I__1574 (
            .O(N__10666),
            .I(N__10630));
    Span4Mux_v I__1573 (
            .O(N__10663),
            .I(N__10630));
    Span4Mux_h I__1572 (
            .O(N__10660),
            .I(N__10627));
    LocalMux I__1571 (
            .O(N__10655),
            .I(N__10624));
    LocalMux I__1570 (
            .O(N__10652),
            .I(N__10621));
    LocalMux I__1569 (
            .O(N__10649),
            .I(N__10618));
    InMux I__1568 (
            .O(N__10648),
            .I(N__10607));
    InMux I__1567 (
            .O(N__10647),
            .I(N__10607));
    InMux I__1566 (
            .O(N__10646),
            .I(N__10607));
    InMux I__1565 (
            .O(N__10645),
            .I(N__10607));
    InMux I__1564 (
            .O(N__10644),
            .I(N__10607));
    InMux I__1563 (
            .O(N__10643),
            .I(N__10594));
    InMux I__1562 (
            .O(N__10642),
            .I(N__10594));
    InMux I__1561 (
            .O(N__10641),
            .I(N__10594));
    InMux I__1560 (
            .O(N__10640),
            .I(N__10594));
    InMux I__1559 (
            .O(N__10639),
            .I(N__10594));
    InMux I__1558 (
            .O(N__10638),
            .I(N__10594));
    LocalMux I__1557 (
            .O(N__10635),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__1556 (
            .O(N__10630),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__1555 (
            .O(N__10627),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__1554 (
            .O(N__10624),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__1553 (
            .O(N__10621),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv12 I__1552 (
            .O(N__10618),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__1551 (
            .O(N__10607),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__1550 (
            .O(N__10594),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    CascadeMux I__1549 (
            .O(N__10577),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0_cascade_ ));
    InMux I__1548 (
            .O(N__10574),
            .I(N__10571));
    LocalMux I__1547 (
            .O(N__10571),
            .I(\this_vga_signals.g2 ));
    InMux I__1546 (
            .O(N__10568),
            .I(N__10565));
    LocalMux I__1545 (
            .O(N__10565),
            .I(\this_vga_signals.g1 ));
    InMux I__1544 (
            .O(N__10562),
            .I(N__10558));
    InMux I__1543 (
            .O(N__10561),
            .I(N__10555));
    LocalMux I__1542 (
            .O(N__10558),
            .I(\this_vga_signals.vaddress_0_6 ));
    LocalMux I__1541 (
            .O(N__10555),
            .I(\this_vga_signals.vaddress_0_6 ));
    InMux I__1540 (
            .O(N__10550),
            .I(N__10547));
    LocalMux I__1539 (
            .O(N__10547),
            .I(\this_vga_signals.g1_0_2 ));
    InMux I__1538 (
            .O(N__10544),
            .I(N__10541));
    LocalMux I__1537 (
            .O(N__10541),
            .I(\this_vga_signals.g0_31_1 ));
    CascadeMux I__1536 (
            .O(N__10538),
            .I(N__10535));
    InMux I__1535 (
            .O(N__10535),
            .I(N__10532));
    LocalMux I__1534 (
            .O(N__10532),
            .I(\this_vga_signals.g1_0_1 ));
    InMux I__1533 (
            .O(N__10529),
            .I(N__10525));
    InMux I__1532 (
            .O(N__10528),
            .I(N__10519));
    LocalMux I__1531 (
            .O(N__10525),
            .I(N__10516));
    InMux I__1530 (
            .O(N__10524),
            .I(N__10513));
    InMux I__1529 (
            .O(N__10523),
            .I(N__10508));
    InMux I__1528 (
            .O(N__10522),
            .I(N__10508));
    LocalMux I__1527 (
            .O(N__10519),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_N_2L1 ));
    Odrv4 I__1526 (
            .O(N__10516),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_N_2L1 ));
    LocalMux I__1525 (
            .O(N__10513),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_N_2L1 ));
    LocalMux I__1524 (
            .O(N__10508),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_N_2L1 ));
    InMux I__1523 (
            .O(N__10499),
            .I(N__10496));
    LocalMux I__1522 (
            .O(N__10496),
            .I(\this_vga_signals.N_5_1_0_0 ));
    InMux I__1521 (
            .O(N__10493),
            .I(N__10490));
    LocalMux I__1520 (
            .O(N__10490),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2_0_1_0 ));
    CascadeMux I__1519 (
            .O(N__10487),
            .I(\this_vga_signals.g0_22_1_cascade_ ));
    InMux I__1518 (
            .O(N__10484),
            .I(N__10481));
    LocalMux I__1517 (
            .O(N__10481),
            .I(N__10478));
    Odrv12 I__1516 (
            .O(N__10478),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0_0_0_0 ));
    InMux I__1515 (
            .O(N__10475),
            .I(N__10471));
    InMux I__1514 (
            .O(N__10474),
            .I(N__10468));
    LocalMux I__1513 (
            .O(N__10471),
            .I(\this_vga_signals.mult1_un61_sum_c3_0 ));
    LocalMux I__1512 (
            .O(N__10468),
            .I(\this_vga_signals.mult1_un61_sum_c3_0 ));
    CascadeMux I__1511 (
            .O(N__10463),
            .I(\this_vga_signals.vaddress_5_5_cascade_ ));
    InMux I__1510 (
            .O(N__10460),
            .I(N__10457));
    LocalMux I__1509 (
            .O(N__10457),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_1 ));
    CascadeMux I__1508 (
            .O(N__10454),
            .I(N__10446));
    CascadeMux I__1507 (
            .O(N__10453),
            .I(N__10443));
    InMux I__1506 (
            .O(N__10452),
            .I(N__10440));
    InMux I__1505 (
            .O(N__10451),
            .I(N__10435));
    InMux I__1504 (
            .O(N__10450),
            .I(N__10435));
    InMux I__1503 (
            .O(N__10449),
            .I(N__10430));
    InMux I__1502 (
            .O(N__10446),
            .I(N__10430));
    InMux I__1501 (
            .O(N__10443),
            .I(N__10427));
    LocalMux I__1500 (
            .O(N__10440),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__1499 (
            .O(N__10435),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__1498 (
            .O(N__10430),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__1497 (
            .O(N__10427),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    CascadeMux I__1496 (
            .O(N__10418),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_1_cascade_ ));
    InMux I__1495 (
            .O(N__10415),
            .I(N__10409));
    InMux I__1494 (
            .O(N__10414),
            .I(N__10409));
    LocalMux I__1493 (
            .O(N__10409),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0_0 ));
    InMux I__1492 (
            .O(N__10406),
            .I(N__10403));
    LocalMux I__1491 (
            .O(N__10403),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_0_0_0 ));
    InMux I__1490 (
            .O(N__10400),
            .I(N__10397));
    LocalMux I__1489 (
            .O(N__10397),
            .I(N__10394));
    Span4Mux_h I__1488 (
            .O(N__10394),
            .I(N__10383));
    InMux I__1487 (
            .O(N__10393),
            .I(N__10380));
    InMux I__1486 (
            .O(N__10392),
            .I(N__10375));
    InMux I__1485 (
            .O(N__10391),
            .I(N__10375));
    InMux I__1484 (
            .O(N__10390),
            .I(N__10372));
    InMux I__1483 (
            .O(N__10389),
            .I(N__10367));
    InMux I__1482 (
            .O(N__10388),
            .I(N__10367));
    InMux I__1481 (
            .O(N__10387),
            .I(N__10362));
    InMux I__1480 (
            .O(N__10386),
            .I(N__10362));
    Odrv4 I__1479 (
            .O(N__10383),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1478 (
            .O(N__10380),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1477 (
            .O(N__10375),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1476 (
            .O(N__10372),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1475 (
            .O(N__10367),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1474 (
            .O(N__10362),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    InMux I__1473 (
            .O(N__10349),
            .I(N__10346));
    LocalMux I__1472 (
            .O(N__10346),
            .I(N__10343));
    Span4Mux_h I__1471 (
            .O(N__10343),
            .I(N__10339));
    InMux I__1470 (
            .O(N__10342),
            .I(N__10336));
    Odrv4 I__1469 (
            .O(N__10339),
            .I(\this_vga_signals.vaddress_2_0_6 ));
    LocalMux I__1468 (
            .O(N__10336),
            .I(\this_vga_signals.vaddress_2_0_6 ));
    CascadeMux I__1467 (
            .O(N__10331),
            .I(N__10328));
    InMux I__1466 (
            .O(N__10328),
            .I(N__10325));
    LocalMux I__1465 (
            .O(N__10325),
            .I(\this_vga_signals.g0_7_0 ));
    CascadeMux I__1464 (
            .O(N__10322),
            .I(N__10315));
    CascadeMux I__1463 (
            .O(N__10321),
            .I(N__10312));
    InMux I__1462 (
            .O(N__10320),
            .I(N__10309));
    InMux I__1461 (
            .O(N__10319),
            .I(N__10306));
    InMux I__1460 (
            .O(N__10318),
            .I(N__10303));
    InMux I__1459 (
            .O(N__10315),
            .I(N__10300));
    InMux I__1458 (
            .O(N__10312),
            .I(N__10297));
    LocalMux I__1457 (
            .O(N__10309),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__1456 (
            .O(N__10306),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__1455 (
            .O(N__10303),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__1454 (
            .O(N__10300),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__1453 (
            .O(N__10297),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    InMux I__1452 (
            .O(N__10286),
            .I(N__10283));
    LocalMux I__1451 (
            .O(N__10283),
            .I(N__10280));
    Odrv4 I__1450 (
            .O(N__10280),
            .I(\this_vga_signals.mult1_un40_sum_axb1_0 ));
    CascadeMux I__1449 (
            .O(N__10277),
            .I(N__10274));
    InMux I__1448 (
            .O(N__10274),
            .I(N__10264));
    InMux I__1447 (
            .O(N__10273),
            .I(N__10264));
    InMux I__1446 (
            .O(N__10272),
            .I(N__10259));
    InMux I__1445 (
            .O(N__10271),
            .I(N__10259));
    InMux I__1444 (
            .O(N__10270),
            .I(N__10256));
    InMux I__1443 (
            .O(N__10269),
            .I(N__10253));
    LocalMux I__1442 (
            .O(N__10264),
            .I(N__10248));
    LocalMux I__1441 (
            .O(N__10259),
            .I(N__10248));
    LocalMux I__1440 (
            .O(N__10256),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__1439 (
            .O(N__10253),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    Odrv4 I__1438 (
            .O(N__10248),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    CascadeMux I__1437 (
            .O(N__10241),
            .I(\this_vga_signals.if_m8_0_a3_1_1_1_cascade_ ));
    CascadeMux I__1436 (
            .O(N__10238),
            .I(N__10235));
    InMux I__1435 (
            .O(N__10235),
            .I(N__10227));
    InMux I__1434 (
            .O(N__10234),
            .I(N__10224));
    InMux I__1433 (
            .O(N__10233),
            .I(N__10221));
    InMux I__1432 (
            .O(N__10232),
            .I(N__10214));
    InMux I__1431 (
            .O(N__10231),
            .I(N__10214));
    InMux I__1430 (
            .O(N__10230),
            .I(N__10214));
    LocalMux I__1429 (
            .O(N__10227),
            .I(N__10209));
    LocalMux I__1428 (
            .O(N__10224),
            .I(N__10209));
    LocalMux I__1427 (
            .O(N__10221),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__1426 (
            .O(N__10214),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    Odrv4 I__1425 (
            .O(N__10209),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    CascadeMux I__1424 (
            .O(N__10202),
            .I(N__10199));
    InMux I__1423 (
            .O(N__10199),
            .I(N__10196));
    LocalMux I__1422 (
            .O(N__10196),
            .I(N__10193));
    Span4Mux_h I__1421 (
            .O(N__10193),
            .I(N__10190));
    Odrv4 I__1420 (
            .O(N__10190),
            .I(\this_vga_signals.vaddress_2_6 ));
    InMux I__1419 (
            .O(N__10187),
            .I(N__10184));
    LocalMux I__1418 (
            .O(N__10184),
            .I(N__10181));
    Span4Mux_h I__1417 (
            .O(N__10181),
            .I(N__10178));
    Odrv4 I__1416 (
            .O(N__10178),
            .I(\this_vga_signals.vaddress_2_5 ));
    InMux I__1415 (
            .O(N__10175),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__1414 (
            .O(N__10172),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__1413 (
            .O(N__10169),
            .I(bfn_11_23_0_));
    CascadeMux I__1412 (
            .O(N__10166),
            .I(\this_vga_signals.un4_hsynclt8_0_cascade_ ));
    IoInMux I__1411 (
            .O(N__10163),
            .I(N__10160));
    LocalMux I__1410 (
            .O(N__10160),
            .I(N__10157));
    IoSpan4Mux I__1409 (
            .O(N__10157),
            .I(N__10154));
    Span4Mux_s1_v I__1408 (
            .O(N__10154),
            .I(N__10151));
    Sp12to4 I__1407 (
            .O(N__10151),
            .I(N__10148));
    Span12Mux_s8_v I__1406 (
            .O(N__10148),
            .I(N__10145));
    Odrv12 I__1405 (
            .O(N__10145),
            .I(this_vga_signals_hsync_1_i));
    InMux I__1404 (
            .O(N__10142),
            .I(N__10135));
    InMux I__1403 (
            .O(N__10141),
            .I(N__10135));
    CascadeMux I__1402 (
            .O(N__10140),
            .I(N__10130));
    LocalMux I__1401 (
            .O(N__10135),
            .I(N__10124));
    InMux I__1400 (
            .O(N__10134),
            .I(N__10117));
    InMux I__1399 (
            .O(N__10133),
            .I(N__10117));
    InMux I__1398 (
            .O(N__10130),
            .I(N__10114));
    CascadeMux I__1397 (
            .O(N__10129),
            .I(N__10110));
    InMux I__1396 (
            .O(N__10128),
            .I(N__10104));
    InMux I__1395 (
            .O(N__10127),
            .I(N__10104));
    Span4Mux_v I__1394 (
            .O(N__10124),
            .I(N__10101));
    InMux I__1393 (
            .O(N__10123),
            .I(N__10098));
    InMux I__1392 (
            .O(N__10122),
            .I(N__10095));
    LocalMux I__1391 (
            .O(N__10117),
            .I(N__10090));
    LocalMux I__1390 (
            .O(N__10114),
            .I(N__10090));
    InMux I__1389 (
            .O(N__10113),
            .I(N__10083));
    InMux I__1388 (
            .O(N__10110),
            .I(N__10083));
    InMux I__1387 (
            .O(N__10109),
            .I(N__10083));
    LocalMux I__1386 (
            .O(N__10104),
            .I(N__10076));
    Span4Mux_h I__1385 (
            .O(N__10101),
            .I(N__10076));
    LocalMux I__1384 (
            .O(N__10098),
            .I(N__10076));
    LocalMux I__1383 (
            .O(N__10095),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1382 (
            .O(N__10090),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1381 (
            .O(N__10083),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1380 (
            .O(N__10076),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__1379 (
            .O(N__10067),
            .I(N__10064));
    LocalMux I__1378 (
            .O(N__10064),
            .I(\this_vga_signals.un3_hsynclt8_0 ));
    CascadeMux I__1377 (
            .O(N__10061),
            .I(\this_vga_signals.un6_vvisibilitylto8_0_cascade_ ));
    CascadeMux I__1376 (
            .O(N__10058),
            .I(\this_vga_signals.un6_vvisibilitylt9_0_cascade_ ));
    InMux I__1375 (
            .O(N__10055),
            .I(N__10052));
    LocalMux I__1374 (
            .O(N__10052),
            .I(N__10049));
    Span4Mux_h I__1373 (
            .O(N__10049),
            .I(N__10044));
    InMux I__1372 (
            .O(N__10048),
            .I(N__10041));
    CascadeMux I__1371 (
            .O(N__10047),
            .I(N__10038));
    Span4Mux_v I__1370 (
            .O(N__10044),
            .I(N__10035));
    LocalMux I__1369 (
            .O(N__10041),
            .I(N__10032));
    InMux I__1368 (
            .O(N__10038),
            .I(N__10029));
    Span4Mux_h I__1367 (
            .O(N__10035),
            .I(N__10026));
    Span12Mux_s11_h I__1366 (
            .O(N__10032),
            .I(N__10023));
    LocalMux I__1365 (
            .O(N__10029),
            .I(N__10020));
    Odrv4 I__1364 (
            .O(N__10026),
            .I(\this_vga_signals.vvisibility ));
    Odrv12 I__1363 (
            .O(N__10023),
            .I(\this_vga_signals.vvisibility ));
    Odrv4 I__1362 (
            .O(N__10020),
            .I(\this_vga_signals.vvisibility ));
    CascadeMux I__1361 (
            .O(N__10013),
            .I(N__10002));
    InMux I__1360 (
            .O(N__10012),
            .I(N__9994));
    InMux I__1359 (
            .O(N__10011),
            .I(N__9991));
    InMux I__1358 (
            .O(N__10010),
            .I(N__9988));
    InMux I__1357 (
            .O(N__10009),
            .I(N__9983));
    InMux I__1356 (
            .O(N__10008),
            .I(N__9983));
    InMux I__1355 (
            .O(N__10007),
            .I(N__9978));
    InMux I__1354 (
            .O(N__10006),
            .I(N__9978));
    InMux I__1353 (
            .O(N__10005),
            .I(N__9973));
    InMux I__1352 (
            .O(N__10002),
            .I(N__9973));
    InMux I__1351 (
            .O(N__10001),
            .I(N__9962));
    InMux I__1350 (
            .O(N__10000),
            .I(N__9962));
    InMux I__1349 (
            .O(N__9999),
            .I(N__9962));
    InMux I__1348 (
            .O(N__9998),
            .I(N__9962));
    InMux I__1347 (
            .O(N__9997),
            .I(N__9962));
    LocalMux I__1346 (
            .O(N__9994),
            .I(\this_vga_signals.mult1_un68_sum_axb1_395 ));
    LocalMux I__1345 (
            .O(N__9991),
            .I(\this_vga_signals.mult1_un68_sum_axb1_395 ));
    LocalMux I__1344 (
            .O(N__9988),
            .I(\this_vga_signals.mult1_un68_sum_axb1_395 ));
    LocalMux I__1343 (
            .O(N__9983),
            .I(\this_vga_signals.mult1_un68_sum_axb1_395 ));
    LocalMux I__1342 (
            .O(N__9978),
            .I(\this_vga_signals.mult1_un68_sum_axb1_395 ));
    LocalMux I__1341 (
            .O(N__9973),
            .I(\this_vga_signals.mult1_un68_sum_axb1_395 ));
    LocalMux I__1340 (
            .O(N__9962),
            .I(\this_vga_signals.mult1_un68_sum_axb1_395 ));
    InMux I__1339 (
            .O(N__9947),
            .I(N__9944));
    LocalMux I__1338 (
            .O(N__9944),
            .I(\this_vga_signals.mult1_un68_sum_ac0_1_x0 ));
    InMux I__1337 (
            .O(N__9941),
            .I(N__9938));
    LocalMux I__1336 (
            .O(N__9938),
            .I(N__9933));
    InMux I__1335 (
            .O(N__9937),
            .I(N__9928));
    InMux I__1334 (
            .O(N__9936),
            .I(N__9928));
    Odrv4 I__1333 (
            .O(N__9933),
            .I(\this_vga_signals.mult1_un61_sum_c3_1 ));
    LocalMux I__1332 (
            .O(N__9928),
            .I(\this_vga_signals.mult1_un61_sum_c3_1 ));
    InMux I__1331 (
            .O(N__9923),
            .I(N__9920));
    LocalMux I__1330 (
            .O(N__9920),
            .I(\this_vga_signals.g0_2_x1 ));
    CascadeMux I__1329 (
            .O(N__9917),
            .I(N__9903));
    CascadeMux I__1328 (
            .O(N__9916),
            .I(N__9899));
    CascadeMux I__1327 (
            .O(N__9915),
            .I(N__9896));
    CascadeMux I__1326 (
            .O(N__9914),
            .I(N__9891));
    CascadeMux I__1325 (
            .O(N__9913),
            .I(N__9888));
    InMux I__1324 (
            .O(N__9912),
            .I(N__9883));
    InMux I__1323 (
            .O(N__9911),
            .I(N__9880));
    InMux I__1322 (
            .O(N__9910),
            .I(N__9869));
    InMux I__1321 (
            .O(N__9909),
            .I(N__9869));
    InMux I__1320 (
            .O(N__9908),
            .I(N__9869));
    InMux I__1319 (
            .O(N__9907),
            .I(N__9869));
    InMux I__1318 (
            .O(N__9906),
            .I(N__9869));
    InMux I__1317 (
            .O(N__9903),
            .I(N__9864));
    InMux I__1316 (
            .O(N__9902),
            .I(N__9864));
    InMux I__1315 (
            .O(N__9899),
            .I(N__9855));
    InMux I__1314 (
            .O(N__9896),
            .I(N__9855));
    InMux I__1313 (
            .O(N__9895),
            .I(N__9855));
    InMux I__1312 (
            .O(N__9894),
            .I(N__9855));
    InMux I__1311 (
            .O(N__9891),
            .I(N__9846));
    InMux I__1310 (
            .O(N__9888),
            .I(N__9846));
    InMux I__1309 (
            .O(N__9887),
            .I(N__9846));
    InMux I__1308 (
            .O(N__9886),
            .I(N__9846));
    LocalMux I__1307 (
            .O(N__9883),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    LocalMux I__1306 (
            .O(N__9880),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    LocalMux I__1305 (
            .O(N__9869),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    LocalMux I__1304 (
            .O(N__9864),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    LocalMux I__1303 (
            .O(N__9855),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    LocalMux I__1302 (
            .O(N__9846),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    InMux I__1301 (
            .O(N__9833),
            .I(N__9830));
    LocalMux I__1300 (
            .O(N__9830),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1 ));
    InMux I__1299 (
            .O(N__9827),
            .I(N__9823));
    CascadeMux I__1298 (
            .O(N__9826),
            .I(N__9815));
    LocalMux I__1297 (
            .O(N__9823),
            .I(N__9812));
    InMux I__1296 (
            .O(N__9822),
            .I(N__9805));
    InMux I__1295 (
            .O(N__9821),
            .I(N__9805));
    InMux I__1294 (
            .O(N__9820),
            .I(N__9805));
    InMux I__1293 (
            .O(N__9819),
            .I(N__9800));
    InMux I__1292 (
            .O(N__9818),
            .I(N__9800));
    InMux I__1291 (
            .O(N__9815),
            .I(N__9797));
    Span4Mux_v I__1290 (
            .O(N__9812),
            .I(N__9791));
    LocalMux I__1289 (
            .O(N__9805),
            .I(N__9791));
    LocalMux I__1288 (
            .O(N__9800),
            .I(N__9786));
    LocalMux I__1287 (
            .O(N__9797),
            .I(N__9786));
    InMux I__1286 (
            .O(N__9796),
            .I(N__9783));
    Span4Mux_h I__1285 (
            .O(N__9791),
            .I(N__9780));
    Span12Mux_s10_h I__1284 (
            .O(N__9786),
            .I(N__9777));
    LocalMux I__1283 (
            .O(N__9783),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1282 (
            .O(N__9780),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv12 I__1281 (
            .O(N__9777),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__1280 (
            .O(N__9770),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    CascadeMux I__1279 (
            .O(N__9767),
            .I(N__9764));
    InMux I__1278 (
            .O(N__9764),
            .I(N__9756));
    InMux I__1277 (
            .O(N__9763),
            .I(N__9756));
    InMux I__1276 (
            .O(N__9762),
            .I(N__9753));
    CascadeMux I__1275 (
            .O(N__9761),
            .I(N__9747));
    LocalMux I__1274 (
            .O(N__9756),
            .I(N__9742));
    LocalMux I__1273 (
            .O(N__9753),
            .I(N__9739));
    CascadeMux I__1272 (
            .O(N__9752),
            .I(N__9736));
    CascadeMux I__1271 (
            .O(N__9751),
            .I(N__9732));
    InMux I__1270 (
            .O(N__9750),
            .I(N__9727));
    InMux I__1269 (
            .O(N__9747),
            .I(N__9727));
    InMux I__1268 (
            .O(N__9746),
            .I(N__9722));
    InMux I__1267 (
            .O(N__9745),
            .I(N__9722));
    Span4Mux_v I__1266 (
            .O(N__9742),
            .I(N__9716));
    Span4Mux_h I__1265 (
            .O(N__9739),
            .I(N__9716));
    InMux I__1264 (
            .O(N__9736),
            .I(N__9709));
    InMux I__1263 (
            .O(N__9735),
            .I(N__9709));
    InMux I__1262 (
            .O(N__9732),
            .I(N__9709));
    LocalMux I__1261 (
            .O(N__9727),
            .I(N__9704));
    LocalMux I__1260 (
            .O(N__9722),
            .I(N__9704));
    InMux I__1259 (
            .O(N__9721),
            .I(N__9700));
    Span4Mux_h I__1258 (
            .O(N__9716),
            .I(N__9697));
    LocalMux I__1257 (
            .O(N__9709),
            .I(N__9692));
    Span4Mux_v I__1256 (
            .O(N__9704),
            .I(N__9692));
    InMux I__1255 (
            .O(N__9703),
            .I(N__9689));
    LocalMux I__1254 (
            .O(N__9700),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1253 (
            .O(N__9697),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1252 (
            .O(N__9692),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1251 (
            .O(N__9689),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__1250 (
            .O(N__9680),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__1249 (
            .O(N__9677),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__1248 (
            .O(N__9674),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__1247 (
            .O(N__9671),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__1246 (
            .O(N__9668),
            .I(N__9665));
    LocalMux I__1245 (
            .O(N__9665),
            .I(N__9662));
    Odrv4 I__1244 (
            .O(N__9662),
            .I(\this_vga_signals.mult1_un54_sum_axb1_1_0_0 ));
    CascadeMux I__1243 (
            .O(N__9659),
            .I(\this_vga_signals.N_5_i_5_cascade_ ));
    InMux I__1242 (
            .O(N__9656),
            .I(N__9653));
    LocalMux I__1241 (
            .O(N__9653),
            .I(\this_vga_signals.N_20_0 ));
    InMux I__1240 (
            .O(N__9650),
            .I(N__9647));
    LocalMux I__1239 (
            .O(N__9647),
            .I(\this_vga_signals.g1_1_1 ));
    InMux I__1238 (
            .O(N__9644),
            .I(N__9641));
    LocalMux I__1237 (
            .O(N__9641),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_0_0 ));
    CascadeMux I__1236 (
            .O(N__9638),
            .I(\this_vga_signals.g0_2_x0_cascade_ ));
    CascadeMux I__1235 (
            .O(N__9635),
            .I(\this_vga_signals.g1_0_0_0_cascade_ ));
    InMux I__1234 (
            .O(N__9632),
            .I(N__9629));
    LocalMux I__1233 (
            .O(N__9629),
            .I(\this_vga_signals.N_5_i_5 ));
    CascadeMux I__1232 (
            .O(N__9626),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_ ));
    InMux I__1231 (
            .O(N__9623),
            .I(N__9620));
    LocalMux I__1230 (
            .O(N__9620),
            .I(\this_vga_signals.g0_i_x2_0_2_0 ));
    InMux I__1229 (
            .O(N__9617),
            .I(N__9614));
    LocalMux I__1228 (
            .O(N__9614),
            .I(N__9611));
    Span4Mux_h I__1227 (
            .O(N__9611),
            .I(N__9608));
    Odrv4 I__1226 (
            .O(N__9608),
            .I(\this_vga_signals.if_i4_mux_0_0_0 ));
    CascadeMux I__1225 (
            .O(N__9605),
            .I(\this_vga_signals.vaddress_6_cascade_ ));
    InMux I__1224 (
            .O(N__9602),
            .I(N__9597));
    CascadeMux I__1223 (
            .O(N__9601),
            .I(N__9593));
    InMux I__1222 (
            .O(N__9600),
            .I(N__9589));
    LocalMux I__1221 (
            .O(N__9597),
            .I(N__9586));
    InMux I__1220 (
            .O(N__9596),
            .I(N__9583));
    InMux I__1219 (
            .O(N__9593),
            .I(N__9578));
    InMux I__1218 (
            .O(N__9592),
            .I(N__9578));
    LocalMux I__1217 (
            .O(N__9589),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    Odrv4 I__1216 (
            .O(N__9586),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__1215 (
            .O(N__9583),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__1214 (
            .O(N__9578),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    InMux I__1213 (
            .O(N__9569),
            .I(N__9566));
    LocalMux I__1212 (
            .O(N__9566),
            .I(N__9563));
    Odrv4 I__1211 (
            .O(N__9563),
            .I(\this_vga_signals.g1_3_0 ));
    CascadeMux I__1210 (
            .O(N__9560),
            .I(N__9554));
    InMux I__1209 (
            .O(N__9559),
            .I(N__9551));
    InMux I__1208 (
            .O(N__9558),
            .I(N__9544));
    InMux I__1207 (
            .O(N__9557),
            .I(N__9544));
    InMux I__1206 (
            .O(N__9554),
            .I(N__9544));
    LocalMux I__1205 (
            .O(N__9551),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__1204 (
            .O(N__9544),
            .I(\this_vga_signals.vaddress_6 ));
    InMux I__1203 (
            .O(N__9539),
            .I(N__9536));
    LocalMux I__1202 (
            .O(N__9536),
            .I(N__9533));
    Odrv4 I__1201 (
            .O(N__9533),
            .I(\this_vga_signals.vaddress_4_0_6 ));
    CascadeMux I__1200 (
            .O(N__9530),
            .I(N__9527));
    InMux I__1199 (
            .O(N__9527),
            .I(N__9524));
    LocalMux I__1198 (
            .O(N__9524),
            .I(\this_vga_signals.vaddress_5_0_5 ));
    CascadeMux I__1197 (
            .O(N__9521),
            .I(\this_vga_signals.g2_0_cascade_ ));
    InMux I__1196 (
            .O(N__9518),
            .I(N__9515));
    LocalMux I__1195 (
            .O(N__9515),
            .I(\this_vga_signals.mult1_un54_sum_axb1_1 ));
    InMux I__1194 (
            .O(N__9512),
            .I(N__9509));
    LocalMux I__1193 (
            .O(N__9509),
            .I(\this_vga_signals.g1_0_0 ));
    InMux I__1192 (
            .O(N__9506),
            .I(N__9500));
    InMux I__1191 (
            .O(N__9505),
            .I(N__9497));
    InMux I__1190 (
            .O(N__9504),
            .I(N__9492));
    InMux I__1189 (
            .O(N__9503),
            .I(N__9492));
    LocalMux I__1188 (
            .O(N__9500),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__1187 (
            .O(N__9497),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__1186 (
            .O(N__9492),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    CascadeMux I__1185 (
            .O(N__9485),
            .I(N__9482));
    InMux I__1184 (
            .O(N__9482),
            .I(N__9477));
    InMux I__1183 (
            .O(N__9481),
            .I(N__9474));
    InMux I__1182 (
            .O(N__9480),
            .I(N__9471));
    LocalMux I__1181 (
            .O(N__9477),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__1180 (
            .O(N__9474),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__1179 (
            .O(N__9471),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    InMux I__1178 (
            .O(N__9464),
            .I(N__9461));
    LocalMux I__1177 (
            .O(N__9461),
            .I(N__9458));
    Odrv4 I__1176 (
            .O(N__9458),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    CascadeMux I__1175 (
            .O(N__9455),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ));
    InMux I__1174 (
            .O(N__9452),
            .I(N__9449));
    LocalMux I__1173 (
            .O(N__9449),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_0 ));
    CascadeMux I__1172 (
            .O(N__9446),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ));
    IoInMux I__1171 (
            .O(N__9443),
            .I(N__9440));
    LocalMux I__1170 (
            .O(N__9440),
            .I(N__9437));
    IoSpan4Mux I__1169 (
            .O(N__9437),
            .I(N__9434));
    Span4Mux_s2_v I__1168 (
            .O(N__9434),
            .I(N__9431));
    Span4Mux_h I__1167 (
            .O(N__9431),
            .I(N__9428));
    Span4Mux_v I__1166 (
            .O(N__9428),
            .I(N__9425));
    Odrv4 I__1165 (
            .O(N__9425),
            .I(this_vga_signals_hvisibility_i));
    InMux I__1164 (
            .O(N__9422),
            .I(N__9418));
    InMux I__1163 (
            .O(N__9421),
            .I(N__9415));
    LocalMux I__1162 (
            .O(N__9418),
            .I(\this_vga_signals.SUM_3_i_0_0_3 ));
    LocalMux I__1161 (
            .O(N__9415),
            .I(\this_vga_signals.SUM_3_i_0_0_3 ));
    InMux I__1160 (
            .O(N__9410),
            .I(N__9407));
    LocalMux I__1159 (
            .O(N__9407),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ));
    InMux I__1158 (
            .O(N__9404),
            .I(N__9396));
    InMux I__1157 (
            .O(N__9403),
            .I(N__9391));
    InMux I__1156 (
            .O(N__9402),
            .I(N__9391));
    InMux I__1155 (
            .O(N__9401),
            .I(N__9388));
    InMux I__1154 (
            .O(N__9400),
            .I(N__9385));
    CascadeMux I__1153 (
            .O(N__9399),
            .I(N__9382));
    LocalMux I__1152 (
            .O(N__9396),
            .I(N__9376));
    LocalMux I__1151 (
            .O(N__9391),
            .I(N__9376));
    LocalMux I__1150 (
            .O(N__9388),
            .I(N__9371));
    LocalMux I__1149 (
            .O(N__9385),
            .I(N__9371));
    InMux I__1148 (
            .O(N__9382),
            .I(N__9368));
    InMux I__1147 (
            .O(N__9381),
            .I(N__9365));
    Span4Mux_h I__1146 (
            .O(N__9376),
            .I(N__9362));
    Span4Mux_v I__1145 (
            .O(N__9371),
            .I(N__9355));
    LocalMux I__1144 (
            .O(N__9368),
            .I(N__9355));
    LocalMux I__1143 (
            .O(N__9365),
            .I(N__9355));
    Span4Mux_v I__1142 (
            .O(N__9362),
            .I(N__9348));
    Span4Mux_h I__1141 (
            .O(N__9355),
            .I(N__9348));
    InMux I__1140 (
            .O(N__9354),
            .I(N__9345));
    InMux I__1139 (
            .O(N__9353),
            .I(N__9342));
    Odrv4 I__1138 (
            .O(N__9348),
            .I(M_this_vga_ramdac_en_0));
    LocalMux I__1137 (
            .O(N__9345),
            .I(M_this_vga_ramdac_en_0));
    LocalMux I__1136 (
            .O(N__9342),
            .I(M_this_vga_ramdac_en_0));
    CascadeMux I__1135 (
            .O(N__9335),
            .I(\this_vga_signals.g0_7_0_0_cascade_ ));
    InMux I__1134 (
            .O(N__9332),
            .I(N__9329));
    LocalMux I__1133 (
            .O(N__9329),
            .I(N__9326));
    Span4Mux_v I__1132 (
            .O(N__9326),
            .I(N__9323));
    Odrv4 I__1131 (
            .O(N__9323),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i_0_1_0 ));
    InMux I__1130 (
            .O(N__9320),
            .I(N__9314));
    InMux I__1129 (
            .O(N__9319),
            .I(N__9314));
    LocalMux I__1128 (
            .O(N__9314),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ));
    InMux I__1127 (
            .O(N__9311),
            .I(N__9304));
    InMux I__1126 (
            .O(N__9310),
            .I(N__9304));
    InMux I__1125 (
            .O(N__9309),
            .I(N__9301));
    LocalMux I__1124 (
            .O(N__9304),
            .I(\this_vga_signals.SUM_2_i_1_2_3 ));
    LocalMux I__1123 (
            .O(N__9301),
            .I(\this_vga_signals.SUM_2_i_1_2_3 ));
    CascadeMux I__1122 (
            .O(N__9296),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i_0_0_cascade_ ));
    InMux I__1121 (
            .O(N__9293),
            .I(N__9286));
    InMux I__1120 (
            .O(N__9292),
            .I(N__9286));
    InMux I__1119 (
            .O(N__9291),
            .I(N__9283));
    LocalMux I__1118 (
            .O(N__9286),
            .I(\this_vga_signals.SUM_2_i_1_0_3 ));
    LocalMux I__1117 (
            .O(N__9283),
            .I(\this_vga_signals.SUM_2_i_1_0_3 ));
    CascadeMux I__1116 (
            .O(N__9278),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_ ));
    InMux I__1115 (
            .O(N__9275),
            .I(N__9269));
    InMux I__1114 (
            .O(N__9274),
            .I(N__9266));
    InMux I__1113 (
            .O(N__9273),
            .I(N__9261));
    InMux I__1112 (
            .O(N__9272),
            .I(N__9261));
    LocalMux I__1111 (
            .O(N__9269),
            .I(N__9258));
    LocalMux I__1110 (
            .O(N__9266),
            .I(N__9255));
    LocalMux I__1109 (
            .O(N__9261),
            .I(N__9252));
    Span4Mux_v I__1108 (
            .O(N__9258),
            .I(N__9247));
    Span4Mux_h I__1107 (
            .O(N__9255),
            .I(N__9247));
    Span4Mux_h I__1106 (
            .O(N__9252),
            .I(N__9244));
    Odrv4 I__1105 (
            .O(N__9247),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_2 ));
    Odrv4 I__1104 (
            .O(N__9244),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_3_2 ));
    InMux I__1103 (
            .O(N__9239),
            .I(N__9236));
    LocalMux I__1102 (
            .O(N__9236),
            .I(N__9232));
    InMux I__1101 (
            .O(N__9235),
            .I(N__9229));
    Odrv12 I__1100 (
            .O(N__9232),
            .I(\this_vga_signals.N_3_2_1 ));
    LocalMux I__1099 (
            .O(N__9229),
            .I(\this_vga_signals.N_3_2_1 ));
    CascadeMux I__1098 (
            .O(N__9224),
            .I(\this_vga_signals.N_3_2_1_cascade_ ));
    InMux I__1097 (
            .O(N__9221),
            .I(N__9217));
    InMux I__1096 (
            .O(N__9220),
            .I(N__9214));
    LocalMux I__1095 (
            .O(N__9217),
            .I(N__9211));
    LocalMux I__1094 (
            .O(N__9214),
            .I(N__9208));
    Sp12to4 I__1093 (
            .O(N__9211),
            .I(N__9203));
    Span4Mux_h I__1092 (
            .O(N__9208),
            .I(N__9200));
    InMux I__1091 (
            .O(N__9207),
            .I(N__9197));
    InMux I__1090 (
            .O(N__9206),
            .I(N__9194));
    Odrv12 I__1089 (
            .O(N__9203),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    Odrv4 I__1088 (
            .O(N__9200),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1087 (
            .O(N__9197),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1086 (
            .O(N__9194),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    InMux I__1085 (
            .O(N__9185),
            .I(N__9180));
    InMux I__1084 (
            .O(N__9184),
            .I(N__9175));
    InMux I__1083 (
            .O(N__9183),
            .I(N__9175));
    LocalMux I__1082 (
            .O(N__9180),
            .I(\this_vga_signals.mult1_un68_sum_axb2_1 ));
    LocalMux I__1081 (
            .O(N__9175),
            .I(\this_vga_signals.mult1_un68_sum_axb2_1 ));
    CascadeMux I__1080 (
            .O(N__9170),
            .I(\this_vga_signals.mult1_un68_sum_axb2_1_cascade_ ));
    InMux I__1079 (
            .O(N__9167),
            .I(N__9161));
    InMux I__1078 (
            .O(N__9166),
            .I(N__9156));
    InMux I__1077 (
            .O(N__9165),
            .I(N__9156));
    InMux I__1076 (
            .O(N__9164),
            .I(N__9153));
    LocalMux I__1075 (
            .O(N__9161),
            .I(N__9150));
    LocalMux I__1074 (
            .O(N__9156),
            .I(N__9147));
    LocalMux I__1073 (
            .O(N__9153),
            .I(N__9144));
    Span4Mux_v I__1072 (
            .O(N__9150),
            .I(N__9141));
    Span4Mux_h I__1071 (
            .O(N__9147),
            .I(N__9138));
    Odrv12 I__1070 (
            .O(N__9144),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    Odrv4 I__1069 (
            .O(N__9141),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    Odrv4 I__1068 (
            .O(N__9138),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    InMux I__1067 (
            .O(N__9131),
            .I(N__9128));
    LocalMux I__1066 (
            .O(N__9128),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1 ));
    CascadeMux I__1065 (
            .O(N__9125),
            .I(N__9122));
    InMux I__1064 (
            .O(N__9122),
            .I(N__9118));
    InMux I__1063 (
            .O(N__9121),
            .I(N__9115));
    LocalMux I__1062 (
            .O(N__9118),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ));
    LocalMux I__1061 (
            .O(N__9115),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ));
    InMux I__1060 (
            .O(N__9110),
            .I(N__9107));
    LocalMux I__1059 (
            .O(N__9107),
            .I(N__9104));
    Span4Mux_v I__1058 (
            .O(N__9104),
            .I(N__9100));
    InMux I__1057 (
            .O(N__9103),
            .I(N__9097));
    Span4Mux_v I__1056 (
            .O(N__9100),
            .I(N__9094));
    LocalMux I__1055 (
            .O(N__9097),
            .I(N__9088));
    Sp12to4 I__1054 (
            .O(N__9094),
            .I(N__9083));
    InMux I__1053 (
            .O(N__9093),
            .I(N__9076));
    InMux I__1052 (
            .O(N__9092),
            .I(N__9076));
    InMux I__1051 (
            .O(N__9091),
            .I(N__9076));
    Span4Mux_v I__1050 (
            .O(N__9088),
            .I(N__9073));
    InMux I__1049 (
            .O(N__9087),
            .I(N__9070));
    InMux I__1048 (
            .O(N__9086),
            .I(N__9067));
    Odrv12 I__1047 (
            .O(N__9083),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1046 (
            .O(N__9076),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    Odrv4 I__1045 (
            .O(N__9073),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1044 (
            .O(N__9070),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1043 (
            .O(N__9067),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    CascadeMux I__1042 (
            .O(N__9056),
            .I(\this_vga_signals.SUM_3_i_0_0_3_cascade_ ));
    InMux I__1041 (
            .O(N__9053),
            .I(N__9050));
    LocalMux I__1040 (
            .O(N__9050),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_0 ));
    InMux I__1039 (
            .O(N__9047),
            .I(N__9044));
    LocalMux I__1038 (
            .O(N__9044),
            .I(\this_vga_signals.vaddress_1_5 ));
    CascadeMux I__1037 (
            .O(N__9041),
            .I(\this_vga_signals.vaddress_1_6_cascade_ ));
    InMux I__1036 (
            .O(N__9038),
            .I(N__9035));
    LocalMux I__1035 (
            .O(N__9035),
            .I(\this_vga_signals.mult1_un54_sum_axb1_1_0_1 ));
    CascadeMux I__1034 (
            .O(N__9032),
            .I(N__9022));
    CascadeMux I__1033 (
            .O(N__9031),
            .I(N__9016));
    CascadeMux I__1032 (
            .O(N__9030),
            .I(N__9013));
    CascadeMux I__1031 (
            .O(N__9029),
            .I(N__9009));
    InMux I__1030 (
            .O(N__9028),
            .I(N__9002));
    InMux I__1029 (
            .O(N__9027),
            .I(N__8997));
    InMux I__1028 (
            .O(N__9026),
            .I(N__8997));
    InMux I__1027 (
            .O(N__9025),
            .I(N__8990));
    InMux I__1026 (
            .O(N__9022),
            .I(N__8990));
    InMux I__1025 (
            .O(N__9021),
            .I(N__8990));
    InMux I__1024 (
            .O(N__9020),
            .I(N__8981));
    InMux I__1023 (
            .O(N__9019),
            .I(N__8981));
    InMux I__1022 (
            .O(N__9016),
            .I(N__8981));
    InMux I__1021 (
            .O(N__9013),
            .I(N__8981));
    InMux I__1020 (
            .O(N__9012),
            .I(N__8976));
    InMux I__1019 (
            .O(N__9009),
            .I(N__8976));
    InMux I__1018 (
            .O(N__9008),
            .I(N__8967));
    InMux I__1017 (
            .O(N__9007),
            .I(N__8967));
    InMux I__1016 (
            .O(N__9006),
            .I(N__8967));
    InMux I__1015 (
            .O(N__9005),
            .I(N__8967));
    LocalMux I__1014 (
            .O(N__9002),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1013 (
            .O(N__8997),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1012 (
            .O(N__8990),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1011 (
            .O(N__8981),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1010 (
            .O(N__8976),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1009 (
            .O(N__8967),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    InMux I__1008 (
            .O(N__8954),
            .I(N__8951));
    LocalMux I__1007 (
            .O(N__8951),
            .I(\this_vga_signals.g0_12_x1 ));
    CascadeMux I__1006 (
            .O(N__8948),
            .I(\this_vga_signals.g0_0_2_1_0_cascade_ ));
    InMux I__1005 (
            .O(N__8945),
            .I(N__8942));
    LocalMux I__1004 (
            .O(N__8942),
            .I(N__8939));
    Odrv4 I__1003 (
            .O(N__8939),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_0 ));
    InMux I__1002 (
            .O(N__8936),
            .I(N__8932));
    InMux I__1001 (
            .O(N__8935),
            .I(N__8929));
    LocalMux I__1000 (
            .O(N__8932),
            .I(\this_vga_signals.g0_0_2 ));
    LocalMux I__999 (
            .O(N__8929),
            .I(\this_vga_signals.g0_0_2 ));
    CascadeMux I__998 (
            .O(N__8924),
            .I(N__8921));
    InMux I__997 (
            .O(N__8921),
            .I(N__8917));
    InMux I__996 (
            .O(N__8920),
            .I(N__8914));
    LocalMux I__995 (
            .O(N__8917),
            .I(N__8911));
    LocalMux I__994 (
            .O(N__8914),
            .I(\this_vga_signals.vaddress_6_5 ));
    Odrv4 I__993 (
            .O(N__8911),
            .I(\this_vga_signals.vaddress_6_5 ));
    CascadeMux I__992 (
            .O(N__8906),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_1_0_cascade_ ));
    InMux I__991 (
            .O(N__8903),
            .I(N__8900));
    LocalMux I__990 (
            .O(N__8900),
            .I(N__8897));
    Odrv4 I__989 (
            .O(N__8897),
            .I(\this_vga_signals.g0_0_2_0 ));
    InMux I__988 (
            .O(N__8894),
            .I(N__8891));
    LocalMux I__987 (
            .O(N__8891),
            .I(\this_vga_signals.N_236 ));
    CascadeMux I__986 (
            .O(N__8888),
            .I(\this_vga_signals.mult1_un68_sum_axb1_395_cascade_ ));
    InMux I__985 (
            .O(N__8885),
            .I(N__8882));
    LocalMux I__984 (
            .O(N__8882),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0 ));
    InMux I__983 (
            .O(N__8879),
            .I(N__8876));
    LocalMux I__982 (
            .O(N__8876),
            .I(N__8869));
    InMux I__981 (
            .O(N__8875),
            .I(N__8864));
    InMux I__980 (
            .O(N__8874),
            .I(N__8864));
    InMux I__979 (
            .O(N__8873),
            .I(N__8859));
    InMux I__978 (
            .O(N__8872),
            .I(N__8859));
    Odrv4 I__977 (
            .O(N__8869),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__976 (
            .O(N__8864),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    LocalMux I__975 (
            .O(N__8859),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    CascadeMux I__974 (
            .O(N__8852),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_cascade_ ));
    CascadeMux I__973 (
            .O(N__8849),
            .I(\this_vga_signals.g0_5_2_cascade_ ));
    InMux I__972 (
            .O(N__8846),
            .I(N__8843));
    LocalMux I__971 (
            .O(N__8843),
            .I(\this_vga_signals.g1_2 ));
    InMux I__970 (
            .O(N__8840),
            .I(N__8837));
    LocalMux I__969 (
            .O(N__8837),
            .I(\this_vga_signals.mult1_un68_sum_ac0_1_x1 ));
    InMux I__968 (
            .O(N__8834),
            .I(N__8831));
    LocalMux I__967 (
            .O(N__8831),
            .I(\this_vga_signals.mult1_un68_sum_ac0_1 ));
    InMux I__966 (
            .O(N__8828),
            .I(N__8825));
    LocalMux I__965 (
            .O(N__8825),
            .I(\this_vga_signals.N_3_1 ));
    InMux I__964 (
            .O(N__8822),
            .I(N__8819));
    LocalMux I__963 (
            .O(N__8819),
            .I(\this_vga_signals.N_7 ));
    CascadeMux I__962 (
            .O(N__8816),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_cascade_ ));
    InMux I__961 (
            .O(N__8813),
            .I(N__8810));
    LocalMux I__960 (
            .O(N__8810),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_0_0 ));
    InMux I__959 (
            .O(N__8807),
            .I(N__8804));
    LocalMux I__958 (
            .O(N__8804),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    CascadeMux I__957 (
            .O(N__8801),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_ ));
    CascadeMux I__956 (
            .O(N__8798),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4_cascade_ ));
    InMux I__955 (
            .O(N__8795),
            .I(N__8792));
    LocalMux I__954 (
            .O(N__8792),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    CascadeMux I__953 (
            .O(N__8789),
            .I(\this_vga_signals.N_1_4_1_cascade_ ));
    CascadeMux I__952 (
            .O(N__8786),
            .I(\this_vga_signals.M_pcounter_q_3_0_cascade_ ));
    InMux I__951 (
            .O(N__8783),
            .I(N__8777));
    InMux I__950 (
            .O(N__8782),
            .I(N__8777));
    LocalMux I__949 (
            .O(N__8777),
            .I(N__8774));
    Span4Mux_h I__948 (
            .O(N__8774),
            .I(N__8771));
    Odrv4 I__947 (
            .O(N__8771),
            .I(\this_vga_signals.N_2_0 ));
    CascadeMux I__946 (
            .O(N__8768),
            .I(\this_vga_signals.N_2_0_cascade_ ));
    InMux I__945 (
            .O(N__8765),
            .I(N__8761));
    InMux I__944 (
            .O(N__8764),
            .I(N__8758));
    LocalMux I__943 (
            .O(N__8761),
            .I(\this_vga_signals.M_pcounter_q_i_3_0 ));
    LocalMux I__942 (
            .O(N__8758),
            .I(\this_vga_signals.M_pcounter_q_i_3_0 ));
    InMux I__941 (
            .O(N__8753),
            .I(N__8747));
    InMux I__940 (
            .O(N__8752),
            .I(N__8747));
    LocalMux I__939 (
            .O(N__8747),
            .I(N__8743));
    InMux I__938 (
            .O(N__8746),
            .I(N__8740));
    Span4Mux_h I__937 (
            .O(N__8743),
            .I(N__8737));
    LocalMux I__936 (
            .O(N__8740),
            .I(\this_vga_signals.N_3_0 ));
    Odrv4 I__935 (
            .O(N__8737),
            .I(\this_vga_signals.N_3_0 ));
    InMux I__934 (
            .O(N__8732),
            .I(N__8725));
    InMux I__933 (
            .O(N__8731),
            .I(N__8725));
    InMux I__932 (
            .O(N__8730),
            .I(N__8722));
    LocalMux I__931 (
            .O(N__8725),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    LocalMux I__930 (
            .O(N__8722),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    CascadeMux I__929 (
            .O(N__8717),
            .I(N__8714));
    InMux I__928 (
            .O(N__8714),
            .I(N__8709));
    InMux I__927 (
            .O(N__8713),
            .I(N__8704));
    InMux I__926 (
            .O(N__8712),
            .I(N__8704));
    LocalMux I__925 (
            .O(N__8709),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    LocalMux I__924 (
            .O(N__8704),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    CascadeMux I__923 (
            .O(N__8699),
            .I(N__8694));
    InMux I__922 (
            .O(N__8698),
            .I(N__8688));
    InMux I__921 (
            .O(N__8697),
            .I(N__8688));
    InMux I__920 (
            .O(N__8694),
            .I(N__8683));
    InMux I__919 (
            .O(N__8693),
            .I(N__8683));
    LocalMux I__918 (
            .O(N__8688),
            .I(\this_vga_signals.M_pcounter_q_i_3_1 ));
    LocalMux I__917 (
            .O(N__8683),
            .I(\this_vga_signals.M_pcounter_q_i_3_1 ));
    InMux I__916 (
            .O(N__8678),
            .I(N__8675));
    LocalMux I__915 (
            .O(N__8675),
            .I(\this_vga_signals.M_pcounter_q_3_1 ));
    CascadeMux I__914 (
            .O(N__8672),
            .I(N__8669));
    InMux I__913 (
            .O(N__8669),
            .I(N__8666));
    LocalMux I__912 (
            .O(N__8666),
            .I(N__8663));
    Span4Mux_h I__911 (
            .O(N__8663),
            .I(N__8660));
    Span4Mux_v I__910 (
            .O(N__8660),
            .I(N__8657));
    Odrv4 I__909 (
            .O(N__8657),
            .I(M_this_vga_signals_address_6));
    CascadeMux I__908 (
            .O(N__8654),
            .I(N__8651));
    InMux I__907 (
            .O(N__8651),
            .I(N__8648));
    LocalMux I__906 (
            .O(N__8648),
            .I(N__8645));
    Span4Mux_v I__905 (
            .O(N__8645),
            .I(N__8640));
    InMux I__904 (
            .O(N__8644),
            .I(N__8635));
    InMux I__903 (
            .O(N__8643),
            .I(N__8635));
    Odrv4 I__902 (
            .O(N__8640),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    LocalMux I__901 (
            .O(N__8635),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    CascadeMux I__900 (
            .O(N__8630),
            .I(N__8627));
    InMux I__899 (
            .O(N__8627),
            .I(N__8624));
    LocalMux I__898 (
            .O(N__8624),
            .I(N__8621));
    Span4Mux_h I__897 (
            .O(N__8621),
            .I(N__8618));
    Span4Mux_v I__896 (
            .O(N__8618),
            .I(N__8615));
    Odrv4 I__895 (
            .O(N__8615),
            .I(M_this_vga_signals_address_3));
    InMux I__894 (
            .O(N__8612),
            .I(N__8609));
    LocalMux I__893 (
            .O(N__8609),
            .I(N__8606));
    Span4Mux_v I__892 (
            .O(N__8606),
            .I(N__8603));
    Odrv4 I__891 (
            .O(N__8603),
            .I(\this_vga_signals.vaddress_1_0_6 ));
    CascadeMux I__890 (
            .O(N__8600),
            .I(\this_vga_signals.g1_2_0_cascade_ ));
    InMux I__889 (
            .O(N__8597),
            .I(N__8594));
    LocalMux I__888 (
            .O(N__8594),
            .I(N__8591));
    Odrv12 I__887 (
            .O(N__8591),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2_0_0 ));
    CascadeMux I__886 (
            .O(N__8588),
            .I(N__8585));
    InMux I__885 (
            .O(N__8585),
            .I(N__8582));
    LocalMux I__884 (
            .O(N__8582),
            .I(N__8579));
    Odrv12 I__883 (
            .O(N__8579),
            .I(\this_vga_signals.g1_3 ));
    CascadeMux I__882 (
            .O(N__8576),
            .I(N__8573));
    InMux I__881 (
            .O(N__8573),
            .I(N__8570));
    LocalMux I__880 (
            .O(N__8570),
            .I(N__8567));
    Span4Mux_h I__879 (
            .O(N__8567),
            .I(N__8564));
    Odrv4 I__878 (
            .O(N__8564),
            .I(\this_vga_signals.M_hcounter_q_RNI8OIBAZ0Z_3 ));
    CascadeMux I__877 (
            .O(N__8561),
            .I(N__8557));
    InMux I__876 (
            .O(N__8560),
            .I(N__8554));
    InMux I__875 (
            .O(N__8557),
            .I(N__8551));
    LocalMux I__874 (
            .O(N__8554),
            .I(N__8548));
    LocalMux I__873 (
            .O(N__8551),
            .I(N__8545));
    Span4Mux_v I__872 (
            .O(N__8548),
            .I(N__8542));
    Span4Mux_h I__871 (
            .O(N__8545),
            .I(N__8539));
    Odrv4 I__870 (
            .O(N__8542),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    Odrv4 I__869 (
            .O(N__8539),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    InMux I__868 (
            .O(N__8534),
            .I(N__8531));
    LocalMux I__867 (
            .O(N__8531),
            .I(N__8528));
    Span4Mux_h I__866 (
            .O(N__8528),
            .I(N__8525));
    Odrv4 I__865 (
            .O(N__8525),
            .I(\this_vga_signals.if_N_8_i_0 ));
    CascadeMux I__864 (
            .O(N__8522),
            .I(\this_vga_signals.g0_9_1_cascade_ ));
    InMux I__863 (
            .O(N__8519),
            .I(N__8516));
    LocalMux I__862 (
            .O(N__8516),
            .I(\this_vga_signals.g0_12_x0 ));
    InMux I__861 (
            .O(N__8513),
            .I(N__8510));
    LocalMux I__860 (
            .O(N__8510),
            .I(\this_vga_signals.g0_5_0 ));
    CascadeMux I__859 (
            .O(N__8507),
            .I(\this_vga_signals.N_6_0_cascade_ ));
    InMux I__858 (
            .O(N__8504),
            .I(N__8501));
    LocalMux I__857 (
            .O(N__8501),
            .I(\this_vga_signals.N_5 ));
    InMux I__856 (
            .O(N__8498),
            .I(N__8495));
    LocalMux I__855 (
            .O(N__8495),
            .I(N__8492));
    Odrv12 I__854 (
            .O(N__8492),
            .I(\this_vga_signals.d_N_3_i_0_0_0 ));
    InMux I__853 (
            .O(N__8489),
            .I(N__8486));
    LocalMux I__852 (
            .O(N__8486),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ));
    CascadeMux I__851 (
            .O(N__8483),
            .I(\this_vga_signals.g0_3_cascade_ ));
    InMux I__850 (
            .O(N__8480),
            .I(N__8476));
    InMux I__849 (
            .O(N__8479),
            .I(N__8473));
    LocalMux I__848 (
            .O(N__8476),
            .I(\this_vga_signals.mult1_un68_sum_axb1 ));
    LocalMux I__847 (
            .O(N__8473),
            .I(\this_vga_signals.mult1_un68_sum_axb1 ));
    CascadeMux I__846 (
            .O(N__8468),
            .I(\this_vga_signals.N_5_1_cascade_ ));
    InMux I__845 (
            .O(N__8465),
            .I(N__8462));
    LocalMux I__844 (
            .O(N__8462),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0 ));
    CascadeMux I__843 (
            .O(N__8459),
            .I(\this_vga_signals.if_i1_mux_0_cascade_ ));
    InMux I__842 (
            .O(N__8456),
            .I(N__8453));
    LocalMux I__841 (
            .O(N__8453),
            .I(\this_vga_signals.g1_6_0 ));
    InMux I__840 (
            .O(N__8450),
            .I(N__8447));
    LocalMux I__839 (
            .O(N__8447),
            .I(\this_vga_signals.mult1_un75_sum_c3_0_0 ));
    InMux I__838 (
            .O(N__8444),
            .I(N__8441));
    LocalMux I__837 (
            .O(N__8441),
            .I(\this_vga_signals.if_m1_3 ));
    InMux I__836 (
            .O(N__8438),
            .I(N__8435));
    LocalMux I__835 (
            .O(N__8435),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3 ));
    CascadeMux I__834 (
            .O(N__8432),
            .I(\this_vga_signals.if_m1_3_cascade_ ));
    InMux I__833 (
            .O(N__8429),
            .I(N__8425));
    InMux I__832 (
            .O(N__8428),
            .I(N__8422));
    LocalMux I__831 (
            .O(N__8425),
            .I(\this_vga_signals.mult1_un68_sum_axbxc2 ));
    LocalMux I__830 (
            .O(N__8422),
            .I(\this_vga_signals.mult1_un68_sum_axbxc2 ));
    CascadeMux I__829 (
            .O(N__8417),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ));
    InMux I__828 (
            .O(N__8414),
            .I(N__8411));
    LocalMux I__827 (
            .O(N__8411),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_i ));
    CascadeMux I__826 (
            .O(N__8408),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_i_cascade_ ));
    InMux I__825 (
            .O(N__8405),
            .I(N__8402));
    LocalMux I__824 (
            .O(N__8402),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0 ));
    InMux I__823 (
            .O(N__8399),
            .I(N__8396));
    LocalMux I__822 (
            .O(N__8396),
            .I(\this_vga_signals.if_N_2_1_0_0 ));
    InMux I__821 (
            .O(N__8393),
            .I(N__8390));
    LocalMux I__820 (
            .O(N__8390),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1 ));
    CascadeMux I__819 (
            .O(N__8387),
            .I(\this_vga_signals.vaddress_1_0_5_cascade_ ));
    CascadeMux I__818 (
            .O(N__8384),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_cascade_ ));
    CascadeMux I__817 (
            .O(N__8381),
            .I(N__8378));
    InMux I__816 (
            .O(N__8378),
            .I(N__8375));
    LocalMux I__815 (
            .O(N__8375),
            .I(N__8372));
    Span4Mux_v I__814 (
            .O(N__8372),
            .I(N__8369));
    Span4Mux_v I__813 (
            .O(N__8369),
            .I(N__8366));
    Odrv4 I__812 (
            .O(N__8366),
            .I(M_this_vga_signals_address_7));
    CascadeMux I__811 (
            .O(N__8363),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_cascade_ ));
    CascadeMux I__810 (
            .O(N__8360),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_cascade_ ));
    CascadeMux I__809 (
            .O(N__8357),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_cascade_ ));
    InMux I__808 (
            .O(N__8354),
            .I(N__8351));
    LocalMux I__807 (
            .O(N__8351),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_0 ));
    CascadeMux I__806 (
            .O(N__8348),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_cascade_ ));
    InMux I__805 (
            .O(N__8345),
            .I(N__8342));
    LocalMux I__804 (
            .O(N__8342),
            .I(\this_vga_signals.mult1_un89_sum_c3 ));
    CascadeMux I__803 (
            .O(N__8339),
            .I(N__8336));
    InMux I__802 (
            .O(N__8336),
            .I(N__8333));
    LocalMux I__801 (
            .O(N__8333),
            .I(N__8330));
    Span4Mux_v I__800 (
            .O(N__8330),
            .I(N__8327));
    Span4Mux_v I__799 (
            .O(N__8327),
            .I(N__8324));
    Odrv4 I__798 (
            .O(N__8324),
            .I(M_this_vga_signals_address_0));
    InMux I__797 (
            .O(N__8321),
            .I(N__8311));
    InMux I__796 (
            .O(N__8320),
            .I(N__8311));
    InMux I__795 (
            .O(N__8319),
            .I(N__8308));
    InMux I__794 (
            .O(N__8318),
            .I(N__8301));
    InMux I__793 (
            .O(N__8317),
            .I(N__8301));
    InMux I__792 (
            .O(N__8316),
            .I(N__8301));
    LocalMux I__791 (
            .O(N__8311),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    LocalMux I__790 (
            .O(N__8308),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    LocalMux I__789 (
            .O(N__8301),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    InMux I__788 (
            .O(N__8294),
            .I(N__8291));
    LocalMux I__787 (
            .O(N__8291),
            .I(\this_vga_signals.d_N_11 ));
    InMux I__786 (
            .O(N__8288),
            .I(N__8285));
    LocalMux I__785 (
            .O(N__8285),
            .I(\this_vga_signals.d_N_12 ));
    CascadeMux I__784 (
            .O(N__8282),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_cascade_ ));
    InMux I__783 (
            .O(N__8279),
            .I(N__8273));
    InMux I__782 (
            .O(N__8278),
            .I(N__8273));
    LocalMux I__781 (
            .O(N__8273),
            .I(\this_vga_signals.mult1_un75_sum_axb1 ));
    InMux I__780 (
            .O(N__8270),
            .I(N__8265));
    InMux I__779 (
            .O(N__8269),
            .I(N__8262));
    CascadeMux I__778 (
            .O(N__8268),
            .I(N__8259));
    LocalMux I__777 (
            .O(N__8265),
            .I(N__8253));
    LocalMux I__776 (
            .O(N__8262),
            .I(N__8253));
    InMux I__775 (
            .O(N__8259),
            .I(N__8248));
    InMux I__774 (
            .O(N__8258),
            .I(N__8248));
    Odrv4 I__773 (
            .O(N__8253),
            .I(\this_vga_signals.mult1_un68_sum_axbxc1 ));
    LocalMux I__772 (
            .O(N__8248),
            .I(\this_vga_signals.mult1_un68_sum_axbxc1 ));
    CascadeMux I__771 (
            .O(N__8243),
            .I(N__8240));
    InMux I__770 (
            .O(N__8240),
            .I(N__8237));
    LocalMux I__769 (
            .O(N__8237),
            .I(N__8234));
    Odrv4 I__768 (
            .O(N__8234),
            .I(M_this_vga_signals_address_5));
    CascadeMux I__767 (
            .O(N__8231),
            .I(N__8228));
    InMux I__766 (
            .O(N__8228),
            .I(N__8225));
    LocalMux I__765 (
            .O(N__8225),
            .I(M_this_vga_signals_address_4));
    CascadeMux I__764 (
            .O(N__8222),
            .I(\this_vga_signals.if_N_9_1_cascade_ ));
    InMux I__763 (
            .O(N__8219),
            .I(N__8216));
    LocalMux I__762 (
            .O(N__8216),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1 ));
    CascadeMux I__761 (
            .O(N__8213),
            .I(\this_vga_signals.if_m1_0_cascade_ ));
    CascadeMux I__760 (
            .O(N__8210),
            .I(\this_vga_signals.mult1_un82_sum_c3_cascade_ ));
    InMux I__759 (
            .O(N__8207),
            .I(N__8204));
    LocalMux I__758 (
            .O(N__8204),
            .I(\this_vga_signals.N_2_7_0 ));
    InMux I__757 (
            .O(N__8201),
            .I(N__8197));
    InMux I__756 (
            .O(N__8200),
            .I(N__8194));
    LocalMux I__755 (
            .O(N__8197),
            .I(\this_vga_signals.mult1_un75_sum_c2_0 ));
    LocalMux I__754 (
            .O(N__8194),
            .I(\this_vga_signals.mult1_un75_sum_c2_0 ));
    InMux I__753 (
            .O(N__8189),
            .I(N__8186));
    LocalMux I__752 (
            .O(N__8186),
            .I(N__8183));
    Span4Mux_h I__751 (
            .O(N__8183),
            .I(N__8180));
    Span4Mux_v I__750 (
            .O(N__8180),
            .I(N__8174));
    InMux I__749 (
            .O(N__8179),
            .I(N__8169));
    InMux I__748 (
            .O(N__8178),
            .I(N__8169));
    InMux I__747 (
            .O(N__8177),
            .I(N__8166));
    Odrv4 I__746 (
            .O(N__8174),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__745 (
            .O(N__8169),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__744 (
            .O(N__8166),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    InMux I__743 (
            .O(N__8159),
            .I(N__8155));
    InMux I__742 (
            .O(N__8158),
            .I(N__8152));
    LocalMux I__741 (
            .O(N__8155),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0 ));
    LocalMux I__740 (
            .O(N__8152),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0 ));
    InMux I__739 (
            .O(N__8147),
            .I(N__8144));
    LocalMux I__738 (
            .O(N__8144),
            .I(N__8141));
    Odrv12 I__737 (
            .O(N__8141),
            .I(\this_vga_ramdac.m19 ));
    InMux I__736 (
            .O(N__8138),
            .I(N__8134));
    CascadeMux I__735 (
            .O(N__8137),
            .I(N__8131));
    LocalMux I__734 (
            .O(N__8134),
            .I(N__8128));
    InMux I__733 (
            .O(N__8131),
            .I(N__8125));
    Odrv12 I__732 (
            .O(N__8128),
            .I(\this_vga_ramdac.N_1766_reto ));
    LocalMux I__731 (
            .O(N__8125),
            .I(\this_vga_ramdac.N_1766_reto ));
    InMux I__730 (
            .O(N__8120),
            .I(N__8117));
    LocalMux I__729 (
            .O(N__8117),
            .I(\this_vga_signals.M_this_vga_signals_pixel_clk_0_0 ));
    CascadeMux I__728 (
            .O(N__8114),
            .I(N__8108));
    CascadeMux I__727 (
            .O(N__8113),
            .I(N__8105));
    InMux I__726 (
            .O(N__8112),
            .I(N__8092));
    InMux I__725 (
            .O(N__8111),
            .I(N__8092));
    InMux I__724 (
            .O(N__8108),
            .I(N__8092));
    InMux I__723 (
            .O(N__8105),
            .I(N__8092));
    InMux I__722 (
            .O(N__8104),
            .I(N__8092));
    InMux I__721 (
            .O(N__8103),
            .I(N__8089));
    LocalMux I__720 (
            .O(N__8092),
            .I(M_pcounter_q_ret_2_RNIRAOL5));
    LocalMux I__719 (
            .O(N__8089),
            .I(M_pcounter_q_ret_2_RNIRAOL5));
    CascadeMux I__718 (
            .O(N__8084),
            .I(M_pcounter_q_ret_2_RNIRAOL5_cascade_));
    InMux I__717 (
            .O(N__8081),
            .I(N__8078));
    LocalMux I__716 (
            .O(N__8078),
            .I(N__8075));
    Odrv12 I__715 (
            .O(N__8075),
            .I(\this_vga_ramdac.i2_mux_0 ));
    InMux I__714 (
            .O(N__8072),
            .I(N__8069));
    LocalMux I__713 (
            .O(N__8069),
            .I(N__8066));
    Span4Mux_v I__712 (
            .O(N__8066),
            .I(N__8062));
    InMux I__711 (
            .O(N__8065),
            .I(N__8059));
    Odrv4 I__710 (
            .O(N__8062),
            .I(\this_vga_ramdac.N_1767_reto ));
    LocalMux I__709 (
            .O(N__8059),
            .I(\this_vga_ramdac.N_1767_reto ));
    InMux I__708 (
            .O(N__8054),
            .I(N__8051));
    LocalMux I__707 (
            .O(N__8051),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    CascadeMux I__706 (
            .O(N__8048),
            .I(N__8045));
    InMux I__705 (
            .O(N__8045),
            .I(N__8042));
    LocalMux I__704 (
            .O(N__8042),
            .I(N__8039));
    Odrv4 I__703 (
            .O(N__8039),
            .I(M_this_vga_signals_address_2));
    CascadeMux I__702 (
            .O(N__8036),
            .I(N__8033));
    InMux I__701 (
            .O(N__8033),
            .I(N__8030));
    LocalMux I__700 (
            .O(N__8030),
            .I(N__8027));
    Span4Mux_v I__699 (
            .O(N__8027),
            .I(N__8024));
    Span4Mux_v I__698 (
            .O(N__8024),
            .I(N__8021));
    Odrv4 I__697 (
            .O(N__8021),
            .I(M_this_vga_signals_address_1));
    CascadeMux I__696 (
            .O(N__8018),
            .I(\this_vga_signals.mult1_un75_sum_c2_0_cascade_ ));
    InMux I__695 (
            .O(N__8015),
            .I(N__8012));
    LocalMux I__694 (
            .O(N__8012),
            .I(\this_vga_signals.if_m7_0_x4_0 ));
    InMux I__693 (
            .O(N__8009),
            .I(N__8004));
    InMux I__692 (
            .O(N__8008),
            .I(N__7999));
    InMux I__691 (
            .O(N__8007),
            .I(N__7999));
    LocalMux I__690 (
            .O(N__8004),
            .I(N__7994));
    LocalMux I__689 (
            .O(N__7999),
            .I(N__7991));
    InMux I__688 (
            .O(N__7998),
            .I(N__7988));
    CascadeMux I__687 (
            .O(N__7997),
            .I(N__7983));
    Span4Mux_v I__686 (
            .O(N__7994),
            .I(N__7980));
    Span4Mux_v I__685 (
            .O(N__7991),
            .I(N__7977));
    LocalMux I__684 (
            .O(N__7988),
            .I(N__7974));
    InMux I__683 (
            .O(N__7987),
            .I(N__7969));
    InMux I__682 (
            .O(N__7986),
            .I(N__7969));
    InMux I__681 (
            .O(N__7983),
            .I(N__7966));
    Odrv4 I__680 (
            .O(N__7980),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    Odrv4 I__679 (
            .O(N__7977),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    Odrv12 I__678 (
            .O(N__7974),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    LocalMux I__677 (
            .O(N__7969),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    LocalMux I__676 (
            .O(N__7966),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    InMux I__675 (
            .O(N__7955),
            .I(N__7952));
    LocalMux I__674 (
            .O(N__7952),
            .I(N__7949));
    Odrv4 I__673 (
            .O(N__7949),
            .I(\this_vga_ramdac.i2_mux ));
    InMux I__672 (
            .O(N__7946),
            .I(N__7942));
    InMux I__671 (
            .O(N__7945),
            .I(N__7939));
    LocalMux I__670 (
            .O(N__7942),
            .I(\this_vga_ramdac.N_1764_reto ));
    LocalMux I__669 (
            .O(N__7939),
            .I(\this_vga_ramdac.N_1764_reto ));
    InMux I__668 (
            .O(N__7934),
            .I(N__7931));
    LocalMux I__667 (
            .O(N__7931),
            .I(N__7928));
    Odrv4 I__666 (
            .O(N__7928),
            .I(\this_vga_ramdac.m16 ));
    InMux I__665 (
            .O(N__7925),
            .I(N__7922));
    LocalMux I__664 (
            .O(N__7922),
            .I(N__7918));
    CascadeMux I__663 (
            .O(N__7921),
            .I(N__7915));
    Span4Mux_v I__662 (
            .O(N__7918),
            .I(N__7912));
    InMux I__661 (
            .O(N__7915),
            .I(N__7909));
    Odrv4 I__660 (
            .O(N__7912),
            .I(\this_vga_ramdac.N_1765_reto ));
    LocalMux I__659 (
            .O(N__7909),
            .I(\this_vga_ramdac.N_1765_reto ));
    InMux I__658 (
            .O(N__7904),
            .I(N__7901));
    LocalMux I__657 (
            .O(N__7901),
            .I(N__7898));
    Odrv12 I__656 (
            .O(N__7898),
            .I(port_clk_c));
    InMux I__655 (
            .O(N__7895),
            .I(N__7892));
    LocalMux I__654 (
            .O(N__7892),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    InMux I__653 (
            .O(N__7889),
            .I(N__7886));
    LocalMux I__652 (
            .O(N__7886),
            .I(N__7883));
    Odrv4 I__651 (
            .O(N__7883),
            .I(\this_vga_ramdac.N_24_mux ));
    InMux I__650 (
            .O(N__7880),
            .I(N__7876));
    CascadeMux I__649 (
            .O(N__7879),
            .I(N__7873));
    LocalMux I__648 (
            .O(N__7876),
            .I(N__7870));
    InMux I__647 (
            .O(N__7873),
            .I(N__7867));
    Odrv4 I__646 (
            .O(N__7870),
            .I(\this_vga_ramdac.N_1762_reto ));
    LocalMux I__645 (
            .O(N__7867),
            .I(\this_vga_ramdac.N_1762_reto ));
    InMux I__644 (
            .O(N__7862),
            .I(N__7859));
    LocalMux I__643 (
            .O(N__7859),
            .I(N__7856));
    Odrv4 I__642 (
            .O(N__7856),
            .I(\this_vga_ramdac.m6 ));
    InMux I__641 (
            .O(N__7853),
            .I(N__7849));
    InMux I__640 (
            .O(N__7852),
            .I(N__7846));
    LocalMux I__639 (
            .O(N__7849),
            .I(\this_vga_ramdac.N_1763_reto ));
    LocalMux I__638 (
            .O(N__7846),
            .I(\this_vga_ramdac.N_1763_reto ));
    IoInMux I__637 (
            .O(N__7841),
            .I(N__7838));
    LocalMux I__636 (
            .O(N__7838),
            .I(N__7835));
    Span12Mux_s7_v I__635 (
            .O(N__7835),
            .I(N__7832));
    Odrv12 I__634 (
            .O(N__7832),
            .I(this_vga_signals_vvisibility_i));
    IoInMux I__633 (
            .O(N__7829),
            .I(N__7826));
    LocalMux I__632 (
            .O(N__7826),
            .I(N__7823));
    IoSpan4Mux I__631 (
            .O(N__7823),
            .I(N__7820));
    Span4Mux_s3_h I__630 (
            .O(N__7820),
            .I(N__7817));
    Odrv4 I__629 (
            .O(N__7817),
            .I(rgb_c_2));
    IoInMux I__628 (
            .O(N__7814),
            .I(N__7811));
    LocalMux I__627 (
            .O(N__7811),
            .I(N__7808));
    IoSpan4Mux I__626 (
            .O(N__7808),
            .I(N__7805));
    Span4Mux_s2_h I__625 (
            .O(N__7805),
            .I(N__7802));
    Odrv4 I__624 (
            .O(N__7802),
            .I(rgb_c_1));
    InMux I__623 (
            .O(N__7799),
            .I(N__7787));
    InMux I__622 (
            .O(N__7798),
            .I(N__7787));
    InMux I__621 (
            .O(N__7797),
            .I(N__7787));
    InMux I__620 (
            .O(N__7796),
            .I(N__7787));
    LocalMux I__619 (
            .O(N__7787),
            .I(N__7782));
    InMux I__618 (
            .O(N__7786),
            .I(N__7777));
    InMux I__617 (
            .O(N__7785),
            .I(N__7777));
    Span4Mux_h I__616 (
            .O(N__7782),
            .I(N__7774));
    LocalMux I__615 (
            .O(N__7777),
            .I(N__7771));
    Sp12to4 I__614 (
            .O(N__7774),
            .I(N__7766));
    Span12Mux_s7_h I__613 (
            .O(N__7771),
            .I(N__7766));
    Odrv12 I__612 (
            .O(N__7766),
            .I(M_this_vram_read_data_0));
    InMux I__611 (
            .O(N__7763),
            .I(N__7753));
    InMux I__610 (
            .O(N__7762),
            .I(N__7753));
    InMux I__609 (
            .O(N__7761),
            .I(N__7744));
    InMux I__608 (
            .O(N__7760),
            .I(N__7744));
    InMux I__607 (
            .O(N__7759),
            .I(N__7744));
    InMux I__606 (
            .O(N__7758),
            .I(N__7744));
    LocalMux I__605 (
            .O(N__7753),
            .I(N__7739));
    LocalMux I__604 (
            .O(N__7744),
            .I(N__7739));
    Span4Mux_v I__603 (
            .O(N__7739),
            .I(N__7736));
    Span4Mux_v I__602 (
            .O(N__7736),
            .I(N__7733));
    Odrv4 I__601 (
            .O(N__7733),
            .I(M_this_vram_read_data_3));
    CascadeMux I__600 (
            .O(N__7730),
            .I(N__7723));
    CascadeMux I__599 (
            .O(N__7729),
            .I(N__7720));
    CascadeMux I__598 (
            .O(N__7728),
            .I(N__7717));
    CascadeMux I__597 (
            .O(N__7727),
            .I(N__7714));
    CascadeMux I__596 (
            .O(N__7726),
            .I(N__7711));
    InMux I__595 (
            .O(N__7723),
            .I(N__7706));
    InMux I__594 (
            .O(N__7720),
            .I(N__7706));
    InMux I__593 (
            .O(N__7717),
            .I(N__7703));
    InMux I__592 (
            .O(N__7714),
            .I(N__7698));
    InMux I__591 (
            .O(N__7711),
            .I(N__7698));
    LocalMux I__590 (
            .O(N__7706),
            .I(N__7691));
    LocalMux I__589 (
            .O(N__7703),
            .I(N__7691));
    LocalMux I__588 (
            .O(N__7698),
            .I(N__7691));
    Span4Mux_v I__587 (
            .O(N__7691),
            .I(N__7688));
    Span4Mux_v I__586 (
            .O(N__7688),
            .I(N__7685));
    Odrv4 I__585 (
            .O(N__7685),
            .I(M_this_vram_read_data_2));
    InMux I__584 (
            .O(N__7682),
            .I(N__7672));
    InMux I__583 (
            .O(N__7681),
            .I(N__7672));
    InMux I__582 (
            .O(N__7680),
            .I(N__7667));
    InMux I__581 (
            .O(N__7679),
            .I(N__7667));
    InMux I__580 (
            .O(N__7678),
            .I(N__7662));
    InMux I__579 (
            .O(N__7677),
            .I(N__7662));
    LocalMux I__578 (
            .O(N__7672),
            .I(N__7655));
    LocalMux I__577 (
            .O(N__7667),
            .I(N__7655));
    LocalMux I__576 (
            .O(N__7662),
            .I(N__7655));
    Span12Mux_v I__575 (
            .O(N__7655),
            .I(N__7652));
    Odrv12 I__574 (
            .O(N__7652),
            .I(M_this_vram_read_data_1));
    IoInMux I__573 (
            .O(N__7649),
            .I(N__7646));
    LocalMux I__572 (
            .O(N__7646),
            .I(\this_vga_signals.N_340_0 ));
    IoInMux I__571 (
            .O(N__7643),
            .I(N__7640));
    LocalMux I__570 (
            .O(N__7640),
            .I(N_198_i));
    IoInMux I__569 (
            .O(N__7637),
            .I(N__7634));
    LocalMux I__568 (
            .O(N__7634),
            .I(N__7631));
    Span4Mux_s2_h I__567 (
            .O(N__7631),
            .I(N__7628));
    Sp12to4 I__566 (
            .O(N__7628),
            .I(N__7625));
    Span12Mux_v I__565 (
            .O(N__7625),
            .I(N__7622));
    Odrv12 I__564 (
            .O(N__7622),
            .I(rgb_c_0));
    IoInMux I__563 (
            .O(N__7619),
            .I(N__7616));
    LocalMux I__562 (
            .O(N__7616),
            .I(N__7613));
    IoSpan4Mux I__561 (
            .O(N__7613),
            .I(N__7610));
    Span4Mux_s2_h I__560 (
            .O(N__7610),
            .I(N__7607));
    Span4Mux_v I__559 (
            .O(N__7607),
            .I(N__7604));
    Odrv4 I__558 (
            .O(N__7604),
            .I(rgb_c_4));
    IoInMux I__557 (
            .O(N__7601),
            .I(N__7598));
    LocalMux I__556 (
            .O(N__7598),
            .I(N__7595));
    Span4Mux_s3_h I__555 (
            .O(N__7595),
            .I(N__7592));
    Odrv4 I__554 (
            .O(N__7592),
            .I(port_nmib_0_i));
    IoInMux I__553 (
            .O(N__7589),
            .I(N__7586));
    LocalMux I__552 (
            .O(N__7586),
            .I(N__7583));
    Span4Mux_s3_h I__551 (
            .O(N__7583),
            .I(N__7580));
    Odrv4 I__550 (
            .O(N__7580),
            .I(rgb_c_3));
    IoInMux I__549 (
            .O(N__7577),
            .I(N__7574));
    LocalMux I__548 (
            .O(N__7574),
            .I(N__7571));
    Span4Mux_s3_h I__547 (
            .O(N__7571),
            .I(N__7568));
    Span4Mux_v I__546 (
            .O(N__7568),
            .I(N__7565));
    Odrv4 I__545 (
            .O(N__7565),
            .I(rgb_c_5));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_21_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_17_0_));
    defparam IN_MUX_bfv_21_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_18_0_ (
            .carryinitin(\this_ppu.sprites_addr_cry_8 ),
            .carryinitout(bfn_21_18_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(un1_M_this_sprites_address_q_cry_7),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_30_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_30_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_30_23_0_));
    defparam IN_MUX_bfv_30_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_30_24_0_ (
            .carryinitin(un1_M_this_external_address_q_cry_7),
            .carryinitout(bfn_30_24_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_17_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_24_0_ (
            .carryinitin(un1_M_this_data_count_q_cry_7),
            .carryinitout(bfn_17_24_0_));
    defparam IN_MUX_bfv_17_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_25_0_ (
            .carryinitin(un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO),
            .carryinitout(bfn_17_25_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNIRO2H5_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__14996),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_515_g ));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNIADVP5_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__7649),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_340_0_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNI6VB7_3  (
            .USERSIGNALTOGLOBALBUFFER(N__14519),
            .GLOBALBUFFEROUTPUT(M_this_state_q_nss_g_0));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIADVP5_9_LC_1_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIADVP5_9_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIADVP5_9_LC_1_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIADVP5_9_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__14263),
            .in2(_gnd_net_),
            .in3(N__11567),
            .lcout(\this_vga_signals.N_340_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_rw_obuf_RNO_LC_1_22_7.C_ON=1'b0;
    defparam port_data_rw_obuf_RNO_LC_1_22_7.SEQ_MODE=4'b0000;
    defparam port_data_rw_obuf_RNO_LC_1_22_7.LUT_INIT=16'b0101010111111111;
    LogicCell40 port_data_rw_obuf_RNO_LC_1_22_7 (
            .in0(N__14431),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13209),
            .lcout(N_198_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_3_20_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_3_20_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_3_20_5  (
            .in0(N__7880),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7998),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_3_21_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_3_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_3_21_7  (
            .in0(_gnd_net_),
            .in1(N__8138),
            .in2(_gnd_net_),
            .in3(N__8009),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA0384_9_LC_4_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA0384_9_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIA0384_9_LC_4_12_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIA0384_9_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(N__13213),
            .in2(_gnd_net_),
            .in3(N__10055),
            .lcout(port_nmib_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_4_22_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_4_22_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_4_22_2  (
            .in0(N__8007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7925),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_22_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_22_6  (
            .in0(N__8008),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8072),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_0_9_LC_5_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_0_9_LC_5_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_0_9_LC_5_19_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_0_9_LC_5_19_6  (
            .in0(N__10048),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_vvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_5_20_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_5_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_5_20_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_5_20_6  (
            .in0(N__7946),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7987),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_5_20_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_5_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_5_20_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_5_20_7  (
            .in0(N__7986),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7853),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_6_17_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_6_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_6_17_2 .LUT_INIT=16'b0001111100011011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_6_17_2  (
            .in0(N__7763),
            .in1(N__7678),
            .in2(N__7730),
            .in3(N__7786),
            .lcout(\this_vga_ramdac.m6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_6_17_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_6_17_6 .LUT_INIT=16'b0001110100100101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_6_17_6  (
            .in0(N__7762),
            .in1(N__7677),
            .in2(N__7729),
            .in3(N__7785),
            .lcout(\this_vga_ramdac.i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_18_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_18_0 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_18_0  (
            .in0(N__7799),
            .in1(N__7758),
            .in2(_gnd_net_),
            .in3(N__7682),
            .lcout(\this_vga_ramdac.N_24_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_18_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_18_1 .LUT_INIT=16'b0010110101110001;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_18_1  (
            .in0(N__7761),
            .in1(N__7680),
            .in2(N__7726),
            .in3(N__7798),
            .lcout(\this_vga_ramdac.m19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_6_18_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_6_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_6_18_5 .LUT_INIT=16'b0000011101100111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_6_18_5  (
            .in0(N__7759),
            .in1(N__7679),
            .in2(N__7727),
            .in3(N__7796),
            .lcout(\this_vga_ramdac.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_6_18_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_6_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_6_18_6 .LUT_INIT=16'b0100000110110111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_6_18_6  (
            .in0(N__7797),
            .in1(N__7760),
            .in2(N__7728),
            .in3(N__7681),
            .lcout(\this_vga_ramdac.m16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_0_LC_6_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_0_LC_6_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_0_LC_6_19_0 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_x4_0_0_LC_6_19_0  (
            .in0(N__8279),
            .in1(_gnd_net_),
            .in2(N__8268),
            .in3(N__8319),
            .lcout(\this_vga_signals.if_m7_0_x4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_6_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_6_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_6_19_3 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_6_19_3  (
            .in0(N__9762),
            .in1(N__8258),
            .in2(N__9826),
            .in3(N__8278),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_6_20_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_6_20_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_6_20_0 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_q_ret_LC_6_20_0  (
            .in0(N__9401),
            .in1(N__8112),
            .in2(N__7997),
            .in3(N__14524),
            .lcout(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_6_20_1 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_6_20_1 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_6_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_6_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7895),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_6_20_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_6_20_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_6_20_3 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_6_20_3  (
            .in0(N__14522),
            .in1(N__7945),
            .in2(N__8114),
            .in3(N__7955),
            .lcout(\this_vga_ramdac.N_1764_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_6_20_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_6_20_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_6_20_4 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_6_20_4  (
            .in0(N__7934),
            .in1(N__8111),
            .in2(N__7921),
            .in3(N__14523),
            .lcout(\this_vga_ramdac.N_1765_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_6_20_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_6_20_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_6_20_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_6_20_5  (
            .in0(N__7904),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_6_20_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_6_20_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_6_20_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_6_20_6  (
            .in0(N__7889),
            .in1(N__8104),
            .in2(N__7879),
            .in3(N__14520),
            .lcout(\this_vga_ramdac.N_1762_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_20_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_20_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_20_7 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_20_7  (
            .in0(N__14521),
            .in1(N__7852),
            .in2(N__8113),
            .in3(N__7862),
            .lcout(\this_vga_ramdac.N_1763_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_6_21_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_6_21_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_6_21_0 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_6_21_0  (
            .in0(N__8147),
            .in1(N__8103),
            .in2(N__8137),
            .in3(N__14533),
            .lcout(\this_vga_ramdac.N_1766_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22231),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_6_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_6_21_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_6_21_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_2_LC_6_21_2  (
            .in0(_gnd_net_),
            .in1(N__8783),
            .in2(_gnd_net_),
            .in3(N__8753),
            .lcout(\this_vga_signals.M_this_vga_signals_pixel_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22231),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_2_RNIRAOL5_LC_6_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_2_RNIRAOL5_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_2_RNIRAOL5_LC_6_21_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_2_RNIRAOL5_LC_6_21_4  (
            .in0(N__8120),
            .in1(N__8782),
            .in2(_gnd_net_),
            .in3(N__8752),
            .lcout(M_pcounter_q_ret_2_RNIRAOL5),
            .ltout(M_pcounter_q_ret_2_RNIRAOL5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_6_21_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_6_21_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_6_21_5 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_6_21_5  (
            .in0(N__14534),
            .in1(N__8065),
            .in2(N__8084),
            .in3(N__8081),
            .lcout(\this_vga_ramdac.N_1767_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22231),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_6_21_6 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_6_21_6 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_6_21_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_6_21_6  (
            .in0(_gnd_net_),
            .in1(N__8054),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22231),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHM2SG2_9_LC_7_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHM2SG2_9_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHM2SG2_9_LC_7_10_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIHM2SG2_9_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__9404),
            .in2(_gnd_net_),
            .in3(N__8189),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNICQMCG5_9_LC_7_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICQMCG5_9_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICQMCG5_9_LC_7_18_0 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNICQMCG5_9_LC_7_18_0  (
            .in0(N__8179),
            .in1(N__8201),
            .in2(N__9399),
            .in3(N__8159),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_7_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_7_18_1 .LUT_INIT=16'b0100010011011101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_7_18_1  (
            .in0(N__9820),
            .in1(N__9763),
            .in2(_gnd_net_),
            .in3(N__8316),
            .lcout(\this_vga_signals.mult1_un75_sum_c2_0 ),
            .ltout(\this_vga_signals.mult1_un75_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_18_2 .LUT_INIT=16'b0111000100010111;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_18_2  (
            .in0(N__11977),
            .in1(N__11936),
            .in2(N__8018),
            .in3(N__8015),
            .lcout(),
            .ltout(\this_vga_signals.if_N_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_18_3 .LUT_INIT=16'b0010011100011011;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_18_3  (
            .in0(N__9822),
            .in1(N__11938),
            .in2(N__8222),
            .in3(N__8178),
            .lcout(\this_vga_signals.mult1_un89_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_7_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_7_18_5 .LUT_INIT=16'b1110000101111000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_7_18_5  (
            .in0(N__8269),
            .in1(N__8317),
            .in2(N__8561),
            .in3(N__8219),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m5_i_LC_7_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m5_i_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m5_i_LC_7_18_6 .LUT_INIT=16'b0011001001001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_m5_i_LC_7_18_6  (
            .in0(N__8318),
            .in1(N__11935),
            .in2(N__9767),
            .in3(N__9821),
            .lcout(\this_vga_signals.N_2_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m1_0_LC_7_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m1_0_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m1_0_LC_7_19_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_haddress_if_m1_0_LC_7_19_0  (
            .in0(N__8643),
            .in1(N__9166),
            .in2(N__9761),
            .in3(N__9272),
            .lcout(),
            .ltout(\this_vga_signals.if_m1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_7_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_7_19_1 .LUT_INIT=16'b0011100000111110;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_7_19_1  (
            .in0(N__11931),
            .in1(N__9818),
            .in2(N__8213),
            .in3(N__8534),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_7_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_7_19_2 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_7_19_2  (
            .in0(N__8270),
            .in1(_gnd_net_),
            .in2(N__8210),
            .in3(N__8320),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_7_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_7_19_3 .LUT_INIT=16'b0000111101000100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_7_19_3  (
            .in0(N__8288),
            .in1(N__8294),
            .in2(N__8576),
            .in3(N__8207),
            .lcout(\this_vga_signals.mult1_un89_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_7_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_7_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_7_19_4  (
            .in0(N__8644),
            .in1(N__9165),
            .in2(_gnd_net_),
            .in3(N__9273),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_7_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_7_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_7_19_5  (
            .in0(N__8200),
            .in1(N__8177),
            .in2(_gnd_net_),
            .in3(N__8158),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIAPUMSC_9_LC_7_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIAPUMSC_9_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIAPUMSC_9_LC_7_19_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIAPUMSC_9_LC_7_19_6  (
            .in0(N__9400),
            .in1(N__8354),
            .in2(N__8348),
            .in3(N__8345),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNICOOCQ_1_LC_7_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNICOOCQ_1_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNICOOCQ_1_LC_7_19_7 .LUT_INIT=16'b1010010101001110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNICOOCQ_1_LC_7_19_7  (
            .in0(N__8321),
            .in1(N__9819),
            .in2(N__11939),
            .in3(N__9750),
            .lcout(\this_vga_signals.d_N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI97PTA_1_LC_7_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI97PTA_1_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI97PTA_1_LC_7_20_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI97PTA_1_LC_7_20_2  (
            .in0(N__11937),
            .in1(N__9827),
            .in2(_gnd_net_),
            .in3(N__8560),
            .lcout(\this_vga_signals.d_N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_c2_LC_7_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_c2_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_c2_LC_7_20_4 .LUT_INIT=16'b0100010011011101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_c2_LC_7_20_4  (
            .in0(N__10141),
            .in1(N__11060),
            .in2(_gnd_net_),
            .in3(N__9220),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_7_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_7_20_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_7_20_5  (
            .in0(N__9746),
            .in1(N__9167),
            .in2(N__8282),
            .in3(N__9274),
            .lcout(\this_vga_signals.mult1_un75_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_7_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_7_20_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_7_20_7  (
            .in0(N__9745),
            .in1(N__10142),
            .in2(_gnd_net_),
            .in3(N__9103),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIT1827_9_LC_9_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIT1827_9_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIT1827_9_LC_9_10_0 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIT1827_9_LC_9_10_0  (
            .in0(N__9403),
            .in1(N__9221),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIRETSA_9_LC_9_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIRETSA_9_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIRETSA_9_LC_9_10_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIRETSA_9_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__9402),
            .in2(_gnd_net_),
            .in3(N__9110),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_9_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_9_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11689),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22211),
            .ce(N__11590),
            .sr(N__11561));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_1_5_LC_9_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_1_5_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_1_5_LC_9_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_1_5_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__12531),
            .in2(_gnd_net_),
            .in3(N__12419),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_1_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_9_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_9_18_1 .LUT_INIT=16'b0000101100001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_26_LC_9_18_1  (
            .in0(N__10806),
            .in1(N__10680),
            .in2(N__8387),
            .in3(N__8612),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_9_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_9_18_4 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_LC_9_18_4  (
            .in0(N__8429),
            .in1(N__8498),
            .in2(N__8588),
            .in3(N__9617),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNISQ5DA02_9_LC_9_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNISQ5DA02_9_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNISQ5DA02_9_LC_9_18_5 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNISQ5DA02_9_LC_9_18_5  (
            .in0(N__9381),
            .in1(N__8450),
            .in2(N__8384),
            .in3(N__8456),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_2_i_m2_LC_9_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_2_i_m2_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_2_i_m2_LC_9_18_6 .LUT_INIT=16'b1000000101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_2_i_m2_LC_9_18_6  (
            .in0(N__12248),
            .in1(N__10807),
            .in2(N__12425),
            .in3(N__10669),
            .lcout(\this_vga_signals.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_9_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_9_19_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_9_19_0  (
            .in0(N__10010),
            .in1(N__9911),
            .in2(_gnd_net_),
            .in3(N__9026),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_ns_LC_9_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_ns_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_ns_LC_9_19_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_ns_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__8885),
            .in2(N__8363),
            .in3(N__8393),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0 ),
            .ltout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_LC_9_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_LC_9_19_2 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_LC_9_19_2  (
            .in0(N__13417),
            .in1(N__8444),
            .in2(N__8360),
            .in3(N__8480),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_9_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_9_19_3 .LUT_INIT=16'b1101010001001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_LC_9_19_3  (
            .in0(N__13302),
            .in1(N__13418),
            .in2(N__8357),
            .in3(N__8414),
            .lcout(),
            .ltout(\this_vga_signals.if_i1_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIOE1NOK_2_LC_9_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIOE1NOK_2_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIOE1NOK_2_LC_9_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIOE1NOK_2_LC_9_19_4  (
            .in0(N__8813),
            .in1(N__9569),
            .in2(N__8459),
            .in3(N__8428),
            .lcout(\this_vga_signals.g1_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_9_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_9_19_5 .LUT_INIT=16'b0011111000101100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_11_LC_9_19_5  (
            .in0(N__13303),
            .in1(N__10484),
            .in2(N__13427),
            .in3(N__8399),
            .lcout(\this_vga_signals.mult1_un75_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m1_3_LC_9_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m1_3_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m1_3_LC_9_19_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m1_3_LC_9_19_6  (
            .in0(N__12836),
            .in1(N__9027),
            .in2(N__12641),
            .in3(N__10012),
            .lcout(\this_vga_signals.if_m1_3 ),
            .ltout(\this_vga_signals.if_m1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_LC_9_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_LC_9_19_7 .LUT_INIT=16'b1111000001001011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_LC_9_19_7  (
            .in0(N__12832),
            .in1(N__8438),
            .in2(N__8432),
            .in3(N__8834),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_x1_LC_9_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_x1_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_x1_LC_9_20_0 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_x1_LC_9_20_0  (
            .in0(N__12775),
            .in1(N__9999),
            .in2(N__13426),
            .in3(N__9894),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_9_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_9_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_9_20_1  (
            .in0(N__10001),
            .in1(N__9020),
            .in2(N__9916),
            .in3(N__8875),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_9_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_9_20_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__8465),
            .in2(N__8417),
            .in3(N__8489),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_i ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_37_LC_9_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_37_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_37_LC_9_20_3 .LUT_INIT=16'b0111100000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_37_LC_9_20_3  (
            .in0(N__13419),
            .in1(N__8846),
            .in2(N__8408),
            .in3(N__8405),
            .lcout(\this_vga_signals.if_N_2_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x1_LC_9_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x1_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x1_LC_9_20_4 .LUT_INIT=16'b1101111011101101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x1_LC_9_20_4  (
            .in0(N__12590),
            .in1(N__12777),
            .in2(N__9030),
            .in3(N__9998),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_9_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_9_20_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_9_20_5  (
            .in0(N__10000),
            .in1(N__9019),
            .in2(N__9915),
            .in3(N__8874),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_9_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_9_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_9_20_6  (
            .in0(N__12776),
            .in1(N__9997),
            .in2(N__9031),
            .in3(N__9895),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_LC_9_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_LC_9_20_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_LC_9_20_7  (
            .in0(N__11521),
            .in1(_gnd_net_),
            .in2(N__11393),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.vaddress_6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_1_LC_9_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_1_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_1_LC_9_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_1_LC_9_21_0  (
            .in0(N__10008),
            .in1(N__9021),
            .in2(N__13247),
            .in3(N__9908),
            .lcout(),
            .ltout(\this_vga_signals.g0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_9_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_9_21_1 .LUT_INIT=16'b1000011111100001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_0_LC_9_21_1  (
            .in0(N__9909),
            .in1(N__12595),
            .in2(N__8483),
            .in3(N__12828),
            .lcout(\this_vga_signals.g0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_LC_9_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_LC_9_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_LC_9_21_2  (
            .in0(N__12827),
            .in1(N__8935),
            .in2(N__12640),
            .in3(N__9025),
            .lcout(),
            .ltout(\this_vga_signals.N_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_m3_LC_9_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_m3_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_m3_LC_9_21_3 .LUT_INIT=16'b0111000001111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_m3_LC_9_21_3  (
            .in0(N__13423),
            .in1(N__8479),
            .in2(N__8468),
            .in3(N__8828),
            .lcout(\this_vga_signals.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_9_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_9_21_4 .LUT_INIT=16'b0100010011011101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_9_21_4  (
            .in0(N__12591),
            .in1(N__12818),
            .in2(_gnd_net_),
            .in3(N__9907),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_12_x0_LC_9_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_12_x0_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_12_x0_LC_9_21_5 .LUT_INIT=16'b1110111111011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_12_x0_LC_9_21_5  (
            .in0(N__9906),
            .in1(N__12826),
            .in2(N__9032),
            .in3(N__10009),
            .lcout(\this_vga_signals.g0_12_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_9_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_9_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_2_LC_9_21_6  (
            .in0(N__9028),
            .in1(N__9602),
            .in2(N__12838),
            .in3(N__9910),
            .lcout(),
            .ltout(\this_vga_signals.g1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_9_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_9_21_7 .LUT_INIT=16'b1111000000101101;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_3_LC_9_21_7  (
            .in0(N__8879),
            .in1(N__12596),
            .in2(N__8600),
            .in3(N__8597),
            .lcout(\this_vga_signals.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI8OIBA_3_LC_9_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI8OIBA_3_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI8OIBA_3_LC_9_22_1 .LUT_INIT=16'b0110110011001001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI8OIBA_3_LC_9_22_1  (
            .in0(N__10134),
            .in1(N__9184),
            .in2(N__9752),
            .in3(N__9093),
            .lcout(\this_vga_signals.M_hcounter_q_RNI8OIBAZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_9_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_9_22_2 .LUT_INIT=16'b0010010011011011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_9_22_2  (
            .in0(N__9091),
            .in1(N__9735),
            .in2(N__10140),
            .in3(N__9185),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_9_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_9_22_3 .LUT_INIT=16'b1001001100110110;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_9_22_3  (
            .in0(N__10133),
            .in1(N__9183),
            .in2(N__9751),
            .in3(N__9092),
            .lcout(\this_vga_signals.if_N_8_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_9_1_LC_9_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_9_1_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_9_1_LC_9_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_9_1_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__12600),
            .in2(N__12837),
            .in3(N__8936),
            .lcout(),
            .ltout(\this_vga_signals.g0_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_12_ns_LC_9_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_12_ns_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_12_ns_LC_9_22_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_12_ns_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__8954),
            .in2(N__8522),
            .in3(N__8519),
            .lcout(),
            .ltout(\this_vga_signals.N_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_9_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_9_22_6 .LUT_INIT=16'b0110100110011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_8_LC_9_22_6  (
            .in0(N__9038),
            .in1(N__8513),
            .in2(N__8507),
            .in3(N__8504),
            .lcout(\this_vga_signals.d_N_3_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIF77A3_1_LC_9_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIF77A3_1_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIF77A3_1_LC_9_23_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNIF77A3_1_LC_9_23_1  (
            .in0(N__8731),
            .in1(N__14261),
            .in2(_gnd_net_),
            .in3(N__8678),
            .lcout(\this_vga_signals.N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_9_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_9_23_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_9_23_2 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_1_LC_9_23_2  (
            .in0(N__14116),
            .in1(N__8732),
            .in2(N__8717),
            .in3(N__8698),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22230),
            .ce(N__14262),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_9_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_9_23_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_0_LC_9_23_5  (
            .in0(N__8697),
            .in1(N__8765),
            .in2(_gnd_net_),
            .in3(N__14115),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22230),
            .ce(N__14262),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNI9C5I1_LC_9_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNI9C5I1_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNI9C5I1_LC_9_24_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_RNI9C5I1_LC_9_24_1  (
            .in0(N__14110),
            .in1(N__8693),
            .in2(_gnd_net_),
            .in3(N__8764),
            .lcout(),
            .ltout(\this_vga_signals.M_pcounter_q_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNII2VA2_0_LC_9_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNII2VA2_0_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNII2VA2_0_LC_9_24_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNII2VA2_0_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(N__8713),
            .in2(N__8786),
            .in3(N__14260),
            .lcout(\this_vga_signals.N_2_0 ),
            .ltout(\this_vga_signals.N_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_9_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_9_24_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_9_24_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8768),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_pcounter_q_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22232),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_LC_9_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_9_24_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_9_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8746),
            .lcout(\this_vga_signals.M_pcounter_q_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22232),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_RNI5GDH2_LC_9_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_RNI5GDH2_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_RNI5GDH2_LC_9_24_6 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_RNI5GDH2_LC_9_24_6  (
            .in0(N__8730),
            .in1(N__8712),
            .in2(N__8699),
            .in3(N__14109),
            .lcout(\this_vga_signals.M_pcounter_q_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHL0E5_9_LC_10_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHL0E5_9_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHL0E5_9_LC_10_16_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIHL0E5_9_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__9354),
            .in2(_gnd_net_),
            .in3(N__9239),
            .lcout(M_this_vga_signals_address_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIN0FTT_9_LC_10_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIN0FTT_9_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIN0FTT_9_LC_10_17_0 .LUT_INIT=16'b0100100010000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIN0FTT_9_LC_10_17_0  (
            .in0(N__9164),
            .in1(N__9353),
            .in2(N__8654),
            .in3(N__9275),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_6_LC_10_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_6_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_6_LC_10_17_4 .LUT_INIT=16'b1010010101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_6_LC_10_17_4  (
            .in0(N__12247),
            .in1(_gnd_net_),
            .in2(N__12421),
            .in3(N__12504),
            .lcout(\this_vga_signals.vaddress_1_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_1_6_LC_10_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_1_6_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_1_6_LC_10_17_5 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_1_6_LC_10_17_5  (
            .in0(N__12503),
            .in1(N__12409),
            .in2(_gnd_net_),
            .in3(N__12246),
            .lcout(\this_vga_signals.vaddress_4_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_10_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_10_17_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__10318),
            .in2(_gnd_net_),
            .in3(N__9505),
            .lcout(\this_vga_signals.vaddress_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_10_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_10_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11266),
            .lcout(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22204),
            .ce(N__11591),
            .sr(N__11562));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_10_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_10_18_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_10_18_1  (
            .in0(N__12953),
            .in1(N__10319),
            .in2(N__10238),
            .in3(N__10269),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_10_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_10_18_2 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_10_18_2  (
            .in0(N__9504),
            .in1(_gnd_net_),
            .in2(N__8801),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ),
            .ltout(\this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_10_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_10_18_3 .LUT_INIT=16'b1100011011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_10_18_3  (
            .in0(N__9291),
            .in1(N__10286),
            .in2(N__8798),
            .in3(N__9309),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_18_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11267),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22204),
            .ce(N__11591),
            .sr(N__11562));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_10_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_10_18_5 .LUT_INIT=16'b0000000000111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__9503),
            .in2(N__10321),
            .in3(N__8795),
            .lcout(),
            .ltout(\this_vga_signals.N_1_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNITEVS_6_LC_10_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNITEVS_6_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNITEVS_6_LC_10_18_6 .LUT_INIT=16'b1100111111101111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNITEVS_6_LC_10_18_6  (
            .in0(N__10234),
            .in1(N__9481),
            .in2(N__8789),
            .in3(N__12952),
            .lcout(\this_vga_signals.SUM_2_i_1_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11693),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22204),
            .ce(N__11591),
            .sr(N__11562));
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_10_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_10_19_0 .LUT_INIT=16'b0100011010010001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_35_LC_10_19_0  (
            .in0(N__10643),
            .in1(N__8920),
            .in2(N__10791),
            .in3(N__11729),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_1_1_LC_10_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_1_1_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_1_1_LC_10_19_1 .LUT_INIT=16'b0000101010110001;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_1_1_LC_10_19_1  (
            .in0(N__11379),
            .in1(N__10400),
            .in2(N__12249),
            .in3(N__10642),
            .lcout(\this_vga_signals.g1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_10_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_10_19_3 .LUT_INIT=16'b0010010010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_14_LC_10_19_3  (
            .in0(N__10187),
            .in1(N__10756),
            .in2(N__10202),
            .in3(N__10641),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_10_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_10_19_4 .LUT_INIT=16'b0101100000100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_10_19_4  (
            .in0(N__10639),
            .in1(N__9558),
            .in2(N__10790),
            .in3(N__11424),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i ),
            .ltout(\this_vga_signals.mult1_un54_sum_axb2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_10_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_10_19_5 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_23_LC_10_19_5  (
            .in0(N__12648),
            .in1(N__8822),
            .in2(N__8816),
            .in3(N__10452),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_10_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_10_19_6 .LUT_INIT=16'b0110010000011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m2_1_LC_10_19_6  (
            .in0(N__10638),
            .in1(N__9557),
            .in2(N__10789),
            .in3(N__11423),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_10_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_10_19_7 .LUT_INIT=16'b0100010101010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_10_19_7  (
            .in0(N__11422),
            .in1(N__10755),
            .in2(N__9560),
            .in3(N__10640),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_10_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_10_20_0 .LUT_INIT=16'b1010101001001101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_10_20_0  (
            .in0(N__11391),
            .in1(N__12769),
            .in2(N__10454),
            .in3(N__10522),
            .lcout(\this_vga_signals.mult1_un61_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_395_LC_10_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_395_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_395_LC_10_20_1 .LUT_INIT=16'b1011010010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_395_LC_10_20_1  (
            .in0(N__8807),
            .in1(N__11389),
            .in2(N__9601),
            .in3(N__8873),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_395 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axb1_395_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x0_LC_10_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x0_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x0_LC_10_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x0_LC_10_20_2  (
            .in0(N__12618),
            .in1(N__12773),
            .in2(N__8888),
            .in3(N__9005),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_10_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_10_20_3 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_10_20_3  (
            .in0(N__9592),
            .in1(N__11390),
            .in2(N__10453),
            .in3(N__8872),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_2_LC_10_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_2_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_2_LC_10_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_2_LC_10_20_4  (
            .in0(N__9596),
            .in1(N__12774),
            .in2(N__8852),
            .in3(N__9006),
            .lcout(),
            .ltout(\this_vga_signals.g0_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_10_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_10_20_5 .LUT_INIT=16'b0001100000100100;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_5_LC_10_20_5  (
            .in0(N__9007),
            .in1(N__9512),
            .in2(N__8849),
            .in3(N__8903),
            .lcout(\this_vga_signals.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_ns_LC_10_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_ns_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_ns_LC_10_20_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_ns_LC_10_20_6  (
            .in0(N__8840),
            .in1(N__9947),
            .in2(_gnd_net_),
            .in3(N__9008),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_10_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_10_20_7 .LUT_INIT=16'b1011101001010001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_17_LC_10_20_7  (
            .in0(N__10523),
            .in1(N__10449),
            .in2(N__12816),
            .in3(N__12617),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_10_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_10_21_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_10_21_0  (
            .in0(N__12619),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12400),
            .lcout(\this_vga_signals.vaddress_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_10_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_10_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_29_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__10006),
            .in2(N__9029),
            .in3(N__9902),
            .lcout(\this_vga_signals.N_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_10_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_10_21_2 .LUT_INIT=16'b1010010101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_10_21_2  (
            .in0(N__12253),
            .in1(_gnd_net_),
            .in2(N__12646),
            .in3(N__12401),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_10_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_10_21_3 .LUT_INIT=16'b0001100011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_9_LC_10_21_3  (
            .in0(N__10810),
            .in1(N__9047),
            .in2(N__9041),
            .in3(N__9332),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_12_x1_LC_10_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_12_x1_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_12_x1_LC_10_21_4 .LUT_INIT=16'b1111111111011110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_12_x1_LC_10_21_4  (
            .in0(N__10007),
            .in1(N__12819),
            .in2(N__9917),
            .in3(N__9012),
            .lcout(\this_vga_signals.g0_12_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_2_1_0_LC_10_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_2_1_0_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_2_1_0_LC_10_21_6 .LUT_INIT=16'b0011010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_2_1_0_LC_10_21_6  (
            .in0(N__11387),
            .in1(N__10809),
            .in2(N__12257),
            .in3(N__10671),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_2_LC_10_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_2_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_2_LC_10_21_7 .LUT_INIT=16'b0001101111100100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_2_LC_10_21_7  (
            .in0(N__12399),
            .in1(N__11388),
            .in2(N__8948),
            .in3(N__8945),
            .lcout(\this_vga_signals.g0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_10_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_10_22_0 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_10_22_0  (
            .in0(N__11122),
            .in1(N__9235),
            .in2(N__11057),
            .in3(N__9121),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_2_9_LC_10_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_2_9_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_2_9_LC_10_22_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_2_9_LC_10_22_1  (
            .in0(N__10909),
            .in1(N__11175),
            .in2(N__11132),
            .in3(N__10974),
            .lcout(\this_vga_signals.N_236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_10_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_10_22_4 .LUT_INIT=16'b0010010011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_LC_10_22_4  (
            .in0(N__11727),
            .in1(N__10808),
            .in2(N__8924),
            .in3(N__10670),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axb2_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_10_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_10_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_0_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(N__12645),
            .in2(N__8906),
            .in3(N__12817),
            .lcout(\this_vga_signals.g0_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_0_LC_10_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_0_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_0_LC_10_22_6 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_0_LC_10_22_6  (
            .in0(N__11123),
            .in1(N__8894),
            .in2(N__11058),
            .in3(N__9422),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_2_LC_10_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_2_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_2_LC_10_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_2_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(N__9207),
            .in2(N__9278),
            .in3(N__9087),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_10_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_10_23_0 .LUT_INIT=16'b0001111010000111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_10_23_0  (
            .in0(N__10972),
            .in1(N__11173),
            .in2(N__11128),
            .in3(N__10907),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_10_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_10_23_1 .LUT_INIT=16'b1011010101010111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_10_23_1  (
            .in0(N__10906),
            .in1(N__11107),
            .in2(N__11186),
            .in3(N__10971),
            .lcout(\this_vga_signals.N_3_2_1 ),
            .ltout(\this_vga_signals.N_3_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_LC_10_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_LC_10_23_2 .LUT_INIT=16'b0101100010000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_LC_10_23_2  (
            .in0(N__11027),
            .in1(N__10109),
            .in2(N__9224),
            .in3(N__11121),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_10_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_10_23_3 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_10_23_3  (
            .in0(N__9206),
            .in1(_gnd_net_),
            .in2(N__10129),
            .in3(N__11028),
            .lcout(\this_vga_signals.mult1_un68_sum_axb2_1 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axb2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_23_4 .LUT_INIT=16'b0100111100001101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_23_4  (
            .in0(N__9703),
            .in1(N__10113),
            .in2(N__9170),
            .in3(N__9086),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_10_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_10_23_5 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_10_23_5  (
            .in0(N__9053),
            .in1(N__9131),
            .in2(N__9125),
            .in3(N__9410),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_10_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_10_23_6 .LUT_INIT=16'b0011111000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_10_23_6  (
            .in0(N__11106),
            .in1(N__11169),
            .in2(N__10983),
            .in3(N__10905),
            .lcout(\this_vga_signals.SUM_3_i_0_0_3 ),
            .ltout(\this_vga_signals.SUM_3_i_0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_0_LC_10_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_0_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_0_LC_10_23_7 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_0_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(N__11111),
            .in2(N__9056),
            .in3(N__11026),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_24_1 .LUT_INIT=16'b1100110111001101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_24_1  (
            .in0(N__11191),
            .in1(N__10982),
            .in2(N__10928),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_hvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_10_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_10_24_7 .LUT_INIT=16'b0000001110100011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_10_24_7  (
            .in0(N__11129),
            .in1(N__10123),
            .in2(N__11059),
            .in3(N__9421),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIE00C4_9_LC_11_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIE00C4_9_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIE00C4_9_LC_11_17_0 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIE00C4_9_LC_11_17_0  (
            .in0(N__10988),
            .in1(N__10927),
            .in2(N__10047),
            .in3(N__11187),
            .lcout(M_this_vga_ramdac_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_7_1_LC_11_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_1_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_1_LC_11_17_3 .LUT_INIT=16'b1010101010010101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_1_LC_11_17_3  (
            .in0(N__12023),
            .in1(N__12413),
            .in2(N__12609),
            .in3(N__12254),
            .lcout(),
            .ltout(\this_vga_signals.g0_7_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_11_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_11_17_4 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_13_LC_11_17_4  (
            .in0(N__9320),
            .in1(N__9293),
            .in2(N__9335),
            .in3(N__9311),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_11_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_11_17_6 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_LC_11_17_6  (
            .in0(N__9319),
            .in1(N__9292),
            .in2(N__10331),
            .in3(N__9310),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_axb1_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_11_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_11_17_7 .LUT_INIT=16'b0010100101001001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_25_LC_11_17_7  (
            .in0(N__11656),
            .in1(N__10349),
            .in2(N__9296),
            .in3(N__10779),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIVA761_6_LC_11_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIVA761_6_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIVA761_6_LC_11_18_0 .LUT_INIT=16'b1010011110101111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIVA761_6_LC_11_18_0  (
            .in0(N__10230),
            .in1(N__10273),
            .in2(N__12964),
            .in3(N__9480),
            .lcout(\this_vga_signals.SUM_2_i_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11756),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22202),
            .ce(N__11593),
            .sr(N__11560));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_11_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_11_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11237),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22202),
            .ce(N__11593),
            .sr(N__11560));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_11_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_11_18_3 .LUT_INIT=16'b0011111100101010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_11_18_3  (
            .in0(N__10388),
            .in1(N__12957),
            .in2(N__10277),
            .in3(N__10231),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_18_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_18_4  (
            .in0(N__10320),
            .in1(N__9506),
            .in2(N__9485),
            .in3(N__9464),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_11_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_11_18_5 .LUT_INIT=16'b0000111000010111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_11_18_5  (
            .in0(N__12958),
            .in1(N__10270),
            .in2(N__9455),
            .in3(N__10232),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_11_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_11_18_6 .LUT_INIT=16'b1011000011010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_11_18_6  (
            .in0(N__9452),
            .in1(N__11769),
            .in2(N__9446),
            .in3(N__10389),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_11_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_11_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11626),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22202),
            .ce(N__11593),
            .sr(N__11560));
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_11_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_11_19_0 .LUT_INIT=16'b0100001010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_24_LC_11_19_0  (
            .in0(N__10765),
            .in1(N__10342),
            .in2(N__11657),
            .in3(N__10646),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_11_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_11_19_1 .LUT_INIT=16'b0110000101001001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_34_LC_11_19_1  (
            .in0(N__10647),
            .in1(N__10817),
            .in2(N__10826),
            .in3(N__10766),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_LC_11_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_LC_11_19_2 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_LC_11_19_2  (
            .in0(N__11508),
            .in1(N__11453),
            .in2(_gnd_net_),
            .in3(N__10391),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(\this_vga_signals.vaddress_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_11_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_11_19_3 .LUT_INIT=16'b0100010101010100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_LC_11_19_3  (
            .in0(N__10837),
            .in1(N__11426),
            .in2(N__9605),
            .in3(N__10760),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_11_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_11_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_19_LC_11_19_4  (
            .in0(N__10764),
            .in1(N__10392),
            .in2(N__11520),
            .in3(N__10645),
            .lcout(\this_vga_signals.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIPQ6L81_2_LC_11_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIPQ6L81_2_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIPQ6L81_2_LC_11_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIPQ6L81_2_LC_11_19_5  (
            .in0(N__10474),
            .in1(N__10568),
            .in2(N__12881),
            .in3(N__9600),
            .lcout(\this_vga_signals.g1_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_N_2L1_LC_11_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_N_2L1_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_N_2L1_LC_11_19_6 .LUT_INIT=16'b0100001010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_N_2L1_LC_11_19_6  (
            .in0(N__9559),
            .in1(N__11425),
            .in2(N__10792),
            .in3(N__10644),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_11_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_11_19_7 .LUT_INIT=16'b0000111000000110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_32_LC_11_19_7  (
            .in0(N__10648),
            .in1(N__9539),
            .in2(N__9530),
            .in3(N__10767),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_2_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_11_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_11_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__12610),
            .in2(_gnd_net_),
            .in3(N__12361),
            .lcout(\this_vga_signals.vaddress_5_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_LC_11_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_LC_11_20_1 .LUT_INIT=16'b1111010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_LC_11_20_1  (
            .in0(N__10673),
            .in1(_gnd_net_),
            .in2(N__10811),
            .in3(N__10561),
            .lcout(\this_vga_signals.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_11_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_11_20_2 .LUT_INIT=16'b1101110110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_0_LC_11_20_2  (
            .in0(N__11728),
            .in1(N__10801),
            .in2(_gnd_net_),
            .in3(N__10672),
            .lcout(),
            .ltout(\this_vga_signals.g2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_11_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_11_20_3 .LUT_INIT=16'b0100110001101111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_4_LC_11_20_3  (
            .in0(N__12362),
            .in1(N__12623),
            .in2(N__9521),
            .in3(N__9518),
            .lcout(\this_vga_signals.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_11_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_11_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_15_LC_11_20_4  (
            .in0(N__9941),
            .in1(N__10011),
            .in2(_gnd_net_),
            .in3(N__9912),
            .lcout(\this_vga_signals.N_5_i_5 ),
            .ltout(\this_vga_signals.N_5_i_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_0_LC_11_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_0_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_0_LC_11_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x2_0_LC_11_20_5  (
            .in0(N__13401),
            .in1(N__9668),
            .in2(N__9659),
            .in3(N__9833),
            .lcout(\this_vga_signals.g0_i_x2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_11_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_11_20_6 .LUT_INIT=16'b0000010001010100;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_1_LC_11_20_6  (
            .in0(N__9656),
            .in1(N__11392),
            .in2(N__11525),
            .in3(N__9650),
            .lcout(\this_vga_signals.g1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_31_1_LC_11_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_1_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_1_LC_11_20_7 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_1_LC_11_20_7  (
            .in0(N__12793),
            .in1(N__9644),
            .in2(N__12644),
            .in3(N__10524),
            .lcout(\this_vga_signals.g0_31_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_x0_LC_11_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_x0_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_x0_LC_11_21_0 .LUT_INIT=16'b0111110111010111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_x0_LC_11_21_0  (
            .in0(N__13403),
            .in1(N__12809),
            .in2(N__9914),
            .in3(N__9937),
            .lcout(),
            .ltout(\this_vga_signals.g0_2_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_ns_LC_11_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_ns_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_ns_LC_11_21_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_ns_LC_11_21_1  (
            .in0(N__10005),
            .in1(_gnd_net_),
            .in2(N__9638),
            .in3(N__9923),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_11_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_11_21_2 .LUT_INIT=16'b1010000011010101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_LC_11_21_2  (
            .in0(N__10499),
            .in1(N__12810),
            .in2(N__9635),
            .in3(N__9632),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_11_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_11_21_3 .LUT_INIT=16'b0000011001100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_0_LC_11_21_3  (
            .in0(N__13301),
            .in1(N__12866),
            .in2(N__9626),
            .in3(N__9623),
            .lcout(\this_vga_signals.if_i4_mux_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_11_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_11_21_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_11_21_4  (
            .in0(N__12122),
            .in1(N__12625),
            .in2(N__12408),
            .in3(N__12965),
            .lcout(\this_vga_signals.vsync_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_x0_LC_11_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_x0_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_x0_LC_11_21_5 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_1_x0_LC_11_21_5  (
            .in0(N__12806),
            .in1(N__13404),
            .in2(N__10013),
            .in3(N__9887),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_1_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_x1_LC_11_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_x1_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_x1_LC_11_21_6 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_x1_LC_11_21_6  (
            .in0(N__13402),
            .in1(N__12808),
            .in2(N__9913),
            .in3(N__9936),
            .lcout(\this_vga_signals.g0_2_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_11_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_11_21_7 .LUT_INIT=16'b0010001010111011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_20_LC_11_21_7  (
            .in0(N__12807),
            .in1(N__12624),
            .in2(_gnd_net_),
            .in3(N__9886),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_22_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__11930),
            .in2(N__11978),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_11_22_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_11_22_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_11_22_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_11_22_1  (
            .in0(N__14267),
            .in1(N__9796),
            .in2(_gnd_net_),
            .in3(N__9770),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__22221),
            .ce(),
            .sr(N__15056));
    defparam \this_vga_signals.M_hcounter_q_3_LC_11_22_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_11_22_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_11_22_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_11_22_2  (
            .in0(N__14264),
            .in1(N__9721),
            .in2(_gnd_net_),
            .in3(N__9680),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__22221),
            .ce(),
            .sr(N__15056));
    defparam \this_vga_signals.M_hcounter_q_4_LC_11_22_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_11_22_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_11_22_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_11_22_3  (
            .in0(N__14268),
            .in1(N__10122),
            .in2(_gnd_net_),
            .in3(N__9677),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__22221),
            .ce(),
            .sr(N__15056));
    defparam \this_vga_signals.M_hcounter_q_5_LC_11_22_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_11_22_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_11_22_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_11_22_4  (
            .in0(N__14265),
            .in1(N__11048),
            .in2(_gnd_net_),
            .in3(N__9674),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__22221),
            .ce(),
            .sr(N__15056));
    defparam \this_vga_signals.M_hcounter_q_6_LC_11_22_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_11_22_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_11_22_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_11_22_5  (
            .in0(N__14269),
            .in1(N__11127),
            .in2(_gnd_net_),
            .in3(N__9671),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__22221),
            .ce(),
            .sr(N__15056));
    defparam \this_vga_signals.M_hcounter_q_7_LC_11_22_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_11_22_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_11_22_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_11_22_6  (
            .in0(N__14266),
            .in1(N__11182),
            .in2(_gnd_net_),
            .in3(N__10175),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__22221),
            .ce(),
            .sr(N__15056));
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_22_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_22_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_22_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_11_22_7  (
            .in0(N__14270),
            .in1(N__10919),
            .in2(_gnd_net_),
            .in3(N__10172),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__22221),
            .ce(),
            .sr(N__15056));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_11_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_11_23_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__10981),
            .in2(_gnd_net_),
            .in3(N__10169),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22223),
            .ce(N__10865),
            .sr(N__15048));
    defparam \this_vga_signals.M_hcounter_q_RNIC1AR_5_LC_11_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIC1AR_5_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIC1AR_5_LC_11_24_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIC1AR_5_LC_11_24_2  (
            .in0(N__11130),
            .in1(N__10127),
            .in2(_gnd_net_),
            .in3(N__11055),
            .lcout(),
            .ltout(\this_vga_signals.un4_hsynclt8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIMBHF2_9_LC_11_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIMBHF2_9_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIMBHF2_9_LC_11_24_3 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIMBHF2_9_LC_11_24_3  (
            .in0(N__10987),
            .in1(N__10067),
            .in2(N__10166),
            .in3(N__10923),
            .lcout(this_vga_signals_hsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIIED41_7_LC_11_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIIED41_7_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIIED41_7_LC_11_24_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIIED41_7_LC_11_24_5  (
            .in0(N__10128),
            .in1(N__11056),
            .in2(N__11192),
            .in3(N__11131),
            .lcout(\this_vga_signals.un3_hsynclt8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_8_LC_12_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_8_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_8_LC_12_17_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIROQM_8_LC_12_17_0  (
            .in0(N__12019),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12118),
            .lcout(),
            .ltout(\this_vga_signals.un6_vvisibilitylto8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_12_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_12_17_1 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_12_17_1  (
            .in0(N__12219),
            .in1(N__12545),
            .in2(N__10061),
            .in3(N__12414),
            .lcout(\this_vga_signals.un6_vvisibilitylt9_0 ),
            .ltout(\this_vga_signals.un6_vvisibilitylt9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_9_LC_12_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_9_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_9_LC_12_17_2 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_9_LC_12_17_2  (
            .in0(N__11806),
            .in1(N__11776),
            .in2(N__10058),
            .in3(N__12949),
            .lcout(\this_vga_signals.vvisibility ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_12_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_12_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_12_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11260),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22189),
            .ce(N__11592),
            .sr(N__11556));
    defparam \this_vga_signals.un5_vaddress_g0_7_0_LC_12_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_0_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_0_LC_12_17_4 .LUT_INIT=16'b1110000111000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_0_LC_12_17_4  (
            .in0(N__11519),
            .in1(N__12218),
            .in2(N__12038),
            .in3(N__11380),
            .lcout(\this_vga_signals.g0_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_12_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_12_18_0 .LUT_INIT=16'b1110110000010011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_12_18_0  (
            .in0(N__11448),
            .in1(N__10386),
            .in2(N__10322),
            .in3(N__10271),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_12_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_12_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11681),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22194),
            .ce(N__11594),
            .sr(N__11558));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_12_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_12_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_12_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11748),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22194),
            .ce(N__11594),
            .sr(N__11558));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_12_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_12_18_3 .LUT_INIT=16'b0110110110110111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_12_18_3  (
            .in0(N__10272),
            .in1(N__10233),
            .in2(N__12962),
            .in3(N__10390),
            .lcout(),
            .ltout(\this_vga_signals.if_m8_0_a3_1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_18_4 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_18_4  (
            .in0(N__11449),
            .in1(_gnd_net_),
            .in2(N__10241),
            .in3(N__11489),
            .lcout(\this_vga_signals.if_N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_12_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_12_18_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_12_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11232),
            .lcout(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22194),
            .ce(N__11594),
            .sr(N__11558));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_0_LC_12_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_0_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_0_LC_12_18_6 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIBS0H_0_LC_12_18_6  (
            .in0(N__11451),
            .in1(N__10387),
            .in2(_gnd_net_),
            .in3(N__11491),
            .lcout(\this_vga_signals.vaddress_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_0_LC_12_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_0_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_0_LC_12_18_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_0_LC_12_18_7  (
            .in0(N__11490),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11450),
            .lcout(\this_vga_signals.vaddress_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_22_1_LC_12_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_22_1_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_22_1_LC_12_19_0 .LUT_INIT=16'b0011001111000110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_22_1_LC_12_19_0  (
            .in0(N__10415),
            .in1(N__12812),
            .in2(N__12643),
            .in3(N__10493),
            .lcout(),
            .ltout(\this_vga_signals.g0_22_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_12_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_12_19_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_22_LC_12_19_1  (
            .in0(N__10460),
            .in1(N__10406),
            .in2(N__10487),
            .in3(N__10475),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_12_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_12_19_2 .LUT_INIT=16'b1111000000101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_LC_12_19_2  (
            .in0(N__12811),
            .in1(N__10451),
            .in2(N__12642),
            .in3(N__10528),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_0_LC_12_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_0_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_0_LC_12_19_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_0_LC_12_19_3  (
            .in0(N__11340),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12386),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_5_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_12_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_12_19_4 .LUT_INIT=16'b0101001010000101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_38_LC_12_19_4  (
            .in0(N__10681),
            .in1(N__11288),
            .in2(N__10463),
            .in3(N__10783),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axb2_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_12_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_12_19_5 .LUT_INIT=16'b1010100010101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_36_LC_12_19_5  (
            .in0(N__10450),
            .in1(N__12602),
            .in2(N__10418),
            .in3(N__10414),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIC07L_LC_12_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIC07L_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIC07L_LC_12_19_6 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIC07L_LC_12_19_6  (
            .in0(N__11512),
            .in1(N__11338),
            .in2(_gnd_net_),
            .in3(N__10393),
            .lcout(\this_vga_signals.vaddress_2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_12_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_12_19_7 .LUT_INIT=16'b0111111011100111;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_1_LC_12_19_7  (
            .in0(N__11339),
            .in1(N__12385),
            .in2(N__12255),
            .in3(N__10773),
            .lcout(\this_vga_signals.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_12_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_12_20_0 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_LC_12_20_0  (
            .in0(N__12728),
            .in1(N__10847),
            .in2(N__12649),
            .in3(N__10841),
            .lcout(\this_vga_signals.g1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_LC_12_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_LC_12_20_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_LC_12_20_1  (
            .in0(N__12338),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11359),
            .lcout(\this_vga_signals.vaddress_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_0_LC_12_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_0_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_0_LC_12_20_2 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_0_LC_12_20_2  (
            .in0(N__11358),
            .in1(N__12339),
            .in2(_gnd_net_),
            .in3(N__12209),
            .lcout(\this_vga_signals.vaddress_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_1_LC_12_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_1_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_1_LC_12_20_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIK3QQ_1_LC_12_20_3  (
            .in0(N__12341),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11357),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_12_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_12_20_4 .LUT_INIT=16'b0100001010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_LC_12_20_4  (
            .in0(N__10562),
            .in1(N__10805),
            .in2(N__10685),
            .in3(N__10682),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_LC_12_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_LC_12_20_5 .LUT_INIT=16'b0100011011001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_LC_12_20_5  (
            .in0(N__12342),
            .in1(N__12635),
            .in2(N__10577),
            .in3(N__10574),
            .lcout(\this_vga_signals.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_LC_12_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_LC_12_20_6 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_LC_12_20_6  (
            .in0(N__11356),
            .in1(N__12340),
            .in2(_gnd_net_),
            .in3(N__12210),
            .lcout(\this_vga_signals.vaddress_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_12_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_12_21_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_12_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11630),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22212),
            .ce(N__11597),
            .sr(N__11563));
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_12_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_12_21_7 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_LC_12_21_7  (
            .in0(N__10550),
            .in1(N__10544),
            .in2(N__10538),
            .in3(N__10529),
            .lcout(\this_vga_signals.N_5_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_22_0 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_22_0  (
            .in0(N__10859),
            .in1(N__11216),
            .in2(N__12256),
            .in3(N__10871),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_12_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_12_22_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_12_22_3  (
            .in0(_gnd_net_),
            .in1(N__11174),
            .in2(_gnd_net_),
            .in3(N__11120),
            .lcout(),
            .ltout(\this_vga_signals.M_hcounter_d7lto7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI704B1_9_LC_12_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI704B1_9_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI704B1_9_LC_12_22_4 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI704B1_9_LC_12_22_4  (
            .in0(N__11047),
            .in1(N__10973),
            .in2(N__10931),
            .in3(N__10908),
            .lcout(\this_vga_signals.M_hcounter_d7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_22_7 .LUT_INIT=16'b0000010100010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_22_7  (
            .in0(N__12650),
            .in1(N__13424),
            .in2(N__12839),
            .in3(N__13304),
            .lcout(\this_vga_signals.un2_vsynclt8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_12_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_12_23_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__14239),
            .in2(_gnd_net_),
            .in3(N__15047),
            .lcout(\this_vga_signals.N_340_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_23_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_23_7  (
            .in0(_gnd_net_),
            .in1(N__13425),
            .in2(_gnd_net_),
            .in3(N__12047),
            .lcout(\this_vga_signals.vsync_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_13_17_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_13_17_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_13_17_0  (
            .in0(N__14256),
            .in1(N__12862),
            .in2(N__14120),
            .in3(N__14114),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__22183),
            .ce(),
            .sr(N__11555));
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_17_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_17_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_13_17_1  (
            .in0(N__14258),
            .in1(N__13285),
            .in2(_gnd_net_),
            .in3(N__10853),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__22183),
            .ce(),
            .sr(N__11555));
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_17_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_17_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_13_17_2  (
            .in0(N__14257),
            .in1(N__13363),
            .in2(_gnd_net_),
            .in3(N__10850),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__22183),
            .ce(),
            .sr(N__11555));
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_17_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_17_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_13_17_3  (
            .in0(N__14259),
            .in1(N__12710),
            .in2(_gnd_net_),
            .in3(N__11279),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__22183),
            .ce(),
            .sr(N__11555));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_17_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__12639),
            .in2(_gnd_net_),
            .in3(N__11276),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_17_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__12418),
            .in2(_gnd_net_),
            .in3(N__11273),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_17_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__12242),
            .in2(_gnd_net_),
            .in3(N__11270),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_17_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__12046),
            .in2(_gnd_net_),
            .in3(N__11246),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_18_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__12112),
            .in2(_gnd_net_),
            .in3(N__11243),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_13_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_13_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_13_18_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__12951),
            .in2(_gnd_net_),
            .in3(N__11240),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22190),
            .ce(N__11595),
            .sr(N__11557));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_8_LC_13_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_8_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_8_LC_13_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_8_LC_13_19_0  (
            .in0(N__12039),
            .in1(N__12948),
            .in2(N__12117),
            .in3(N__12184),
            .lcout(\this_vga_signals.vaddress_ac0_9_0_a0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_13_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_13_19_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_13_19_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__11233),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22195),
            .ce(N__11596),
            .sr(N__11559));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_13_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_13_19_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_13_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11752),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22195),
            .ce(N__11596),
            .sr(N__11559));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_LC_13_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_LC_13_19_3 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIE35R_LC_13_19_3  (
            .in0(N__12183),
            .in1(N__11342),
            .in2(_gnd_net_),
            .in3(N__11488),
            .lcout(\this_vga_signals.vaddress_5_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_LC_13_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_LC_13_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11688),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22195),
            .ce(N__11596),
            .sr(N__11559));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_0_LC_13_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_0_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_0_LC_13_19_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIIONF_0_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__11341),
            .in2(_gnd_net_),
            .in3(N__11487),
            .lcout(\this_vga_signals.vaddress_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_13_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_13_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11614),
            .lcout(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22195),
            .ce(N__11596),
            .sr(N__11559));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_LC_13_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_LC_13_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIHKHB_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__11486),
            .in2(_gnd_net_),
            .in3(N__11452),
            .lcout(\this_vga_signals.vaddress_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_1_LC_13_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_1_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_1_LC_13_20_0 .LUT_INIT=16'b1010010101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep2_esr_RNIGE761_1_LC_13_20_0  (
            .in0(N__12186),
            .in1(_gnd_net_),
            .in2(N__12379),
            .in3(N__11360),
            .lcout(\this_vga_signals.vaddress_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_0_8_LC_13_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_0_8_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_0_8_LC_13_20_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_0_8_LC_13_20_3  (
            .in0(N__12048),
            .in1(N__12334),
            .in2(N__12116),
            .in3(N__12185),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_d7lto8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_13_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_13_20_4 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_13_20_4  (
            .in0(N__12278),
            .in1(N__12601),
            .in2(N__11282),
            .in3(N__12963),
            .lcout(\this_vga_signals.M_vcounter_d8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_13_20_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_13_20_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_13_20_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_13_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_13_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_13_21_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_13_21_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_13_21_3  (
            .in0(N__11964),
            .in1(N__11900),
            .in2(_gnd_net_),
            .in3(N__14231),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22205),
            .ce(),
            .sr(N__15037));
    defparam \this_delay_clk.M_pipe_q_4_LC_13_22_1 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_13_22_1 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_13_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11861),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22213),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_address_delay.out_LC_13_22_2 .C_ON=1'b0;
    defparam \this_start_address_delay.out_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \this_start_address_delay.out_LC_13_22_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \this_start_address_delay.out_LC_13_22_2  (
            .in0(N__11854),
            .in1(_gnd_net_),
            .in2(N__11819),
            .in3(N__11841),
            .lcout(M_this_start_address_delay_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_13_22_4 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_13_22_4 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_13_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11876),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22213),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_13_22_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_13_22_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBJQQ_LC_13_22_5  (
            .in0(N__11843),
            .in1(N__11815),
            .in2(_gnd_net_),
            .in3(N__11853),
            .lcout(M_this_start_data_delay_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_13_22_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_13_22_6 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_13_22_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_13_22_6  (
            .in0(N__11855),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11842),
            .lcout(this_start_data_delay_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22213),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIQ80L_2_LC_13_23_4.C_ON=1'b0;
    defparam M_this_state_q_RNIQ80L_2_LC_13_23_4.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIQ80L_2_LC_13_23_4.LUT_INIT=16'b0000000000010001;
    LogicCell40 M_this_state_q_RNIQ80L_2_LC_13_23_4 (
            .in0(N__20922),
            .in1(N__16213),
            .in2(_gnd_net_),
            .in3(N__20388),
            .lcout(port_dmab_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBILS3_6_LC_14_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBILS3_6_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBILS3_6_LC_14_17_2 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIBILS3_6_LC_14_17_2  (
            .in0(N__11807),
            .in1(N__11789),
            .in2(N__13208),
            .in3(N__11780),
            .lcout(M_this_ppu_vga_is_drawing_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_14_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_14_18_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_14_18_1  (
            .in0(N__14336),
            .in1(N__14366),
            .in2(_gnd_net_),
            .in3(N__12950),
            .lcout(\this_vga_signals.line_clk_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIV19S_2_LC_14_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIV19S_2_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIV19S_2_LC_14_18_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIV19S_2_LC_14_18_4  (
            .in0(N__12681),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13339),
            .lcout(\this_vga_signals.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_18_7 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_18_7  (
            .in0(N__13272),
            .in1(N__12852),
            .in2(N__13364),
            .in3(N__12680),
            .lcout(\this_vga_signals.M_vcounter_d7lt8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_14_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_14_19_3 .LUT_INIT=16'b0000000000110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_14_19_3  (
            .in0(N__12647),
            .in1(N__12420),
            .in2(N__12277),
            .in3(N__12211),
            .lcout(\this_vga_signals.un4_lvisibility_1 ),
            .ltout(\this_vga_signals.un4_lvisibility_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICHRV3_8_LC_14_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICHRV3_8_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICHRV3_8_LC_14_19_4 .LUT_INIT=16'b1010001010001010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICHRV3_8_LC_14_19_4  (
            .in0(N__12067),
            .in1(N__12110),
            .in2(N__12125),
            .in3(N__12049),
            .lcout(M_this_vga_signals_line_clk_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_LC_14_19_7 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_LC_14_19_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.line_clk.M_last_q_LC_14_19_7 .LUT_INIT=16'b1100010010001100;
    LogicCell40 \this_ppu.line_clk.M_last_q_LC_14_19_7  (
            .in0(N__12111),
            .in1(N__12068),
            .in2(N__12059),
            .in3(N__12050),
            .lcout(\this_ppu.line_clk.M_last_qZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22191),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_0_LC_14_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_14_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_14_20_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__11963),
            .in2(_gnd_net_),
            .in3(N__14235),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22196),
            .ce(),
            .sr(N__15055));
    defparam M_this_sprites_address_q_RNO_0_5_LC_14_21_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_5_LC_14_21_0.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_5_LC_14_21_0.LUT_INIT=16'b0010011100110011;
    LogicCell40 M_this_sprites_address_q_RNO_0_5_LC_14_21_0 (
            .in0(N__16418),
            .in1(N__13635),
            .in2(N__21472),
            .in3(N__20255),
            .lcout(M_this_sprites_address_q_3_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_3_LC_14_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_3_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_3_LC_14_21_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_3_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__13400),
            .in2(_gnd_net_),
            .in3(N__13300),
            .lcout(\this_vga_signals.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_4_LC_14_21_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_4_LC_14_21_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_4_LC_14_21_2.LUT_INIT=16'b0010011100110011;
    LogicCell40 M_this_sprites_address_q_RNO_0_4_LC_14_21_2 (
            .in0(N__16417),
            .in1(N__13770),
            .in2(N__20120),
            .in3(N__20254),
            .lcout(M_this_sprites_address_q_3_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_2_4_LC_14_22_1.C_ON=1'b0;
    defparam M_this_state_q_RNO_2_4_LC_14_22_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_2_4_LC_14_22_1.LUT_INIT=16'b0000010000000000;
    LogicCell40 M_this_state_q_RNO_2_4_LC_14_22_1 (
            .in0(N__21992),
            .in1(N__13173),
            .in2(N__22447),
            .in3(N__20256),
            .lcout(),
            .ltout(N_206_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_14_22_2.C_ON=1'b0;
    defparam M_this_state_q_4_LC_14_22_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_14_22_2.LUT_INIT=16'b1111110011111110;
    LogicCell40 M_this_state_q_4_LC_14_22_2 (
            .in0(N__13223),
            .in1(N__13229),
            .in2(N__13232),
            .in3(N__14417),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22206),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_3_4_LC_14_22_3.C_ON=1'b0;
    defparam M_this_state_q_RNO_3_4_LC_14_22_3.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_3_4_LC_14_22_3.LUT_INIT=16'b0100010000000000;
    LogicCell40 M_this_state_q_RNO_3_4_LC_14_22_3 (
            .in0(N__21993),
            .in1(N__16277),
            .in2(_gnd_net_),
            .in3(N__16217),
            .lcout(N_207),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_0_4_LC_14_22_6.C_ON=1'b0;
    defparam M_this_state_q_RNO_0_4_LC_14_22_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_0_4_LC_14_22_6.LUT_INIT=16'b0000000000000010;
    LogicCell40 M_this_state_q_RNO_0_4_LC_14_22_6 (
            .in0(N__14407),
            .in1(N__20377),
            .in2(N__20975),
            .in3(N__21991),
            .lcout(M_this_state_q_srsts_0_a2_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIQ80L_0_2_LC_14_23_1.C_ON=1'b0;
    defparam M_this_state_q_RNIQ80L_0_2_LC_14_23_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIQ80L_0_2_LC_14_23_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 M_this_state_q_RNIQ80L_0_2_LC_14_23_1 (
            .in0(N__13174),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(port_dmab_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_0_2_LC_14_23_6.C_ON=1'b0;
    defparam M_this_state_q_RNO_0_2_LC_14_23_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_0_2_LC_14_23_6.LUT_INIT=16'b0000000011101100;
    LogicCell40 M_this_state_q_RNO_0_2_LC_14_23_6 (
            .in0(N__16214),
            .in1(N__20389),
            .in2(N__16249),
            .in3(N__21995),
            .lcout(M_this_state_q_srsts_i_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_3_ns_1_11_LC_14_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_3_ns_1_11_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_3_ns_1_11_LC_14_24_7 .LUT_INIT=16'b0001101100110011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_3_ns_1_11_LC_14_24_7  (
            .in0(N__16411),
            .in1(N__21016),
            .in2(N__20119),
            .in3(N__20290),
            .lcout(\this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNI5CEE4_LC_15_18_6 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNI5CEE4_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNI5CEE4_LC_15_18_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNI5CEE4_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__15101),
            .in2(_gnd_net_),
            .in3(N__15137),
            .lcout(\this_ppu.M_line_clk_out_0 ),
            .ltout(\this_ppu.M_line_clk_out_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIDFVT8_LC_15_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIDFVT8_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIDFVT8_LC_15_18_7 .LUT_INIT=16'b0000000011101111;
    LogicCell40 \this_ppu.M_state_q_RNIDFVT8_LC_15_18_7  (
            .in0(N__19368),
            .in1(N__13460),
            .in2(N__13454),
            .in3(N__21990),
            .lcout(\this_ppu.N_258_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_5_LC_15_21_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_5_LC_15_21_2.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_5_LC_15_21_2.LUT_INIT=16'b0010011100100010;
    LogicCell40 M_this_sprites_address_q_5_LC_15_21_2 (
            .in0(N__17512),
            .in1(N__13451),
            .in2(N__22420),
            .in3(N__13616),
            .lcout(M_this_sprites_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22197),
            .ce(),
            .sr(N__21941));
    defparam M_this_sprites_address_q_4_LC_15_21_3.C_ON=1'b0;
    defparam M_this_sprites_address_q_4_LC_15_21_3.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_4_LC_15_21_3.LUT_INIT=16'b0010011100100010;
    LogicCell40 M_this_sprites_address_q_4_LC_15_21_3 (
            .in0(N__17511),
            .in1(N__13445),
            .in2(N__22419),
            .in3(N__13751),
            .lcout(M_this_sprites_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22197),
            .ce(),
            .sr(N__21941));
    defparam M_this_sprites_address_q_RNO_0_7_LC_15_21_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_7_LC_15_21_4.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_7_LC_15_21_4.LUT_INIT=16'b0001101100110011;
    LogicCell40 M_this_sprites_address_q_RNO_0_7_LC_15_21_4 (
            .in0(N__16415),
            .in1(N__13503),
            .in2(N__20163),
            .in3(N__20335),
            .lcout(),
            .ltout(M_this_sprites_address_q_3_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_7_LC_15_21_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_7_LC_15_21_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_7_LC_15_21_5.LUT_INIT=16'b0001110100001100;
    LogicCell40 M_this_sprites_address_q_7_LC_15_21_5 (
            .in0(N__22365),
            .in1(N__17513),
            .in2(N__13439),
            .in3(N__13484),
            .lcout(M_this_sprites_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22197),
            .ce(),
            .sr(N__21941));
    defparam M_this_sprites_address_q_RNO_1_0_LC_15_22_0.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_0_LC_15_22_0.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_0_LC_15_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_0_LC_15_22_0 (
            .in0(_gnd_net_),
            .in1(N__15283),
            .in2(N__14387),
            .in3(N__14386),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_0),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(un1_M_this_sprites_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_1_LC_15_22_1.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_1_LC_15_22_1.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_1_LC_15_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_1_LC_15_22_1 (
            .in0(_gnd_net_),
            .in1(N__14569),
            .in2(_gnd_net_),
            .in3(N__13436),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_1),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_0),
            .carryout(un1_M_this_sprites_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_2_LC_15_22_2.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_2_LC_15_22_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_2_LC_15_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_2_LC_15_22_2 (
            .in0(_gnd_net_),
            .in1(N__16716),
            .in2(_gnd_net_),
            .in3(N__13433),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_2),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_1),
            .carryout(un1_M_this_sprites_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_3_LC_15_22_3.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_3_LC_15_22_3.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_3_LC_15_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_3_LC_15_22_3 (
            .in0(_gnd_net_),
            .in1(N__17323),
            .in2(_gnd_net_),
            .in3(N__13430),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_3),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_2),
            .carryout(un1_M_this_sprites_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_4_LC_15_22_4.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_4_LC_15_22_4.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_4_LC_15_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_4_LC_15_22_4 (
            .in0(_gnd_net_),
            .in1(N__13771),
            .in2(_gnd_net_),
            .in3(N__13745),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_4),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_3),
            .carryout(un1_M_this_sprites_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_5_LC_15_22_5.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_5_LC_15_22_5.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_5_LC_15_22_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_5_LC_15_22_5 (
            .in0(_gnd_net_),
            .in1(N__13636),
            .in2(_gnd_net_),
            .in3(N__13610),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_5),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_4),
            .carryout(un1_M_this_sprites_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_6_LC_15_22_6.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_6_LC_15_22_6.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_6_LC_15_22_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_6_LC_15_22_6 (
            .in0(_gnd_net_),
            .in1(N__14830),
            .in2(_gnd_net_),
            .in3(N__13607),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_6),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_5),
            .carryout(un1_M_this_sprites_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_7_LC_15_22_7.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_7_LC_15_22_7.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_7_LC_15_22_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_7_LC_15_22_7 (
            .in0(_gnd_net_),
            .in1(N__13504),
            .in2(_gnd_net_),
            .in3(N__13478),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_7),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_6),
            .carryout(un1_M_this_sprites_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_8_LC_15_23_0.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_8_LC_15_23_0.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_8_LC_15_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_8_LC_15_23_0 (
            .in0(_gnd_net_),
            .in1(N__13924),
            .in2(_gnd_net_),
            .in3(N__13475),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_8),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(un1_M_this_sprites_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_9_LC_15_23_1.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_9_LC_15_23_1.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_9_LC_15_23_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_9_LC_15_23_1 (
            .in0(_gnd_net_),
            .in1(N__14704),
            .in2(_gnd_net_),
            .in3(N__13472),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_9),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_8),
            .carryout(un1_M_this_sprites_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_1_10_LC_15_23_2.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNO_1_10_LC_15_23_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_1_10_LC_15_23_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNO_1_10_LC_15_23_2 (
            .in0(_gnd_net_),
            .in1(N__16444),
            .in2(_gnd_net_),
            .in3(N__13469),
            .lcout(M_this_sprites_address_q_RNO_1Z0Z_10),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_9),
            .carryout(un1_M_this_sprites_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_15_23_3.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_15_23_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_15_23_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_15_23_3 (
            .in0(_gnd_net_),
            .in1(N__21015),
            .in2(_gnd_net_),
            .in3(N__13466),
            .lcout(un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_10),
            .carryout(un1_M_this_sprites_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_15_23_4.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_15_23_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_15_23_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_15_23_4 (
            .in0(_gnd_net_),
            .in1(N__21281),
            .in2(_gnd_net_),
            .in3(N__13463),
            .lcout(un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_11),
            .carryout(un1_M_this_sprites_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_15_23_5.C_ON=1'b0;
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_15_23_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_15_23_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_15_23_5 (
            .in0(_gnd_net_),
            .in1(N__21092),
            .in2(_gnd_net_),
            .in3(N__14042),
            .lcout(un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_3_ns_1_12_LC_15_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_3_ns_1_12_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_3_ns_1_12_LC_15_23_6 .LUT_INIT=16'b0000100001111111;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_3_ns_1_12_LC_15_23_6  (
            .in0(N__20325),
            .in1(N__16413),
            .in2(N__21473),
            .in3(N__21282),
            .lcout(\this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_8_LC_15_24_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_8_LC_15_24_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_8_LC_15_24_2.LUT_INIT=16'b0001101100110011;
    LogicCell40 M_this_sprites_address_q_RNO_0_8_LC_15_24_2 (
            .in0(N__16414),
            .in1(N__13923),
            .in2(N__21542),
            .in3(N__20331),
            .lcout(),
            .ltout(M_this_sprites_address_q_3_ns_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_8_LC_15_24_3.C_ON=1'b0;
    defparam M_this_sprites_address_q_8_LC_15_24_3.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_8_LC_15_24_3.LUT_INIT=16'b0000101001001110;
    LogicCell40 M_this_sprites_address_q_8_LC_15_24_3 (
            .in0(N__17509),
            .in1(N__14039),
            .in2(N__14033),
            .in3(N__22422),
            .lcout(M_this_sprites_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22214),
            .ce(),
            .sr(N__21940));
    defparam M_this_sprites_address_q_11_LC_15_24_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_11_LC_15_24_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_11_LC_15_24_5.LUT_INIT=16'b0010011100100010;
    LogicCell40 M_this_sprites_address_q_11_LC_15_24_5 (
            .in0(N__17507),
            .in1(N__13904),
            .in2(N__22448),
            .in3(N__13898),
            .lcout(M_this_sprites_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22214),
            .ce(),
            .sr(N__21940));
    defparam M_this_sprites_address_q_12_LC_15_24_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_12_LC_15_24_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_12_LC_15_24_7.LUT_INIT=16'b0010011100100010;
    LogicCell40 M_this_sprites_address_q_12_LC_15_24_7 (
            .in0(N__17508),
            .in1(N__13892),
            .in2(N__22449),
            .in3(N__13886),
            .lcout(M_this_sprites_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22214),
            .ce(),
            .sr(N__21940));
    defparam M_this_sprites_address_q_1_LC_15_25_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_1_LC_15_25_2.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_1_LC_15_25_2.LUT_INIT=16'b0010011100100010;
    LogicCell40 M_this_sprites_address_q_1_LC_15_25_2 (
            .in0(N__17510),
            .in1(N__14543),
            .in2(N__22450),
            .in3(N__13880),
            .lcout(M_this_sprites_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22217),
            .ce(),
            .sr(N__21937));
    defparam \this_vga_signals.M_lcounter_q_RNIGRI95_1_LC_16_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNIGRI95_1_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNIGRI95_1_LC_16_18_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNIGRI95_1_LC_16_18_1  (
            .in0(N__14334),
            .in1(N__15077),
            .in2(_gnd_net_),
            .in3(N__14118),
            .lcout(\this_vga_signals.un1_M_hcounter_d7_1_0 ),
            .ltout(\this_vga_signals.un1_M_hcounter_d7_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_0_LC_16_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_0_LC_16_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_0_LC_16_18_2 .LUT_INIT=16'b0000011011001100;
    LogicCell40 \this_vga_signals.M_lcounter_q_0_LC_16_18_2  (
            .in0(N__14119),
            .in1(N__14365),
            .in2(N__13871),
            .in3(N__14205),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22176),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_16_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_16_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_1_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__14364),
            .in2(_gnd_net_),
            .in3(N__14117),
            .lcout(),
            .ltout(\this_vga_signals.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_1_LC_16_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_1_LC_16_18_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_1_LC_16_18_4 .LUT_INIT=16'b0011011101000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_1_LC_16_18_4  (
            .in0(N__14345),
            .in1(N__14204),
            .in2(N__14339),
            .in3(N__14335),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22176),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_0_LC_16_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_0_LC_16_18_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_0_LC_16_18_5 .LUT_INIT=16'b1010011000000000;
    LogicCell40 \this_ppu.M_vaddress_q_0_LC_16_18_5  (
            .in0(N__17943),
            .in1(N__14318),
            .in2(N__19385),
            .in3(N__16863),
            .lcout(M_this_ppu_vram_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22176),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_16_20_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_16_20_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_16_20_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__14304),
            .in2(_gnd_net_),
            .in3(N__14312),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22182),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_16_20_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_16_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14303),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22182),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_16_20_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_16_20_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_16_20_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_16_20_3  (
            .in0(N__14306),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14276),
            .lcout(M_this_state_q_nss_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22182),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_16_20_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_16_20_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_16_20_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__14305),
            .in2(_gnd_net_),
            .in3(N__14282),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22182),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_RNIFKS8_1_LC_16_21_0 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_RNIFKS8_1_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \this_pixel_clk.M_counter_q_RNIFKS8_1_LC_16_21_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_pixel_clk.M_counter_q_RNIFKS8_1_LC_16_21_0  (
            .in0(N__14473),
            .in1(N__14964),
            .in2(_gnd_net_),
            .in3(N__21987),
            .lcout(M_counter_q_RNIFKS8_1),
            .ltout(M_counter_q_RNIFKS8_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIMK0K1_9_LC_16_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIMK0K1_9_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIMK0K1_9_LC_16_21_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIMK0K1_9_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14123),
            .in3(N__14101),
            .lcout(\this_vga_signals.M_vcounter_q_249_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_0_LC_16_21_3.C_ON=1'b0;
    defparam M_this_state_q_0_LC_16_21_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_0_LC_16_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_state_q_0_LC_16_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14501),
            .lcout(M_this_state_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22188),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_1_LC_16_21_6 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_1_LC_16_21_6 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_1_LC_16_21_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clk.M_counter_q_1_LC_16_21_6  (
            .in0(N__14474),
            .in1(N__14965),
            .in2(_gnd_net_),
            .in3(N__21988),
            .lcout(\this_pixel_clk.M_counter_q_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22188),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_2_LC_16_22_0.C_ON=1'b0;
    defparam M_this_state_q_2_LC_16_22_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_16_22_0.LUT_INIT=16'b0010000001110000;
    LogicCell40 M_this_state_q_2_LC_16_22_0 (
            .in0(N__16216),
            .in1(N__16276),
            .in2(N__14465),
            .in3(N__20289),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22193),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_6_LC_16_22_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_6_LC_16_22_1.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_6_LC_16_22_1.LUT_INIT=16'b0000001011011111;
    LogicCell40 M_this_sprites_address_q_RNO_0_6_LC_16_22_1 (
            .in0(N__20288),
            .in1(N__16386),
            .in2(N__19796),
            .in3(N__14829),
            .lcout(M_this_sprites_address_q_3_ns_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_rw_iobuf_RNIILOC1_LC_16_22_2.C_ON=1'b0;
    defparam port_rw_iobuf_RNIILOC1_LC_16_22_2.SEQ_MODE=4'b0000;
    defparam port_rw_iobuf_RNIILOC1_LC_16_22_2.LUT_INIT=16'b0000000000001000;
    LogicCell40 port_rw_iobuf_RNIILOC1_LC_16_22_2 (
            .in0(N__14406),
            .in1(N__16248),
            .in2(N__14450),
            .in3(N__21989),
            .lcout(N_218),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_4_4_LC_16_22_4.C_ON=1'b0;
    defparam M_this_state_q_RNO_4_4_LC_16_22_4.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_4_4_LC_16_22_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 M_this_state_q_RNO_4_4_LC_16_22_4 (
            .in0(N__14446),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16247),
            .lcout(),
            .ltout(N_171_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_1_4_LC_16_22_5.C_ON=1'b0;
    defparam M_this_state_q_RNO_1_4_LC_16_22_5.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_1_4_LC_16_22_5.LUT_INIT=16'b0010000010100000;
    LogicCell40 M_this_state_q_RNO_1_4_LC_16_22_5 (
            .in0(N__21764),
            .in1(N__16019),
            .in2(N__14420),
            .in3(N__16045),
            .lcout(N_176_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI95RM1_4_LC_16_22_6.C_ON=1'b0;
    defparam M_this_state_q_RNI95RM1_4_LC_16_22_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI95RM1_4_LC_16_22_6.LUT_INIT=16'b0000010100000100;
    LogicCell40 M_this_state_q_RNI95RM1_4_LC_16_22_6 (
            .in0(N__16215),
            .in1(N__19169),
            .in2(N__14408),
            .in3(N__20287),
            .lcout(N_153_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_2_LC_16_23_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_2_LC_16_23_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_2_LC_16_23_1.LUT_INIT=16'b0001101100001010;
    LogicCell40 M_this_sprites_address_q_2_LC_16_23_1 (
            .in0(N__17494),
            .in1(N__22427),
            .in2(N__16694),
            .in3(N__14372),
            .lcout(M_this_sprites_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22201),
            .ce(),
            .sr(N__21939));
    defparam M_this_sprites_address_q_9_LC_16_23_3.C_ON=1'b0;
    defparam M_this_sprites_address_q_9_LC_16_23_3.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_9_LC_16_23_3.LUT_INIT=16'b0001101100001010;
    LogicCell40 M_this_sprites_address_q_9_LC_16_23_3 (
            .in0(N__17495),
            .in1(N__22428),
            .in2(N__14684),
            .in3(N__14951),
            .lcout(M_this_sprites_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22201),
            .ce(),
            .sr(N__21939));
    defparam M_this_sprites_address_q_13_LC_16_23_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_13_LC_16_23_6.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_13_LC_16_23_6.LUT_INIT=16'b0010011100100010;
    LogicCell40 M_this_sprites_address_q_13_LC_16_23_6 (
            .in0(N__17482),
            .in1(N__16826),
            .in2(N__22452),
            .in3(N__14945),
            .lcout(M_this_sprites_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22201),
            .ce(),
            .sr(N__21939));
    defparam M_this_sprites_address_q_6_LC_16_23_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_6_LC_16_23_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_6_LC_16_23_7.LUT_INIT=16'b0100011101000100;
    LogicCell40 M_this_sprites_address_q_6_LC_16_23_7 (
            .in0(N__14939),
            .in1(N__17483),
            .in2(N__22453),
            .in3(N__14933),
            .lcout(M_this_sprites_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22201),
            .ce(),
            .sr(N__21939));
    defparam M_this_state_q_RNI20CE_0_LC_16_24_1.C_ON=1'b0;
    defparam M_this_state_q_RNI20CE_0_LC_16_24_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI20CE_0_LC_16_24_1.LUT_INIT=16'b1111111110101010;
    LogicCell40 M_this_state_q_RNI20CE_0_LC_16_24_1 (
            .in0(N__22375),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21996),
            .lcout(M_this_state_q_RNI20CEZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_9_LC_16_24_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_9_LC_16_24_5.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_9_LC_16_24_5.LUT_INIT=16'b0001101100110011;
    LogicCell40 M_this_sprites_address_q_RNO_0_9_LC_16_24_5 (
            .in0(N__16410),
            .in1(N__14703),
            .in2(N__19843),
            .in3(N__20327),
            .lcout(M_this_sprites_address_q_3_ns_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_1_LC_16_25_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_1_LC_16_25_6.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_1_LC_16_25_6.LUT_INIT=16'b0000001011011111;
    LogicCell40 M_this_sprites_address_q_RNO_0_1_LC_16_25_6 (
            .in0(N__20326),
            .in1(N__16412),
            .in2(N__21538),
            .in3(N__14562),
            .lcout(M_this_sprites_address_q_3_ns_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI9PQ_4_LC_17_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI9PQ_4_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI9PQ_4_LC_17_17_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \this_ppu.M_haddress_q_RNI9PQ_4_LC_17_17_0  (
            .in0(N__18585),
            .in1(N__17100),
            .in2(N__18430),
            .in3(N__15155),
            .lcout(\this_ppu.un1_M_line_clk_out_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNO_0_4_LC_17_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNO_0_4_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNO_0_4_LC_17_17_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNO_0_4_LC_17_17_4  (
            .in0(N__18901),
            .in1(N__17026),
            .in2(N__17107),
            .in3(N__16120),
            .lcout(),
            .ltout(\this_ppu.un1_M_haddress_q_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_4_LC_17_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_4_LC_17_17_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_4_LC_17_17_5 .LUT_INIT=16'b0110101000000000;
    LogicCell40 \this_ppu.M_haddress_q_4_LC_17_17_5  (
            .in0(N__18433),
            .in1(N__18586),
            .in2(N__14537),
            .in3(N__16174),
            .lcout(M_this_ppu_vram_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22177),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNITAF_6_LC_17_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNITAF_6_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNITAF_6_LC_17_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNITAF_6_LC_17_17_7  (
            .in0(N__18265),
            .in1(N__17021),
            .in2(N__18115),
            .in3(N__18900),
            .lcout(\this_ppu.M_haddress_d8lto6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNI5NOQ4_LC_17_18_3 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNI5NOQ4_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNI5NOQ4_LC_17_18_3 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNI5NOQ4_LC_17_18_3  (
            .in0(N__19367),
            .in1(N__15149),
            .in2(N__15116),
            .in3(N__15143),
            .lcout(\this_ppu.M_last_q_RNI5NOQ4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_1_LC_17_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_1_LC_17_18_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_1_LC_17_18_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_vaddress_q_1_LC_17_18_5  (
            .in0(N__17796),
            .in1(N__16850),
            .in2(_gnd_net_),
            .in3(N__16072),
            .lcout(\this_ppu.M_vaddress_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22180),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIMT2V4_LC_17_19_2 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIMT2V4_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIMT2V4_LC_17_19_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIMT2V4_LC_17_19_2  (
            .in0(N__17939),
            .in1(N__19372),
            .in2(N__15114),
            .in3(N__15138),
            .lcout(\this_ppu.un1_M_vaddress_q_c1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNI2T915_LC_17_19_6 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNI2T915_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNI2T915_LC_17_19_6 .LUT_INIT=16'b0000000011111011;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNI2T915_LC_17_19_6  (
            .in0(N__19373),
            .in1(N__15139),
            .in2(N__15115),
            .in3(N__21994),
            .lcout(\this_ppu.N_250_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRO2H5_9_LC_17_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRO2H5_9_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRO2H5_9_LC_17_20_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIRO2H5_9_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(N__15073),
            .in2(_gnd_net_),
            .in3(N__15019),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNIRO2H5Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_0_LC_17_21_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_0_LC_17_21_0.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_0_LC_17_21_0.LUT_INIT=16'b0010011100100010;
    LogicCell40 M_this_sprites_address_q_0_LC_17_21_0 (
            .in0(N__17506),
            .in1(N__15251),
            .in2(N__22421),
            .in3(N__14978),
            .lcout(M_this_sprites_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22198),
            .ce(),
            .sr(N__21942));
    defparam \this_pixel_clk.M_counter_q_0_LC_17_21_1 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_0_LC_17_21_1 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_0_LC_17_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clk.M_counter_q_0_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14966),
            .lcout(\this_pixel_clk.M_counter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22198),
            .ce(),
            .sr(N__21942));
    defparam M_this_data_count_q_RNIBTAK_10_LC_17_22_1.C_ON=1'b0;
    defparam M_this_data_count_q_RNIBTAK_10_LC_17_22_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIBTAK_10_LC_17_22_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNIBTAK_10_LC_17_22_1 (
            .in0(N__15187),
            .in1(N__15169),
            .in2(N__15419),
            .in3(N__15205),
            .lcout(M_this_state_q_srsts_i_a2_1_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_0_LC_17_22_3.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_0_LC_17_22_3.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_0_LC_17_22_3.LUT_INIT=16'b0100011101010101;
    LogicCell40 M_this_sprites_address_q_RNO_0_0_LC_17_22_3 (
            .in0(N__15270),
            .in1(N__16396),
            .in2(N__20174),
            .in3(N__20281),
            .lcout(M_this_sprites_address_q_3_ns_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIAVRI_11_LC_17_22_4.C_ON=1'b0;
    defparam M_this_data_count_q_RNIAVRI_11_LC_17_22_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIAVRI_11_LC_17_22_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNIAVRI_11_LC_17_22_4 (
            .in0(N__15394),
            .in1(N__15439),
            .in2(N__15956),
            .in3(N__15460),
            .lcout(),
            .ltout(M_this_state_q_srsts_i_a2_1_7_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIDFF62_10_LC_17_22_5.C_ON=1'b0;
    defparam M_this_data_count_q_RNIDFF62_10_LC_17_22_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIDFF62_10_LC_17_22_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_data_count_q_RNIDFF62_10_LC_17_22_5 (
            .in0(N__15236),
            .in1(N__15245),
            .in2(N__15239),
            .in3(N__15230),
            .lcout(N_233),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIAQQL_4_LC_17_22_6.C_ON=1'b0;
    defparam M_this_data_count_q_RNIAQQL_4_LC_17_22_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIAQQL_4_LC_17_22_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNIAQQL_4_LC_17_22_6 (
            .in0(N__15493),
            .in1(N__15511),
            .in2(N__15535),
            .in3(N__15475),
            .lcout(M_this_state_q_srsts_i_a2_1_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIEOD9_13_LC_17_22_7.C_ON=1'b0;
    defparam M_this_data_count_q_RNIEOD9_13_LC_17_22_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIEOD9_13_LC_17_22_7.LUT_INIT=16'b0000000000110011;
    LogicCell40 M_this_data_count_q_RNIEOD9_13_LC_17_22_7 (
            .in0(_gnd_net_),
            .in1(N__15220),
            .in2(_gnd_net_),
            .in3(N__15557),
            .lcout(M_this_state_q_srsts_i_a2_1_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_0_LC_17_23_0.C_ON=1'b1;
    defparam M_this_data_count_q_0_LC_17_23_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_17_23_0.LUT_INIT=16'b0011110000111100;
    LogicCell40 M_this_data_count_q_0_LC_17_23_0 (
            .in0(_gnd_net_),
            .in1(N__20923),
            .in2(N__15224),
            .in3(_gnd_net_),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(un1_M_this_data_count_q_cry_0),
            .clk(N__22207),
            .ce(),
            .sr(N__15932));
    defparam M_this_data_count_q_1_LC_17_23_1.C_ON=1'b1;
    defparam M_this_data_count_q_1_LC_17_23_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_17_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_1_LC_17_23_1 (
            .in0(_gnd_net_),
            .in1(N__20927),
            .in2(N__15209),
            .in3(N__15194),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_0),
            .carryout(un1_M_this_data_count_q_cry_1),
            .clk(N__22207),
            .ce(),
            .sr(N__15932));
    defparam M_this_data_count_q_2_LC_17_23_2.C_ON=1'b1;
    defparam M_this_data_count_q_2_LC_17_23_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_17_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_2_LC_17_23_2 (
            .in0(_gnd_net_),
            .in1(N__20924),
            .in2(N__15191),
            .in3(N__15176),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_1),
            .carryout(un1_M_this_data_count_q_cry_2),
            .clk(N__22207),
            .ce(),
            .sr(N__15932));
    defparam M_this_data_count_q_3_LC_17_23_3.C_ON=1'b1;
    defparam M_this_data_count_q_3_LC_17_23_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_17_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_3_LC_17_23_3 (
            .in0(_gnd_net_),
            .in1(N__20928),
            .in2(N__15173),
            .in3(N__15158),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_2),
            .carryout(un1_M_this_data_count_q_cry_3),
            .clk(N__22207),
            .ce(),
            .sr(N__15932));
    defparam M_this_data_count_q_4_LC_17_23_4.C_ON=1'b1;
    defparam M_this_data_count_q_4_LC_17_23_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_17_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_4_LC_17_23_4 (
            .in0(_gnd_net_),
            .in1(N__20925),
            .in2(N__15536),
            .in3(N__15518),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_3),
            .carryout(un1_M_this_data_count_q_cry_4),
            .clk(N__22207),
            .ce(),
            .sr(N__15932));
    defparam M_this_data_count_q_5_LC_17_23_5.C_ON=1'b1;
    defparam M_this_data_count_q_5_LC_17_23_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_17_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_5_LC_17_23_5 (
            .in0(_gnd_net_),
            .in1(N__20929),
            .in2(N__15515),
            .in3(N__15500),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_4),
            .carryout(un1_M_this_data_count_q_cry_5),
            .clk(N__22207),
            .ce(),
            .sr(N__15932));
    defparam M_this_data_count_q_6_LC_17_23_6.C_ON=1'b1;
    defparam M_this_data_count_q_6_LC_17_23_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_17_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_6_LC_17_23_6 (
            .in0(_gnd_net_),
            .in1(N__20926),
            .in2(N__15497),
            .in3(N__15482),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_5),
            .carryout(un1_M_this_data_count_q_cry_6),
            .clk(N__22207),
            .ce(),
            .sr(N__15932));
    defparam M_this_data_count_q_7_LC_17_23_7.C_ON=1'b1;
    defparam M_this_data_count_q_7_LC_17_23_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_17_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_7_LC_17_23_7 (
            .in0(_gnd_net_),
            .in1(N__20930),
            .in2(N__15479),
            .in3(N__15464),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_6),
            .carryout(un1_M_this_data_count_q_cry_7),
            .clk(N__22207),
            .ce(),
            .sr(N__15932));
    defparam M_this_data_count_q_8_LC_17_24_0.C_ON=1'b1;
    defparam M_this_data_count_q_8_LC_17_24_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_17_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_8_LC_17_24_0 (
            .in0(_gnd_net_),
            .in1(N__20958),
            .in2(N__15461),
            .in3(N__15443),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(bfn_17_24_0_),
            .carryout(un1_M_this_data_count_q_cry_8),
            .clk(N__22215),
            .ce(),
            .sr(N__15925));
    defparam M_this_data_count_q_9_LC_17_24_1.C_ON=1'b1;
    defparam M_this_data_count_q_9_LC_17_24_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_17_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_9_LC_17_24_1 (
            .in0(_gnd_net_),
            .in1(N__20961),
            .in2(N__15440),
            .in3(N__15422),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_8),
            .carryout(un1_M_this_data_count_q_cry_9),
            .clk(N__22215),
            .ce(),
            .sr(N__15925));
    defparam M_this_data_count_q_10_LC_17_24_2.C_ON=1'b1;
    defparam M_this_data_count_q_10_LC_17_24_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_17_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_10_LC_17_24_2 (
            .in0(_gnd_net_),
            .in1(N__20959),
            .in2(N__15418),
            .in3(N__15398),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_9),
            .carryout(un1_M_this_data_count_q_cry_10),
            .clk(N__22215),
            .ce(),
            .sr(N__15925));
    defparam M_this_data_count_q_11_LC_17_24_3.C_ON=1'b1;
    defparam M_this_data_count_q_11_LC_17_24_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_17_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_11_LC_17_24_3 (
            .in0(_gnd_net_),
            .in1(N__20962),
            .in2(N__15395),
            .in3(N__15377),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_10),
            .carryout(un1_M_this_data_count_q_cry_11),
            .clk(N__22215),
            .ce(),
            .sr(N__15925));
    defparam M_this_data_count_q_12_LC_17_24_4.C_ON=1'b1;
    defparam M_this_data_count_q_12_LC_17_24_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_17_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_12_LC_17_24_4 (
            .in0(_gnd_net_),
            .in1(N__20960),
            .in2(N__15955),
            .in3(N__15935),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_11),
            .carryout(un1_M_this_data_count_q_cry_12),
            .clk(N__22215),
            .ce(),
            .sr(N__15925));
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_17_24_5.C_ON=1'b1;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_17_24_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_17_24_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_17_24_5 (
            .in0(_gnd_net_),
            .in1(N__15668),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_12),
            .carryout(un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_17_24_6.C_ON=1'b1;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_17_24_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_17_24_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_17_24_6 (
            .in0(_gnd_net_),
            .in1(N__15670),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO),
            .carryout(un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_17_24_7.C_ON=1'b1;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_17_24_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_17_24_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_17_24_7 (
            .in0(_gnd_net_),
            .in1(N__15669),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO),
            .carryout(un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_17_25_0.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_17_25_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_17_25_0.LUT_INIT=16'b1110101110111110;
    LogicCell40 M_this_data_count_q_13_LC_17_25_0 (
            .in0(N__22435),
            .in1(N__15556),
            .in2(N__20973),
            .in3(N__15560),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22218),
            .ce(),
            .sr(N__21938));
    defparam \this_ppu.M_haddress_q_RNIU60R4_1_LC_18_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIU60R4_1_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIU60R4_1_LC_18_17_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNIU60R4_1_LC_18_17_1  (
            .in0(N__17085),
            .in1(N__18903),
            .in2(_gnd_net_),
            .in3(N__16119),
            .lcout(\this_ppu.un1_M_haddress_q_c2 ),
            .ltout(\this_ppu.un1_M_haddress_q_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIBMBR4_4_LC_18_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIBMBR4_4_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIBMBR4_4_LC_18_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNIBMBR4_4_LC_18_17_2  (
            .in0(N__18432),
            .in1(N__18590),
            .in2(N__15542),
            .in3(N__17025),
            .lcout(\this_ppu.un1_M_haddress_q_c5 ),
            .ltout(\this_ppu.un1_M_haddress_q_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_6_LC_18_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_6_LC_18_17_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_6_LC_18_17_3 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \this_ppu.M_haddress_q_6_LC_18_17_3  (
            .in0(N__16161),
            .in1(N__18114),
            .in2(N__15539),
            .in3(N__18270),
            .lcout(M_this_ppu_vram_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22181),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_2_LC_18_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_2_LC_18_17_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_2_LC_18_17_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_haddress_q_2_LC_18_17_4  (
            .in0(N__17027),
            .in1(N__16158),
            .in2(_gnd_net_),
            .in3(N__16081),
            .lcout(M_this_ppu_vram_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22181),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_5_LC_18_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_5_LC_18_17_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_5_LC_18_17_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_ppu.M_haddress_q_5_LC_18_17_5  (
            .in0(N__16159),
            .in1(N__18269),
            .in2(_gnd_net_),
            .in3(N__16088),
            .lcout(M_this_ppu_vram_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22181),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_3_LC_18_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_3_LC_18_17_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_3_LC_18_17_6 .LUT_INIT=16'b0100100010001000;
    LogicCell40 \this_ppu.M_haddress_q_3_LC_18_17_6  (
            .in0(N__18591),
            .in1(N__16160),
            .in2(N__17035),
            .in3(N__16082),
            .lcout(M_this_ppu_vram_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22181),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_4_LC_18_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_4_LC_18_18_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_4_LC_18_18_5 .LUT_INIT=16'b0100100011000000;
    LogicCell40 \this_ppu.M_vaddress_q_4_LC_18_18_5  (
            .in0(N__19127),
            .in1(N__16865),
            .in2(N__18989),
            .in3(N__16103),
            .lcout(\this_ppu.M_vaddress_qZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22184),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_2_LC_18_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_2_LC_18_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_2_LC_18_18_7 .LUT_INIT=16'b0100100011000000;
    LogicCell40 \this_ppu.M_vaddress_q_2_LC_18_18_7  (
            .in0(N__17797),
            .in1(N__16864),
            .in2(N__17654),
            .in3(N__16073),
            .lcout(\this_ppu.M_vaddress_qZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22184),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNID0D95_2_LC_18_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNID0D95_2_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNID0D95_2_LC_18_19_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNID0D95_2_LC_18_19_3  (
            .in0(N__17646),
            .in1(N__17792),
            .in2(_gnd_net_),
            .in3(N__16071),
            .lcout(\this_ppu.un1_M_vaddress_q_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_5_LC_18_22_0.C_ON=1'b0;
    defparam M_this_state_q_5_LC_18_22_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_18_22_0.LUT_INIT=16'b1100110011011100;
    LogicCell40 M_this_state_q_5_LC_18_22_0 (
            .in0(N__20286),
            .in1(N__15962),
            .in2(N__16404),
            .in3(N__22000),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22208),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_0_7_LC_18_22_3.C_ON=1'b0;
    defparam M_this_state_q_RNO_0_7_LC_18_22_3.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_0_7_LC_18_22_3.LUT_INIT=16'b0100000000000000;
    LogicCell40 M_this_state_q_RNO_0_7_LC_18_22_3 (
            .in0(N__16055),
            .in1(N__16018),
            .in2(N__21767),
            .in3(N__15977),
            .lcout(N_200),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_0_6_LC_18_22_5.C_ON=1'b0;
    defparam M_this_state_q_RNO_0_6_LC_18_22_5.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_0_6_LC_18_22_5.LUT_INIT=16'b0010000000000000;
    LogicCell40 M_this_state_q_RNO_0_6_LC_18_22_5 (
            .in0(N__16054),
            .in1(N__16017),
            .in2(N__21766),
            .in3(N__15976),
            .lcout(N_202),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_0_5_LC_18_22_7.C_ON=1'b0;
    defparam M_this_state_q_RNO_0_5_LC_18_22_7.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_0_5_LC_18_22_7.LUT_INIT=16'b0001000000000000;
    LogicCell40 M_this_state_q_RNO_0_5_LC_18_22_7 (
            .in0(N__16053),
            .in1(N__16016),
            .in2(N__21765),
            .in3(N__15975),
            .lcout(N_204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_6_LC_18_23_1.C_ON=1'b0;
    defparam M_this_state_q_6_LC_18_23_1.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_18_23_1.LUT_INIT=16'b1100110111001100;
    LogicCell40 M_this_state_q_6_LC_18_23_1 (
            .in0(N__21999),
            .in1(N__16292),
            .in2(N__20336),
            .in3(N__16286),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22216),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIVD0L_6_LC_18_23_3.C_ON=1'b0;
    defparam M_this_state_q_RNIVD0L_6_LC_18_23_3.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIVD0L_6_LC_18_23_3.LUT_INIT=16'b0000000011101110;
    LogicCell40 M_this_state_q_RNIVD0L_6_LC_18_23_3 (
            .in0(N__16375),
            .in1(N__16285),
            .in2(_gnd_net_),
            .in3(N__22395),
            .lcout(M_this_sprites_address_q_3_sm0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_0_1_LC_18_23_5.C_ON=1'b0;
    defparam M_this_state_q_RNO_0_1_LC_18_23_5.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_0_1_LC_18_23_5.LUT_INIT=16'b0001000100000000;
    LogicCell40 M_this_state_q_RNO_0_1_LC_18_23_5 (
            .in0(N__16275),
            .in1(N__16256),
            .in2(_gnd_net_),
            .in3(N__16204),
            .lcout(),
            .ltout(M_this_state_q_srsts_i_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_1_LC_18_23_6.C_ON=1'b0;
    defparam M_this_state_q_1_LC_18_23_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_18_23_6.LUT_INIT=16'b0000000011111110;
    LogicCell40 M_this_state_q_1_LC_18_23_6 (
            .in0(N__22396),
            .in1(N__20952),
            .in2(N__16220),
            .in3(N__21998),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22216),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_1_LC_19_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_1_LC_19_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_1_LC_19_17_2 .LUT_INIT=16'b0110000011000000;
    LogicCell40 \this_ppu.M_haddress_q_1_LC_19_17_2  (
            .in0(N__18896),
            .in1(N__17086),
            .in2(N__16175),
            .in3(N__16133),
            .lcout(M_this_ppu_vram_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22185),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_0_LC_19_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_0_LC_19_17_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_0_LC_19_17_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_haddress_q_0_LC_19_17_3  (
            .in0(N__16132),
            .in1(N__16170),
            .in2(_gnd_net_),
            .in3(N__18895),
            .lcout(M_this_ppu_vram_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22185),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_LC_19_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_LC_19_17_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_LC_19_17_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_state_q_LC_19_17_6  (
            .in0(_gnd_net_),
            .in1(N__16131),
            .in2(_gnd_net_),
            .in3(N__21997),
            .lcout(M_this_ppu_vram_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22185),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_6_LC_19_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_6_LC_19_18_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_6_LC_19_18_0 .LUT_INIT=16'b0010100010100000;
    LogicCell40 \this_ppu.M_vaddress_q_6_LC_19_18_0  (
            .in0(N__16868),
            .in1(N__18962),
            .in2(N__18941),
            .in3(N__16874),
            .lcout(\this_ppu.M_vaddress_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22192),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_3_LC_19_18_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_3_LC_19_18_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_3_LC_19_18_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_vaddress_q_3_LC_19_18_3  (
            .in0(N__19124),
            .in1(N__16866),
            .in2(_gnd_net_),
            .in3(N__16102),
            .lcout(\this_ppu.M_vaddress_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22192),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNI87NJ5_4_LC_19_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNI87NJ5_4_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNI87NJ5_4_LC_19_18_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNI87NJ5_4_LC_19_18_5  (
            .in0(N__18981),
            .in1(N__19126),
            .in2(_gnd_net_),
            .in3(N__16101),
            .lcout(\this_ppu.un1_M_vaddress_q_c5 ),
            .ltout(\this_ppu.un1_M_vaddress_q_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_5_LC_19_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_5_LC_19_18_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_5_LC_19_18_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \this_ppu.M_vaddress_q_5_LC_19_18_6  (
            .in0(N__16867),
            .in1(_gnd_net_),
            .in2(N__16829),
            .in3(N__18961),
            .lcout(\this_ppu.M_vaddress_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22192),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_3_ns_1_13_LC_19_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_3_ns_1_13_LC_19_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_3_ns_1_13_LC_19_23_3 .LUT_INIT=16'b0001110101010101;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_3_ns_1_13_LC_19_23_3  (
            .in0(N__21106),
            .in1(N__16371),
            .in2(N__19795),
            .in3(N__20322),
            .lcout(\this_vga_signals.M_this_sprites_address_q_3_ns_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_2_LC_19_24_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_2_LC_19_24_1.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_2_LC_19_24_1.LUT_INIT=16'b0010011100110011;
    LogicCell40 M_this_sprites_address_q_RNO_0_2_LC_19_24_1 (
            .in0(N__16385),
            .in1(N__16726),
            .in2(N__19844),
            .in3(N__20321),
            .lcout(M_this_sprites_address_q_3_ns_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI84774_LC_20_11_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI84774_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI84774_LC_20_11_3 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \this_ppu.M_state_q_RNI84774_LC_20_11_3  (
            .in0(N__19378),
            .in1(N__18617),
            .in2(N__19278),
            .in3(N__17216),
            .lcout(M_this_ppu_vram_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIPF7_1_LC_20_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIPF7_1_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIPF7_1_LC_20_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_haddress_q_RNIPF7_1_LC_20_17_3  (
            .in0(_gnd_net_),
            .in1(N__17081),
            .in2(_gnd_net_),
            .in3(N__18894),
            .lcout(M_this_ppu_sprites_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_10_LC_20_22_3.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_10_LC_20_22_3.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_10_LC_20_22_3.LUT_INIT=16'b0001110101010101;
    LogicCell40 M_this_sprites_address_q_RNO_0_10_LC_20_22_3 (
            .in0(N__16437),
            .in1(N__16400),
            .in2(N__19985),
            .in3(N__20282),
            .lcout(M_this_sprites_address_q_3_ns_1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_10_LC_20_23_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_10_LC_20_23_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_10_LC_20_23_1.LUT_INIT=16'b0010011100100010;
    LogicCell40 M_this_sprites_address_q_10_LC_20_23_1 (
            .in0(N__17504),
            .in1(N__16556),
            .in2(N__22451),
            .in3(N__16550),
            .lcout(M_this_sprites_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22222),
            .ce(),
            .sr(N__21943));
    defparam M_this_sprites_address_q_RNO_0_3_LC_20_23_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_3_LC_20_23_4.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_3_LC_20_23_4.LUT_INIT=16'b0001101100001111;
    LogicCell40 M_this_sprites_address_q_RNO_0_3_LC_20_23_4 (
            .in0(N__16416),
            .in1(N__19971),
            .in2(N__17313),
            .in3(N__20323),
            .lcout(),
            .ltout(M_this_sprites_address_q_3_ns_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_3_LC_20_23_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_3_LC_20_23_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_3_LC_20_23_5.LUT_INIT=16'b0001101100001010;
    LogicCell40 M_this_sprites_address_q_3_LC_20_23_5 (
            .in0(N__17505),
            .in1(N__22423),
            .in2(N__17432),
            .in3(N__17429),
            .lcout(M_this_sprites_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22222),
            .ce(),
            .sr(N__21943));
    defparam M_this_state_q_3_LC_20_23_6.C_ON=1'b0;
    defparam M_this_state_q_3_LC_20_23_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_20_23_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 M_this_state_q_3_LC_20_23_6 (
            .in0(_gnd_net_),
            .in1(N__20390),
            .in2(_gnd_net_),
            .in3(N__20324),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22222),
            .ce(),
            .sr(N__21943));
    defparam \this_sprites_ram.mem_mem_1_1_RNIJBQ01_0_LC_21_10_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNIJBQ01_0_LC_21_10_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNIJBQ01_0_LC_21_10_3 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNIJBQ01_0_LC_21_10_3  (
            .in0(N__20495),
            .in1(N__17285),
            .in2(N__20672),
            .in3(N__17267),
            .lcout(\this_sprites_ram.mem_DOUT_6_i_m2_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIDT2Q1_0_LC_21_11_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIDT2Q1_0_LC_21_11_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIDT2Q1_0_LC_21_11_7 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIDT2Q1_0_LC_21_11_7  (
            .in0(N__17255),
            .in1(N__20530),
            .in2(N__17240),
            .in3(N__17222),
            .lcout(this_sprites_ram_mem_N_102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI04774_LC_21_13_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI04774_LC_21_13_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI04774_LC_21_13_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \this_ppu.M_state_q_RNI04774_LC_21_13_5  (
            .in0(N__19374),
            .in1(N__18683),
            .in2(N__19268),
            .in3(N__17156),
            .lcout(M_this_ppu_vram_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNI5LUP1_0_LC_21_14_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNI5LUP1_0_LC_21_14_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNI5LUP1_0_LC_21_14_3 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNI5LUP1_0_LC_21_14_3  (
            .in0(N__17192),
            .in1(N__20546),
            .in2(N__17177),
            .in3(N__17120),
            .lcout(this_sprites_ram_mem_N_91),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIF7O01_0_LC_21_15_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIF7O01_0_LC_21_15_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIF7O01_0_LC_21_15_1 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIF7O01_0_LC_21_15_1  (
            .in0(N__20496),
            .in1(N__17150),
            .in2(N__20657),
            .in3(N__17138),
            .lcout(\this_sprites_ram.mem_DOUT_3_i_m2_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_cry_1_c_LC_21_17_0 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_cry_1_c_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_cry_1_c_LC_21_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.sprites_addr_cry_1_c_LC_21_17_0  (
            .in0(_gnd_net_),
            .in1(N__18902),
            .in2(N__17099),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_21_17_0_),
            .carryout(\this_ppu.sprites_addr_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_cry_1_c_RNIB25D_LC_21_17_1 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_cry_1_c_RNIB25D_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_cry_1_c_RNIB25D_LC_21_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.sprites_addr_cry_1_c_RNIB25D_LC_21_17_1  (
            .in0(_gnd_net_),
            .in1(N__17031),
            .in2(_gnd_net_),
            .in3(N__18605),
            .lcout(M_this_ppu_sprites_addr_2),
            .ltout(),
            .carryin(\this_ppu.sprites_addr_cry_1 ),
            .carryout(\this_ppu.sprites_addr_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_cry_2_c_RNID56D_LC_21_17_2 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_cry_2_c_RNID56D_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_cry_2_c_RNID56D_LC_21_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.sprites_addr_cry_2_c_RNID56D_LC_21_17_2  (
            .in0(_gnd_net_),
            .in1(N__18595),
            .in2(_gnd_net_),
            .in3(N__18446),
            .lcout(M_this_ppu_sprites_addr_3),
            .ltout(),
            .carryin(\this_ppu.sprites_addr_cry_2 ),
            .carryout(\this_ppu.sprites_addr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_cry_3_c_RNIF87D_LC_21_17_3 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_cry_3_c_RNIF87D_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_cry_3_c_RNIF87D_LC_21_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.sprites_addr_cry_3_c_RNIF87D_LC_21_17_3  (
            .in0(_gnd_net_),
            .in1(N__18431),
            .in2(_gnd_net_),
            .in3(N__18284),
            .lcout(M_this_ppu_sprites_addr_4),
            .ltout(),
            .carryin(\this_ppu.sprites_addr_cry_3 ),
            .carryout(\this_ppu.sprites_addr_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_cry_4_c_RNIHB8D_LC_21_17_4 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_cry_4_c_RNIHB8D_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_cry_4_c_RNIHB8D_LC_21_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.sprites_addr_cry_4_c_RNIHB8D_LC_21_17_4  (
            .in0(_gnd_net_),
            .in1(N__18274),
            .in2(_gnd_net_),
            .in3(N__18131),
            .lcout(M_this_ppu_sprites_addr_5),
            .ltout(),
            .carryin(\this_ppu.sprites_addr_cry_4 ),
            .carryout(\this_ppu.sprites_addr_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_cry_5_c_RNIJE9D_LC_21_17_5 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_cry_5_c_RNIJE9D_LC_21_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_cry_5_c_RNIJE9D_LC_21_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.sprites_addr_cry_5_c_RNIJE9D_LC_21_17_5  (
            .in0(_gnd_net_),
            .in1(N__18113),
            .in2(_gnd_net_),
            .in3(N__17969),
            .lcout(M_this_ppu_sprites_addr_6),
            .ltout(),
            .carryin(\this_ppu.sprites_addr_cry_5 ),
            .carryout(\this_ppu.sprites_addr_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_cry_6_c_RNISIBI_LC_21_17_6 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_cry_6_c_RNISIBI_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_cry_6_c_RNISIBI_LC_21_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.sprites_addr_cry_6_c_RNISIBI_LC_21_17_6  (
            .in0(_gnd_net_),
            .in1(N__17959),
            .in2(_gnd_net_),
            .in3(N__17804),
            .lcout(M_this_ppu_sprites_addr_7),
            .ltout(),
            .carryin(\this_ppu.sprites_addr_cry_6 ),
            .carryout(\this_ppu.sprites_addr_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_cry_7_c_RNIULCI_LC_21_17_7 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_cry_7_c_RNIULCI_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_cry_7_c_RNIULCI_LC_21_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.sprites_addr_cry_7_c_RNIULCI_LC_21_17_7  (
            .in0(_gnd_net_),
            .in1(N__17801),
            .in2(_gnd_net_),
            .in3(N__17657),
            .lcout(M_this_ppu_sprites_addr_8),
            .ltout(),
            .carryin(\this_ppu.sprites_addr_cry_7 ),
            .carryout(\this_ppu.sprites_addr_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_cry_8_c_RNI0PDI_LC_21_18_0 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_cry_8_c_RNI0PDI_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_cry_8_c_RNI0PDI_LC_21_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.sprites_addr_cry_8_c_RNI0PDI_LC_21_18_0  (
            .in0(_gnd_net_),
            .in1(N__17653),
            .in2(_gnd_net_),
            .in3(N__17516),
            .lcout(M_this_ppu_sprites_addr_9),
            .ltout(),
            .carryin(bfn_21_18_0_),
            .carryout(\this_ppu.sprites_addr_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_cry_9_c_RNI2SEI_LC_21_18_1 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_cry_9_c_RNI2SEI_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_cry_9_c_RNI2SEI_LC_21_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.sprites_addr_cry_9_c_RNI2SEI_LC_21_18_1  (
            .in0(_gnd_net_),
            .in1(N__19125),
            .in2(_gnd_net_),
            .in3(N__18992),
            .lcout(M_this_ppu_sprites_addr_10),
            .ltout(),
            .carryin(\this_ppu.sprites_addr_cry_9 ),
            .carryout(\this_ppu.sprites_addr_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_11_LC_21_18_2 .C_ON=1'b1;
    defparam \this_sprites_ram.mem_radreg_11_LC_21_18_2 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_11_LC_21_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_sprites_ram.mem_radreg_11_LC_21_18_2  (
            .in0(_gnd_net_),
            .in1(N__18988),
            .in2(_gnd_net_),
            .in3(N__18965),
            .lcout(this_sprites_ram_mem_radreg_11),
            .ltout(),
            .carryin(\this_ppu.sprites_addr_cry_10 ),
            .carryout(\this_ppu.sprites_addr_cry_11 ),
            .clk(N__22203),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_12_LC_21_18_3 .C_ON=1'b1;
    defparam \this_sprites_ram.mem_radreg_12_LC_21_18_3 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_12_LC_21_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_sprites_ram.mem_radreg_12_LC_21_18_3  (
            .in0(_gnd_net_),
            .in1(N__18960),
            .in2(_gnd_net_),
            .in3(N__18944),
            .lcout(\this_sprites_ram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(\this_ppu.sprites_addr_cry_11 ),
            .carryout(\this_ppu.sprites_addr_cry_12 ),
            .clk(N__22203),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_13_LC_21_18_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_13_LC_21_18_4 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_13_LC_21_18_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_sprites_ram.mem_radreg_13_LC_21_18_4  (
            .in0(_gnd_net_),
            .in1(N__18937),
            .in2(_gnd_net_),
            .in3(N__18923),
            .lcout(\this_sprites_ram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22203),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNICN3_0_LC_21_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNICN3_0_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNICN3_0_LC_21_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.M_haddress_q_RNICN3_0_LC_21_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18910),
            .lcout(M_this_ppu_vram_addr_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNIHBQ01_0_LC_22_13_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNIHBQ01_0_LC_22_13_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNIHBQ01_0_LC_22_13_2 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNIHBQ01_0_LC_22_13_2  (
            .in0(N__20535),
            .in1(N__18743),
            .in2(N__20683),
            .in3(N__18731),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_6_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNI9T2Q1_0_LC_22_13_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNI9T2Q1_0_LC_22_13_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNI9T2Q1_0_LC_22_13_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNI9T2Q1_0_LC_22_13_3  (
            .in0(N__18716),
            .in1(N__18695),
            .in2(N__18686),
            .in3(N__20536),
            .lcout(this_sprites_ram_mem_N_88),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_22_13_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_22_13_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_22_13_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_wclke_3_LC_22_13_6  (
            .in0(N__21338),
            .in1(N__21076),
            .in2(N__21183),
            .in3(N__21257),
            .lcout(\this_sprites_ram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNI9LUP1_0_LC_22_15_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNI9LUP1_0_LC_22_15_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNI9LUP1_0_LC_22_15_5 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNI9LUP1_0_LC_22_15_5  (
            .in0(N__18647),
            .in1(N__20534),
            .in2(N__18635),
            .in3(N__19190),
            .lcout(this_sprites_ram_mem_N_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_22_22_0.C_ON=1'b0;
    defparam M_this_state_q_7_LC_22_22_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_22_22_0.LUT_INIT=16'b1111000011110100;
    LogicCell40 M_this_state_q_7_LC_22_22_0 (
            .in0(N__20258),
            .in1(N__19184),
            .in2(N__19421),
            .in3(N__22001),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22224),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIB2RF1_3_LC_22_22_3.C_ON=1'b0;
    defparam M_this_state_q_RNIB2RF1_3_LC_22_22_3.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIB2RF1_3_LC_22_22_3.LUT_INIT=16'b0100010001010101;
    LogicCell40 M_this_state_q_RNIB2RF1_3_LC_22_22_3 (
            .in0(N__20953),
            .in1(N__19165),
            .in2(_gnd_net_),
            .in3(N__20257),
            .lcout(M_this_sprites_ram_write_en_1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI84774_0_LC_23_9_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI84774_0_LC_23_9_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI84774_0_LC_23_9_3 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \this_ppu.M_state_q_RNI84774_0_LC_23_9_3  (
            .in0(N__19391),
            .in1(N__19619),
            .in2(N__19289),
            .in3(N__20447),
            .lcout(M_this_ppu_vram_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI04774_0_LC_23_10_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI04774_0_LC_23_10_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI04774_0_LC_23_10_3 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \this_ppu.M_state_q_RNI04774_0_LC_23_10_3  (
            .in0(N__19387),
            .in1(N__19493),
            .in2(N__19285),
            .in3(N__19556),
            .lcout(M_this_ppu_vram_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIH7O01_0_LC_23_15_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIH7O01_0_LC_23_15_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIH7O01_0_LC_23_15_1 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIH7O01_0_LC_23_15_1  (
            .in0(N__20531),
            .in1(N__19217),
            .in2(N__20674),
            .in3(N__19205),
            .lcout(\this_sprites_ram.mem_DOUT_3_i_m2_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIDVQ81_7_LC_23_22_1.C_ON=1'b0;
    defparam M_this_state_q_RNIDVQ81_7_LC_23_22_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIDVQ81_7_LC_23_22_1.LUT_INIT=16'b0001000100110011;
    LogicCell40 M_this_state_q_RNIDVQ81_7_LC_23_22_1 (
            .in0(N__19183),
            .in1(N__20954),
            .in2(_gnd_net_),
            .in3(N__20262),
            .lcout(un1_M_this_state_q_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI1B0E_7_LC_23_22_2.C_ON=1'b0;
    defparam M_this_state_q_RNI1B0E_7_LC_23_22_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI1B0E_7_LC_23_22_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 M_this_state_q_RNI1B0E_7_LC_23_22_2 (
            .in0(_gnd_net_),
            .in1(N__19182),
            .in2(_gnd_net_),
            .in3(N__20373),
            .lcout(N_170_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_23_24_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_23_24_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_23_24_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_sprites_ram.mem_mem_7_0_wclke_3_LC_23_24_3  (
            .in0(N__21300),
            .in1(N__21029),
            .in2(N__21156),
            .in3(N__21234),
            .lcout(\this_sprites_ram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIH7O01_LC_24_10_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIH7O01_LC_24_10_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIH7O01_LC_24_10_0 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIH7O01_LC_24_10_0  (
            .in0(N__20547),
            .in1(N__19676),
            .in2(N__20673),
            .in3(N__19661),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_3_i_m2_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNI9LUP1_LC_24_10_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNI9LUP1_LC_24_10_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNI9LUP1_LC_24_10_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNI9LUP1_LC_24_10_1  (
            .in0(N__19649),
            .in1(N__19631),
            .in2(N__19622),
            .in3(N__20548),
            .lcout(this_sprites_ram_mem_N_98),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNIHBQ01_LC_24_11_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNIHBQ01_LC_24_11_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNIHBQ01_LC_24_11_1 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNIHBQ01_LC_24_11_1  (
            .in0(N__20549),
            .in1(N__19613),
            .in2(N__20684),
            .in3(N__19598),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_6_i_m2_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNI9T2Q1_LC_24_11_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNI9T2Q1_LC_24_11_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNI9T2Q1_LC_24_11_2 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNI9T2Q1_LC_24_11_2  (
            .in0(N__19586),
            .in1(N__19577),
            .in2(N__19559),
            .in3(N__20551),
            .lcout(this_sprites_ram_mem_N_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIF7O01_LC_24_11_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIF7O01_LC_24_11_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIF7O01_LC_24_11_4 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIF7O01_LC_24_11_4  (
            .in0(N__19550),
            .in1(N__20682),
            .in2(N__19535),
            .in3(N__20550),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_3_i_m2_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNI5LUP1_LC_24_11_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNI5LUP1_LC_24_11_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNI5LUP1_LC_24_11_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNI5LUP1_LC_24_11_5  (
            .in0(N__20552),
            .in1(N__19517),
            .in2(N__19502),
            .in3(N__19499),
            .lcout(this_sprites_ram_mem_N_112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_14_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_14_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_14_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_14_0  (
            .in0(N__21326),
            .in1(N__21072),
            .in2(N__21185),
            .in3(N__21259),
            .lcout(\this_sprites_ram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_14_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_14_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_14_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_14_1  (
            .in0(N__21260),
            .in1(N__21182),
            .in2(N__21077),
            .in3(N__21327),
            .lcout(\this_sprites_ram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_14_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_14_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_14_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_14_2  (
            .in0(N__21325),
            .in1(N__21071),
            .in2(N__21184),
            .in3(N__21258),
            .lcout(\this_sprites_ram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNIJBQ01_LC_24_15_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNIJBQ01_LC_24_15_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNIJBQ01_LC_24_15_5 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNIJBQ01_LC_24_15_5  (
            .in0(N__20532),
            .in1(N__20696),
            .in2(N__20678),
            .in3(N__20588),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_6_i_m2_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIDT2Q1_LC_24_15_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIDT2Q1_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIDT2Q1_LC_24_15_6 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIDT2Q1_LC_24_15_6  (
            .in0(N__20576),
            .in1(N__20561),
            .in2(N__20555),
            .in3(N__20533),
            .lcout(this_sprites_ram_mem_N_95),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_18_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_18_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_18_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_18_0  (
            .in0(N__21324),
            .in1(N__21060),
            .in2(N__21175),
            .in3(N__21249),
            .lcout(\this_sprites_ram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_21_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_21_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_21_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_21_6  (
            .in0(N__21331),
            .in1(N__21050),
            .in2(N__21161),
            .in3(N__21247),
            .lcout(\this_sprites_ram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI9MQ11_2_LC_24_22_4.C_ON=1'b0;
    defparam M_this_state_q_RNI9MQ11_2_LC_24_22_4.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI9MQ11_2_LC_24_22_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 M_this_state_q_RNI9MQ11_2_LC_24_22_4 (
            .in0(_gnd_net_),
            .in1(N__20387),
            .in2(_gnd_net_),
            .in3(N__20291),
            .lcout(M_this_sprites_ram_write_data_0_sqmuxa),
            .ltout(M_this_sprites_ram_write_data_0_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_ibuf_RNIGSD53_0_LC_24_22_5.C_ON=1'b0;
    defparam port_data_ibuf_RNIGSD53_0_LC_24_22_5.SEQ_MODE=4'b0000;
    defparam port_data_ibuf_RNIGSD53_0_LC_24_22_5.LUT_INIT=16'b1100000011101010;
    LogicCell40 port_data_ibuf_RNIGSD53_0_LC_24_22_5 (
            .in0(N__20173),
            .in1(N__20118),
            .in2(N__20075),
            .in3(N__21488),
            .lcout(M_this_sprites_ram_write_data_0_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_ibuf_RNIM2E53_7_LC_24_22_7.C_ON=1'b0;
    defparam port_data_ibuf_RNIM2E53_7_LC_24_22_7.SEQ_MODE=4'b0000;
    defparam port_data_ibuf_RNIM2E53_7_LC_24_22_7.LUT_INIT=16'b1111001000100010;
    LogicCell40 port_data_ibuf_RNIM2E53_7_LC_24_22_7 (
            .in0(N__19978),
            .in1(N__21489),
            .in2(N__19940),
            .in3(N__21423),
            .lcout(M_this_sprites_ram_write_data_0_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_ibuf_RNIK0E53_2_LC_24_23_0.C_ON=1'b0;
    defparam port_data_ibuf_RNIK0E53_2_LC_24_23_0.SEQ_MODE=4'b0000;
    defparam port_data_ibuf_RNIK0E53_2_LC_24_23_0.LUT_INIT=16'b1111001000100010;
    LogicCell40 port_data_ibuf_RNIK0E53_2_LC_24_23_0 (
            .in0(N__19827),
            .in1(N__21491),
            .in2(N__19788),
            .in3(N__21425),
            .lcout(M_this_sprites_ram_write_data_0_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_ibuf_RNIIUD53_1_LC_24_23_4.C_ON=1'b0;
    defparam port_data_ibuf_RNIIUD53_1_LC_24_23_4.SEQ_MODE=4'b0000;
    defparam port_data_ibuf_RNIIUD53_1_LC_24_23_4.LUT_INIT=16'b1111001000100010;
    LogicCell40 port_data_ibuf_RNIIUD53_1_LC_24_23_4 (
            .in0(N__21531),
            .in1(N__21490),
            .in2(N__21465),
            .in3(N__21424),
            .lcout(M_this_sprites_ram_write_data_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_24_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_24_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_24_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_24_5  (
            .in0(N__21320),
            .in1(N__21248),
            .in2(N__21160),
            .in3(N__21030),
            .lcout(\this_sprites_ram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_0_LC_30_23_0.C_ON=1'b1;
    defparam M_this_external_address_q_0_LC_30_23_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_0_LC_30_23_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_0_LC_30_23_0 (
            .in0(N__22482),
            .in1(N__20824),
            .in2(N__20974),
            .in3(N__20969),
            .lcout(M_this_external_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_30_23_0_),
            .carryout(un1_M_this_external_address_q_cry_0),
            .clk(N__22239),
            .ce(),
            .sr(N__21945));
    defparam M_this_external_address_q_1_LC_30_23_1.C_ON=1'b1;
    defparam M_this_external_address_q_1_LC_30_23_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_1_LC_30_23_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_1_LC_30_23_1 (
            .in0(N__22488),
            .in1(N__20803),
            .in2(_gnd_net_),
            .in3(N__20792),
            .lcout(M_this_external_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_0),
            .carryout(un1_M_this_external_address_q_cry_1),
            .clk(N__22239),
            .ce(),
            .sr(N__21945));
    defparam M_this_external_address_q_2_LC_30_23_2.C_ON=1'b1;
    defparam M_this_external_address_q_2_LC_30_23_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_2_LC_30_23_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_2_LC_30_23_2 (
            .in0(N__22483),
            .in1(N__20773),
            .in2(_gnd_net_),
            .in3(N__20762),
            .lcout(M_this_external_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_1),
            .carryout(un1_M_this_external_address_q_cry_2),
            .clk(N__22239),
            .ce(),
            .sr(N__21945));
    defparam M_this_external_address_q_3_LC_30_23_3.C_ON=1'b1;
    defparam M_this_external_address_q_3_LC_30_23_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_3_LC_30_23_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_3_LC_30_23_3 (
            .in0(N__22489),
            .in1(N__20749),
            .in2(_gnd_net_),
            .in3(N__20738),
            .lcout(M_this_external_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_2),
            .carryout(un1_M_this_external_address_q_cry_3),
            .clk(N__22239),
            .ce(),
            .sr(N__21945));
    defparam M_this_external_address_q_4_LC_30_23_4.C_ON=1'b1;
    defparam M_this_external_address_q_4_LC_30_23_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_4_LC_30_23_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_4_LC_30_23_4 (
            .in0(N__22484),
            .in1(N__20731),
            .in2(_gnd_net_),
            .in3(N__20720),
            .lcout(M_this_external_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_3),
            .carryout(un1_M_this_external_address_q_cry_4),
            .clk(N__22239),
            .ce(),
            .sr(N__21945));
    defparam M_this_external_address_q_5_LC_30_23_5.C_ON=1'b1;
    defparam M_this_external_address_q_5_LC_30_23_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_5_LC_30_23_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_5_LC_30_23_5 (
            .in0(N__22486),
            .in1(N__20710),
            .in2(_gnd_net_),
            .in3(N__20699),
            .lcout(M_this_external_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_4),
            .carryout(un1_M_this_external_address_q_cry_5),
            .clk(N__22239),
            .ce(),
            .sr(N__21945));
    defparam M_this_external_address_q_6_LC_30_23_6.C_ON=1'b1;
    defparam M_this_external_address_q_6_LC_30_23_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_6_LC_30_23_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_6_LC_30_23_6 (
            .in0(N__22485),
            .in1(N__21727),
            .in2(_gnd_net_),
            .in3(N__21716),
            .lcout(M_this_external_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_5),
            .carryout(un1_M_this_external_address_q_cry_6),
            .clk(N__22239),
            .ce(),
            .sr(N__21945));
    defparam M_this_external_address_q_7_LC_30_23_7.C_ON=1'b1;
    defparam M_this_external_address_q_7_LC_30_23_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_7_LC_30_23_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_7_LC_30_23_7 (
            .in0(N__22487),
            .in1(N__21700),
            .in2(_gnd_net_),
            .in3(N__21689),
            .lcout(M_this_external_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_6),
            .carryout(un1_M_this_external_address_q_cry_7),
            .clk(N__22239),
            .ce(),
            .sr(N__21945));
    defparam M_this_external_address_q_8_LC_30_24_0.C_ON=1'b1;
    defparam M_this_external_address_q_8_LC_30_24_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_8_LC_30_24_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_8_LC_30_24_0 (
            .in0(N__22507),
            .in1(N__21667),
            .in2(_gnd_net_),
            .in3(N__21656),
            .lcout(M_this_external_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_30_24_0_),
            .carryout(un1_M_this_external_address_q_cry_8),
            .clk(N__22242),
            .ce(),
            .sr(N__21944));
    defparam M_this_external_address_q_9_LC_30_24_1.C_ON=1'b1;
    defparam M_this_external_address_q_9_LC_30_24_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_9_LC_30_24_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_9_LC_30_24_1 (
            .in0(N__22492),
            .in1(N__21646),
            .in2(_gnd_net_),
            .in3(N__21635),
            .lcout(M_this_external_address_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_8),
            .carryout(un1_M_this_external_address_q_cry_9),
            .clk(N__22242),
            .ce(),
            .sr(N__21944));
    defparam M_this_external_address_q_10_LC_30_24_2.C_ON=1'b1;
    defparam M_this_external_address_q_10_LC_30_24_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_10_LC_30_24_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_10_LC_30_24_2 (
            .in0(N__22504),
            .in1(N__21616),
            .in2(_gnd_net_),
            .in3(N__21605),
            .lcout(M_this_external_address_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_9),
            .carryout(un1_M_this_external_address_q_cry_10),
            .clk(N__22242),
            .ce(),
            .sr(N__21944));
    defparam M_this_external_address_q_11_LC_30_24_3.C_ON=1'b1;
    defparam M_this_external_address_q_11_LC_30_24_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_11_LC_30_24_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_11_LC_30_24_3 (
            .in0(N__22490),
            .in1(N__21598),
            .in2(_gnd_net_),
            .in3(N__21587),
            .lcout(M_this_external_address_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_10),
            .carryout(un1_M_this_external_address_q_cry_11),
            .clk(N__22242),
            .ce(),
            .sr(N__21944));
    defparam M_this_external_address_q_12_LC_30_24_4.C_ON=1'b1;
    defparam M_this_external_address_q_12_LC_30_24_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_12_LC_30_24_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_12_LC_30_24_4 (
            .in0(N__22505),
            .in1(N__21580),
            .in2(_gnd_net_),
            .in3(N__21569),
            .lcout(M_this_external_address_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_11),
            .carryout(un1_M_this_external_address_q_cry_12),
            .clk(N__22242),
            .ce(),
            .sr(N__21944));
    defparam M_this_external_address_q_13_LC_30_24_5.C_ON=1'b1;
    defparam M_this_external_address_q_13_LC_30_24_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_13_LC_30_24_5.LUT_INIT=16'b1011101111101110;
    LogicCell40 M_this_external_address_q_13_LC_30_24_5 (
            .in0(N__22491),
            .in1(N__21556),
            .in2(_gnd_net_),
            .in3(N__21545),
            .lcout(M_this_external_address_qZ0Z_13),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_12),
            .carryout(un1_M_this_external_address_q_cry_13),
            .clk(N__22242),
            .ce(),
            .sr(N__21944));
    defparam M_this_external_address_q_14_LC_30_24_6.C_ON=1'b1;
    defparam M_this_external_address_q_14_LC_30_24_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_14_LC_30_24_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_14_LC_30_24_6 (
            .in0(N__22506),
            .in1(N__22522),
            .in2(_gnd_net_),
            .in3(N__22511),
            .lcout(M_this_external_address_qZ0Z_14),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_13),
            .carryout(un1_M_this_external_address_q_cry_14),
            .clk(N__22242),
            .ce(),
            .sr(N__21944));
    defparam M_this_external_address_q_15_LC_30_24_7.C_ON=1'b0;
    defparam M_this_external_address_q_15_LC_30_24_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_15_LC_30_24_7.LUT_INIT=16'b1101110111101110;
    LogicCell40 M_this_external_address_q_15_LC_30_24_7 (
            .in0(N__22255),
            .in1(N__22508),
            .in2(_gnd_net_),
            .in3(N__22271),
            .lcout(M_this_external_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22242),
            .ce(),
            .sr(N__21944));
    defparam port_address_iobuf_RNI6NG6_2_LC_32_22_1.C_ON=1'b0;
    defparam port_address_iobuf_RNI6NG6_2_LC_32_22_1.SEQ_MODE=4'b0000;
    defparam port_address_iobuf_RNI6NG6_2_LC_32_22_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 port_address_iobuf_RNI6NG6_2_LC_32_22_1 (
            .in0(N__21857),
            .in1(N__21845),
            .in2(N__21839),
            .in3(N__21830),
            .lcout(),
            .ltout(M_this_state_d36_2_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_address_iobuf_RNIV8P9_6_LC_32_22_2.C_ON=1'b0;
    defparam port_address_iobuf_RNIV8P9_6_LC_32_22_2.SEQ_MODE=4'b0000;
    defparam port_address_iobuf_RNIV8P9_6_LC_32_22_2.LUT_INIT=16'b0000000001010000;
    LogicCell40 port_address_iobuf_RNIV8P9_6_LC_32_22_2 (
            .in0(N__21806),
            .in1(_gnd_net_),
            .in2(N__21782),
            .in3(N__21779),
            .lcout(M_this_state_d37_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
