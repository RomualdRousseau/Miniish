// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 28 2022 16:04:31

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    led,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    input [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output [7:0] led;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__36351;
    wire N__36350;
    wire N__36349;
    wire N__36340;
    wire N__36339;
    wire N__36338;
    wire N__36331;
    wire N__36330;
    wire N__36329;
    wire N__36322;
    wire N__36321;
    wire N__36320;
    wire N__36313;
    wire N__36312;
    wire N__36311;
    wire N__36304;
    wire N__36303;
    wire N__36302;
    wire N__36295;
    wire N__36294;
    wire N__36293;
    wire N__36286;
    wire N__36285;
    wire N__36284;
    wire N__36277;
    wire N__36276;
    wire N__36275;
    wire N__36268;
    wire N__36267;
    wire N__36266;
    wire N__36259;
    wire N__36258;
    wire N__36257;
    wire N__36250;
    wire N__36249;
    wire N__36248;
    wire N__36241;
    wire N__36240;
    wire N__36239;
    wire N__36232;
    wire N__36231;
    wire N__36230;
    wire N__36223;
    wire N__36222;
    wire N__36221;
    wire N__36214;
    wire N__36213;
    wire N__36212;
    wire N__36205;
    wire N__36204;
    wire N__36203;
    wire N__36196;
    wire N__36195;
    wire N__36194;
    wire N__36187;
    wire N__36186;
    wire N__36185;
    wire N__36178;
    wire N__36177;
    wire N__36176;
    wire N__36169;
    wire N__36168;
    wire N__36167;
    wire N__36160;
    wire N__36159;
    wire N__36158;
    wire N__36151;
    wire N__36150;
    wire N__36149;
    wire N__36142;
    wire N__36141;
    wire N__36140;
    wire N__36133;
    wire N__36132;
    wire N__36131;
    wire N__36124;
    wire N__36123;
    wire N__36122;
    wire N__36115;
    wire N__36114;
    wire N__36113;
    wire N__36106;
    wire N__36105;
    wire N__36104;
    wire N__36097;
    wire N__36096;
    wire N__36095;
    wire N__36088;
    wire N__36087;
    wire N__36086;
    wire N__36079;
    wire N__36078;
    wire N__36077;
    wire N__36070;
    wire N__36069;
    wire N__36068;
    wire N__36061;
    wire N__36060;
    wire N__36059;
    wire N__36052;
    wire N__36051;
    wire N__36050;
    wire N__36043;
    wire N__36042;
    wire N__36041;
    wire N__36034;
    wire N__36033;
    wire N__36032;
    wire N__36025;
    wire N__36024;
    wire N__36023;
    wire N__36016;
    wire N__36015;
    wire N__36014;
    wire N__36007;
    wire N__36006;
    wire N__36005;
    wire N__35998;
    wire N__35997;
    wire N__35996;
    wire N__35989;
    wire N__35988;
    wire N__35987;
    wire N__35980;
    wire N__35979;
    wire N__35978;
    wire N__35971;
    wire N__35970;
    wire N__35969;
    wire N__35962;
    wire N__35961;
    wire N__35960;
    wire N__35953;
    wire N__35952;
    wire N__35951;
    wire N__35944;
    wire N__35943;
    wire N__35942;
    wire N__35935;
    wire N__35934;
    wire N__35933;
    wire N__35926;
    wire N__35925;
    wire N__35924;
    wire N__35917;
    wire N__35916;
    wire N__35915;
    wire N__35908;
    wire N__35907;
    wire N__35906;
    wire N__35899;
    wire N__35898;
    wire N__35897;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35871;
    wire N__35868;
    wire N__35867;
    wire N__35866;
    wire N__35865;
    wire N__35864;
    wire N__35863;
    wire N__35862;
    wire N__35861;
    wire N__35860;
    wire N__35859;
    wire N__35858;
    wire N__35857;
    wire N__35856;
    wire N__35855;
    wire N__35854;
    wire N__35853;
    wire N__35852;
    wire N__35851;
    wire N__35850;
    wire N__35847;
    wire N__35846;
    wire N__35829;
    wire N__35814;
    wire N__35813;
    wire N__35812;
    wire N__35811;
    wire N__35810;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35793;
    wire N__35788;
    wire N__35787;
    wire N__35786;
    wire N__35785;
    wire N__35784;
    wire N__35783;
    wire N__35782;
    wire N__35781;
    wire N__35780;
    wire N__35779;
    wire N__35778;
    wire N__35775;
    wire N__35766;
    wire N__35765;
    wire N__35764;
    wire N__35763;
    wire N__35756;
    wire N__35755;
    wire N__35750;
    wire N__35747;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35718;
    wire N__35717;
    wire N__35716;
    wire N__35715;
    wire N__35714;
    wire N__35713;
    wire N__35708;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35680;
    wire N__35673;
    wire N__35666;
    wire N__35661;
    wire N__35640;
    wire N__35639;
    wire N__35638;
    wire N__35637;
    wire N__35636;
    wire N__35635;
    wire N__35634;
    wire N__35619;
    wire N__35618;
    wire N__35617;
    wire N__35616;
    wire N__35615;
    wire N__35614;
    wire N__35613;
    wire N__35612;
    wire N__35611;
    wire N__35610;
    wire N__35609;
    wire N__35606;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35580;
    wire N__35579;
    wire N__35578;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35538;
    wire N__35535;
    wire N__35532;
    wire N__35529;
    wire N__35526;
    wire N__35523;
    wire N__35520;
    wire N__35519;
    wire N__35516;
    wire N__35515;
    wire N__35512;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35487;
    wire N__35486;
    wire N__35485;
    wire N__35484;
    wire N__35483;
    wire N__35482;
    wire N__35481;
    wire N__35480;
    wire N__35479;
    wire N__35470;
    wire N__35469;
    wire N__35468;
    wire N__35467;
    wire N__35466;
    wire N__35463;
    wire N__35460;
    wire N__35453;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35445;
    wire N__35444;
    wire N__35443;
    wire N__35442;
    wire N__35441;
    wire N__35440;
    wire N__35439;
    wire N__35436;
    wire N__35435;
    wire N__35432;
    wire N__35431;
    wire N__35430;
    wire N__35429;
    wire N__35428;
    wire N__35427;
    wire N__35424;
    wire N__35423;
    wire N__35422;
    wire N__35421;
    wire N__35420;
    wire N__35419;
    wire N__35418;
    wire N__35415;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35400;
    wire N__35399;
    wire N__35398;
    wire N__35397;
    wire N__35392;
    wire N__35383;
    wire N__35380;
    wire N__35377;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35359;
    wire N__35356;
    wire N__35345;
    wire N__35342;
    wire N__35341;
    wire N__35340;
    wire N__35337;
    wire N__35334;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35316;
    wire N__35313;
    wire N__35306;
    wire N__35303;
    wire N__35292;
    wire N__35289;
    wire N__35284;
    wire N__35279;
    wire N__35274;
    wire N__35261;
    wire N__35250;
    wire N__35249;
    wire N__35248;
    wire N__35247;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35239;
    wire N__35238;
    wire N__35237;
    wire N__35236;
    wire N__35235;
    wire N__35234;
    wire N__35233;
    wire N__35232;
    wire N__35231;
    wire N__35230;
    wire N__35229;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35213;
    wire N__35210;
    wire N__35201;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35190;
    wire N__35189;
    wire N__35188;
    wire N__35187;
    wire N__35186;
    wire N__35185;
    wire N__35184;
    wire N__35183;
    wire N__35180;
    wire N__35177;
    wire N__35176;
    wire N__35175;
    wire N__35174;
    wire N__35171;
    wire N__35170;
    wire N__35169;
    wire N__35166;
    wire N__35165;
    wire N__35164;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35129;
    wire N__35126;
    wire N__35123;
    wire N__35122;
    wire N__35121;
    wire N__35120;
    wire N__35119;
    wire N__35116;
    wire N__35111;
    wire N__35106;
    wire N__35099;
    wire N__35098;
    wire N__35095;
    wire N__35090;
    wire N__35081;
    wire N__35080;
    wire N__35071;
    wire N__35064;
    wire N__35061;
    wire N__35058;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35027;
    wire N__35020;
    wire N__35015;
    wire N__35004;
    wire N__35003;
    wire N__35002;
    wire N__35001;
    wire N__35000;
    wire N__34999;
    wire N__34998;
    wire N__34997;
    wire N__34996;
    wire N__34995;
    wire N__34994;
    wire N__34991;
    wire N__34990;
    wire N__34989;
    wire N__34988;
    wire N__34987;
    wire N__34986;
    wire N__34983;
    wire N__34982;
    wire N__34981;
    wire N__34980;
    wire N__34979;
    wire N__34978;
    wire N__34975;
    wire N__34966;
    wire N__34963;
    wire N__34962;
    wire N__34959;
    wire N__34954;
    wire N__34953;
    wire N__34952;
    wire N__34951;
    wire N__34950;
    wire N__34947;
    wire N__34940;
    wire N__34939;
    wire N__34938;
    wire N__34937;
    wire N__34936;
    wire N__34935;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34923;
    wire N__34922;
    wire N__34921;
    wire N__34920;
    wire N__34911;
    wire N__34908;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34894;
    wire N__34893;
    wire N__34892;
    wire N__34891;
    wire N__34890;
    wire N__34889;
    wire N__34882;
    wire N__34879;
    wire N__34874;
    wire N__34867;
    wire N__34862;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34843;
    wire N__34836;
    wire N__34833;
    wire N__34828;
    wire N__34817;
    wire N__34814;
    wire N__34803;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34766;
    wire N__34763;
    wire N__34762;
    wire N__34761;
    wire N__34758;
    wire N__34757;
    wire N__34754;
    wire N__34751;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34741;
    wire N__34740;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34707;
    wire N__34706;
    wire N__34705;
    wire N__34702;
    wire N__34699;
    wire N__34696;
    wire N__34695;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34684;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34665;
    wire N__34664;
    wire N__34659;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34635;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34612;
    wire N__34605;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34595;
    wire N__34594;
    wire N__34593;
    wire N__34592;
    wire N__34591;
    wire N__34590;
    wire N__34589;
    wire N__34588;
    wire N__34587;
    wire N__34586;
    wire N__34585;
    wire N__34584;
    wire N__34583;
    wire N__34582;
    wire N__34581;
    wire N__34580;
    wire N__34579;
    wire N__34578;
    wire N__34577;
    wire N__34576;
    wire N__34575;
    wire N__34574;
    wire N__34573;
    wire N__34572;
    wire N__34571;
    wire N__34570;
    wire N__34569;
    wire N__34568;
    wire N__34567;
    wire N__34566;
    wire N__34565;
    wire N__34564;
    wire N__34563;
    wire N__34562;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34557;
    wire N__34556;
    wire N__34555;
    wire N__34554;
    wire N__34553;
    wire N__34552;
    wire N__34551;
    wire N__34550;
    wire N__34549;
    wire N__34548;
    wire N__34547;
    wire N__34546;
    wire N__34545;
    wire N__34544;
    wire N__34543;
    wire N__34542;
    wire N__34541;
    wire N__34540;
    wire N__34539;
    wire N__34538;
    wire N__34537;
    wire N__34536;
    wire N__34535;
    wire N__34534;
    wire N__34533;
    wire N__34532;
    wire N__34531;
    wire N__34530;
    wire N__34529;
    wire N__34528;
    wire N__34527;
    wire N__34526;
    wire N__34525;
    wire N__34524;
    wire N__34523;
    wire N__34522;
    wire N__34521;
    wire N__34520;
    wire N__34519;
    wire N__34518;
    wire N__34517;
    wire N__34516;
    wire N__34515;
    wire N__34514;
    wire N__34513;
    wire N__34512;
    wire N__34511;
    wire N__34510;
    wire N__34509;
    wire N__34508;
    wire N__34507;
    wire N__34506;
    wire N__34505;
    wire N__34504;
    wire N__34503;
    wire N__34502;
    wire N__34501;
    wire N__34500;
    wire N__34499;
    wire N__34498;
    wire N__34497;
    wire N__34496;
    wire N__34495;
    wire N__34494;
    wire N__34493;
    wire N__34492;
    wire N__34491;
    wire N__34490;
    wire N__34489;
    wire N__34488;
    wire N__34487;
    wire N__34486;
    wire N__34485;
    wire N__34484;
    wire N__34483;
    wire N__34482;
    wire N__34481;
    wire N__34480;
    wire N__34479;
    wire N__34478;
    wire N__34477;
    wire N__34476;
    wire N__34475;
    wire N__34474;
    wire N__34473;
    wire N__34472;
    wire N__34471;
    wire N__34470;
    wire N__34469;
    wire N__34468;
    wire N__34467;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34199;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34188;
    wire N__34187;
    wire N__34184;
    wire N__34179;
    wire N__34176;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34164;
    wire N__34163;
    wire N__34162;
    wire N__34159;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34138;
    wire N__34135;
    wire N__34130;
    wire N__34125;
    wire N__34124;
    wire N__34123;
    wire N__34122;
    wire N__34121;
    wire N__34120;
    wire N__34119;
    wire N__34118;
    wire N__34117;
    wire N__34116;
    wire N__34115;
    wire N__34114;
    wire N__34113;
    wire N__34112;
    wire N__34111;
    wire N__34110;
    wire N__34109;
    wire N__34108;
    wire N__34107;
    wire N__34106;
    wire N__34105;
    wire N__34104;
    wire N__34101;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34041;
    wire N__34040;
    wire N__34039;
    wire N__34038;
    wire N__34037;
    wire N__34036;
    wire N__34035;
    wire N__34034;
    wire N__34033;
    wire N__34032;
    wire N__34031;
    wire N__34030;
    wire N__34029;
    wire N__34028;
    wire N__34027;
    wire N__34026;
    wire N__34025;
    wire N__34024;
    wire N__34023;
    wire N__34022;
    wire N__34021;
    wire N__34020;
    wire N__34019;
    wire N__34018;
    wire N__34017;
    wire N__34016;
    wire N__34015;
    wire N__34014;
    wire N__34013;
    wire N__34012;
    wire N__34011;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33995;
    wire N__33992;
    wire N__33989;
    wire N__33986;
    wire N__33983;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33953;
    wire N__33852;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33826;
    wire N__33825;
    wire N__33822;
    wire N__33819;
    wire N__33818;
    wire N__33815;
    wire N__33814;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33801;
    wire N__33800;
    wire N__33799;
    wire N__33796;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33757;
    wire N__33754;
    wire N__33751;
    wire N__33750;
    wire N__33745;
    wire N__33742;
    wire N__33739;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33717;
    wire N__33714;
    wire N__33711;
    wire N__33708;
    wire N__33705;
    wire N__33696;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33672;
    wire N__33671;
    wire N__33670;
    wire N__33669;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33658;
    wire N__33657;
    wire N__33654;
    wire N__33651;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33630;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33589;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33546;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33524;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33506;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33491;
    wire N__33488;
    wire N__33487;
    wire N__33484;
    wire N__33483;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33472;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33458;
    wire N__33455;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33444;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33434;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33422;
    wire N__33421;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33383;
    wire N__33380;
    wire N__33375;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33360;
    wire N__33357;
    wire N__33348;
    wire N__33345;
    wire N__33342;
    wire N__33337;
    wire N__33330;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33318;
    wire N__33317;
    wire N__33314;
    wire N__33311;
    wire N__33306;
    wire N__33303;
    wire N__33300;
    wire N__33297;
    wire N__33296;
    wire N__33293;
    wire N__33290;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33262;
    wire N__33259;
    wire N__33256;
    wire N__33253;
    wire N__33250;
    wire N__33247;
    wire N__33244;
    wire N__33241;
    wire N__33234;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33222;
    wire N__33221;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33174;
    wire N__33173;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33149;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33129;
    wire N__33126;
    wire N__33125;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33101;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33084;
    wire N__33083;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33039;
    wire N__33038;
    wire N__33035;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32987;
    wire N__32986;
    wire N__32985;
    wire N__32982;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32955;
    wire N__32954;
    wire N__32951;
    wire N__32946;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32930;
    wire N__32927;
    wire N__32926;
    wire N__32923;
    wire N__32918;
    wire N__32917;
    wire N__32916;
    wire N__32913;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32878;
    wire N__32873;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32856;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32834;
    wire N__32833;
    wire N__32832;
    wire N__32831;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32802;
    wire N__32801;
    wire N__32800;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32782;
    wire N__32779;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32759;
    wire N__32756;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32731;
    wire N__32728;
    wire N__32725;
    wire N__32720;
    wire N__32717;
    wire N__32714;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32700;
    wire N__32691;
    wire N__32688;
    wire N__32685;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32643;
    wire N__32640;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32617;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32598;
    wire N__32595;
    wire N__32594;
    wire N__32593;
    wire N__32592;
    wire N__32589;
    wire N__32588;
    wire N__32585;
    wire N__32582;
    wire N__32579;
    wire N__32578;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32568;
    wire N__32565;
    wire N__32562;
    wire N__32559;
    wire N__32556;
    wire N__32551;
    wire N__32548;
    wire N__32547;
    wire N__32544;
    wire N__32543;
    wire N__32538;
    wire N__32533;
    wire N__32530;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32502;
    wire N__32499;
    wire N__32494;
    wire N__32489;
    wire N__32486;
    wire N__32481;
    wire N__32480;
    wire N__32477;
    wire N__32474;
    wire N__32471;
    wire N__32468;
    wire N__32465;
    wire N__32462;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32408;
    wire N__32407;
    wire N__32404;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32393;
    wire N__32390;
    wire N__32389;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32365;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32353;
    wire N__32352;
    wire N__32349;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32335;
    wire N__32332;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32305;
    wire N__32302;
    wire N__32299;
    wire N__32290;
    wire N__32287;
    wire N__32282;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32190;
    wire N__32189;
    wire N__32188;
    wire N__32185;
    wire N__32184;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32143;
    wire N__32140;
    wire N__32137;
    wire N__32134;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31988;
    wire N__31985;
    wire N__31984;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31974;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31968;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31948;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31940;
    wire N__31937;
    wire N__31932;
    wire N__31929;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31890;
    wire N__31887;
    wire N__31886;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31875;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31863;
    wire N__31862;
    wire N__31861;
    wire N__31858;
    wire N__31853;
    wire N__31850;
    wire N__31847;
    wire N__31846;
    wire N__31845;
    wire N__31844;
    wire N__31843;
    wire N__31840;
    wire N__31835;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31800;
    wire N__31799;
    wire N__31796;
    wire N__31795;
    wire N__31792;
    wire N__31791;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31783;
    wire N__31780;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31754;
    wire N__31753;
    wire N__31750;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31724;
    wire N__31721;
    wire N__31718;
    wire N__31711;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31699;
    wire N__31696;
    wire N__31693;
    wire N__31686;
    wire N__31671;
    wire N__31668;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31660;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31649;
    wire N__31646;
    wire N__31645;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31627;
    wire N__31626;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31593;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31541;
    wire N__31540;
    wire N__31537;
    wire N__31536;
    wire N__31535;
    wire N__31534;
    wire N__31529;
    wire N__31526;
    wire N__31519;
    wire N__31516;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31438;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31416;
    wire N__31415;
    wire N__31412;
    wire N__31409;
    wire N__31406;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31373;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31282;
    wire N__31279;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31257;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31249;
    wire N__31248;
    wire N__31247;
    wire N__31244;
    wire N__31239;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31205;
    wire N__31202;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31180;
    wire N__31177;
    wire N__31172;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31127;
    wire N__31124;
    wire N__31121;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31094;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30929;
    wire N__30928;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30916;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30879;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30871;
    wire N__30870;
    wire N__30865;
    wire N__30862;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30830;
    wire N__30827;
    wire N__30824;
    wire N__30819;
    wire N__30816;
    wire N__30815;
    wire N__30812;
    wire N__30811;
    wire N__30808;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30789;
    wire N__30786;
    wire N__30783;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30775;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30690;
    wire N__30689;
    wire N__30686;
    wire N__30685;
    wire N__30684;
    wire N__30683;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30639;
    wire N__30636;
    wire N__30635;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30622;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30602;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30590;
    wire N__30587;
    wire N__30586;
    wire N__30585;
    wire N__30582;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30569;
    wire N__30566;
    wire N__30563;
    wire N__30552;
    wire N__30551;
    wire N__30550;
    wire N__30547;
    wire N__30542;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30507;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30465;
    wire N__30464;
    wire N__30461;
    wire N__30460;
    wire N__30459;
    wire N__30458;
    wire N__30457;
    wire N__30456;
    wire N__30455;
    wire N__30454;
    wire N__30453;
    wire N__30450;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30431;
    wire N__30426;
    wire N__30425;
    wire N__30424;
    wire N__30423;
    wire N__30420;
    wire N__30419;
    wire N__30418;
    wire N__30415;
    wire N__30404;
    wire N__30397;
    wire N__30394;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30357;
    wire N__30356;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30318;
    wire N__30315;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30300;
    wire N__30297;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30282;
    wire N__30279;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30264;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30181;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30165;
    wire N__30164;
    wire N__30163;
    wire N__30162;
    wire N__30161;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30153;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30145;
    wire N__30142;
    wire N__30137;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30113;
    wire N__30112;
    wire N__30109;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30083;
    wire N__30082;
    wire N__30081;
    wire N__30078;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30064;
    wire N__30059;
    wire N__30056;
    wire N__30055;
    wire N__30052;
    wire N__30045;
    wire N__30038;
    wire N__30033;
    wire N__30024;
    wire N__30021;
    wire N__30020;
    wire N__30019;
    wire N__30018;
    wire N__30017;
    wire N__30016;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30006;
    wire N__30003;
    wire N__30002;
    wire N__30001;
    wire N__30000;
    wire N__29999;
    wire N__29998;
    wire N__29997;
    wire N__29992;
    wire N__29991;
    wire N__29990;
    wire N__29987;
    wire N__29982;
    wire N__29979;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29942;
    wire N__29941;
    wire N__29938;
    wire N__29931;
    wire N__29928;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29910;
    wire N__29907;
    wire N__29904;
    wire N__29899;
    wire N__29896;
    wire N__29883;
    wire N__29882;
    wire N__29879;
    wire N__29876;
    wire N__29875;
    wire N__29874;
    wire N__29871;
    wire N__29870;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29862;
    wire N__29859;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29851;
    wire N__29848;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29822;
    wire N__29819;
    wire N__29816;
    wire N__29815;
    wire N__29814;
    wire N__29809;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29798;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29759;
    wire N__29756;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29678;
    wire N__29675;
    wire N__29670;
    wire N__29665;
    wire N__29662;
    wire N__29657;
    wire N__29650;
    wire N__29641;
    wire N__29634;
    wire N__29633;
    wire N__29632;
    wire N__29631;
    wire N__29630;
    wire N__29629;
    wire N__29628;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29601;
    wire N__29600;
    wire N__29595;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29564;
    wire N__29561;
    wire N__29558;
    wire N__29557;
    wire N__29556;
    wire N__29555;
    wire N__29552;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29507;
    wire N__29506;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29474;
    wire N__29473;
    wire N__29472;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29460;
    wire N__29457;
    wire N__29456;
    wire N__29451;
    wire N__29448;
    wire N__29443;
    wire N__29436;
    wire N__29435;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29413;
    wire N__29410;
    wire N__29407;
    wire N__29404;
    wire N__29403;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29388;
    wire N__29379;
    wire N__29376;
    wire N__29373;
    wire N__29372;
    wire N__29371;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29359;
    wire N__29358;
    wire N__29357;
    wire N__29352;
    wire N__29349;
    wire N__29344;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29327;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29306;
    wire N__29305;
    wire N__29304;
    wire N__29303;
    wire N__29302;
    wire N__29299;
    wire N__29296;
    wire N__29291;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29265;
    wire N__29264;
    wire N__29261;
    wire N__29258;
    wire N__29255;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29199;
    wire N__29198;
    wire N__29197;
    wire N__29194;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29158;
    wire N__29155;
    wire N__29148;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29133;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29118;
    wire N__29117;
    wire N__29116;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29076;
    wire N__29073;
    wire N__29070;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29058;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29003;
    wire N__29000;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28989;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28977;
    wire N__28974;
    wire N__28967;
    wire N__28964;
    wire N__28961;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28949;
    wire N__28948;
    wire N__28945;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28920;
    wire N__28919;
    wire N__28918;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28889;
    wire N__28888;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28878;
    wire N__28875;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28851;
    wire N__28850;
    wire N__28845;
    wire N__28842;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28830;
    wire N__28827;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28791;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28739;
    wire N__28736;
    wire N__28731;
    wire N__28722;
    wire N__28721;
    wire N__28720;
    wire N__28717;
    wire N__28716;
    wire N__28715;
    wire N__28712;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28694;
    wire N__28689;
    wire N__28686;
    wire N__28677;
    wire N__28676;
    wire N__28673;
    wire N__28672;
    wire N__28669;
    wire N__28668;
    wire N__28665;
    wire N__28664;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28646;
    wire N__28643;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28617;
    wire N__28614;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28583;
    wire N__28580;
    wire N__28579;
    wire N__28576;
    wire N__28571;
    wire N__28568;
    wire N__28567;
    wire N__28562;
    wire N__28561;
    wire N__28558;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28534;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28520;
    wire N__28519;
    wire N__28516;
    wire N__28511;
    wire N__28506;
    wire N__28503;
    wire N__28502;
    wire N__28501;
    wire N__28500;
    wire N__28495;
    wire N__28490;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28478;
    wire N__28475;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28454;
    wire N__28451;
    wire N__28450;
    wire N__28447;
    wire N__28442;
    wire N__28441;
    wire N__28436;
    wire N__28433;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28415;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28407;
    wire N__28404;
    wire N__28399;
    wire N__28396;
    wire N__28395;
    wire N__28394;
    wire N__28391;
    wire N__28386;
    wire N__28383;
    wire N__28382;
    wire N__28379;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28364;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28284;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28269;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28257;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28245;
    wire N__28242;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28191;
    wire N__28188;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28133;
    wire N__28130;
    wire N__28127;
    wire N__28126;
    wire N__28121;
    wire N__28120;
    wire N__28119;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28109;
    wire N__28106;
    wire N__28103;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28032;
    wire N__28031;
    wire N__28030;
    wire N__28027;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28007;
    wire N__28004;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27992;
    wire N__27989;
    wire N__27986;
    wire N__27981;
    wire N__27980;
    wire N__27977;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27962;
    wire N__27959;
    wire N__27954;
    wire N__27951;
    wire N__27948;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27936;
    wire N__27933;
    wire N__27932;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27913;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27897;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27882;
    wire N__27881;
    wire N__27880;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27864;
    wire N__27861;
    wire N__27858;
    wire N__27857;
    wire N__27854;
    wire N__27853;
    wire N__27852;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27809;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27764;
    wire N__27761;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27728;
    wire N__27727;
    wire N__27726;
    wire N__27725;
    wire N__27724;
    wire N__27723;
    wire N__27722;
    wire N__27721;
    wire N__27716;
    wire N__27707;
    wire N__27704;
    wire N__27703;
    wire N__27702;
    wire N__27697;
    wire N__27692;
    wire N__27689;
    wire N__27686;
    wire N__27685;
    wire N__27684;
    wire N__27683;
    wire N__27680;
    wire N__27677;
    wire N__27670;
    wire N__27663;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27612;
    wire N__27611;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27599;
    wire N__27596;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27584;
    wire N__27581;
    wire N__27580;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27561;
    wire N__27556;
    wire N__27553;
    wire N__27550;
    wire N__27549;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27538;
    wire N__27533;
    wire N__27530;
    wire N__27529;
    wire N__27526;
    wire N__27523;
    wire N__27522;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27493;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27466;
    wire N__27461;
    wire N__27456;
    wire N__27449;
    wire N__27446;
    wire N__27445;
    wire N__27442;
    wire N__27441;
    wire N__27438;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27415;
    wire N__27412;
    wire N__27405;
    wire N__27404;
    wire N__27401;
    wire N__27400;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27379;
    wire N__27376;
    wire N__27369;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27361;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27321;
    wire N__27318;
    wire N__27317;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27309;
    wire N__27306;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27295;
    wire N__27292;
    wire N__27289;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27273;
    wire N__27268;
    wire N__27265;
    wire N__27264;
    wire N__27263;
    wire N__27260;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27227;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27203;
    wire N__27202;
    wire N__27201;
    wire N__27200;
    wire N__27197;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27165;
    wire N__27164;
    wire N__27161;
    wire N__27158;
    wire N__27155;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27131;
    wire N__27128;
    wire N__27123;
    wire N__27120;
    wire N__27119;
    wire N__27116;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27084;
    wire N__27081;
    wire N__27080;
    wire N__27077;
    wire N__27072;
    wire N__27069;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27013;
    wire N__27006;
    wire N__26997;
    wire N__26996;
    wire N__26993;
    wire N__26992;
    wire N__26991;
    wire N__26990;
    wire N__26987;
    wire N__26986;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26978;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26947;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26897;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26863;
    wire N__26860;
    wire N__26859;
    wire N__26856;
    wire N__26851;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26831;
    wire N__26826;
    wire N__26823;
    wire N__26818;
    wire N__26813;
    wire N__26810;
    wire N__26803;
    wire N__26798;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26735;
    wire N__26732;
    wire N__26731;
    wire N__26728;
    wire N__26727;
    wire N__26726;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26709;
    wire N__26708;
    wire N__26703;
    wire N__26698;
    wire N__26695;
    wire N__26690;
    wire N__26687;
    wire N__26682;
    wire N__26681;
    wire N__26678;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26666;
    wire N__26663;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26609;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26598;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26584;
    wire N__26581;
    wire N__26580;
    wire N__26579;
    wire N__26578;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26563;
    wire N__26562;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26528;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26491;
    wire N__26486;
    wire N__26481;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26453;
    wire N__26448;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26434;
    wire N__26433;
    wire N__26430;
    wire N__26427;
    wire N__26420;
    wire N__26419;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26385;
    wire N__26384;
    wire N__26383;
    wire N__26380;
    wire N__26379;
    wire N__26378;
    wire N__26377;
    wire N__26376;
    wire N__26375;
    wire N__26374;
    wire N__26373;
    wire N__26370;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26358;
    wire N__26357;
    wire N__26356;
    wire N__26353;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26335;
    wire N__26330;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26318;
    wire N__26315;
    wire N__26310;
    wire N__26307;
    wire N__26298;
    wire N__26293;
    wire N__26292;
    wire N__26291;
    wire N__26290;
    wire N__26287;
    wire N__26284;
    wire N__26281;
    wire N__26276;
    wire N__26273;
    wire N__26268;
    wire N__26265;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26215;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26201;
    wire N__26200;
    wire N__26199;
    wire N__26198;
    wire N__26197;
    wire N__26196;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26178;
    wire N__26177;
    wire N__26176;
    wire N__26173;
    wire N__26170;
    wire N__26167;
    wire N__26164;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26148;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26140;
    wire N__26139;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26104;
    wire N__26101;
    wire N__26098;
    wire N__26097;
    wire N__26090;
    wire N__26087;
    wire N__26082;
    wire N__26079;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26057;
    wire N__26052;
    wire N__26045;
    wire N__26044;
    wire N__26039;
    wire N__26036;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26016;
    wire N__26013;
    wire N__26012;
    wire N__26011;
    wire N__26010;
    wire N__26007;
    wire N__26000;
    wire N__25995;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25952;
    wire N__25951;
    wire N__25948;
    wire N__25947;
    wire N__25944;
    wire N__25937;
    wire N__25932;
    wire N__25931;
    wire N__25930;
    wire N__25927;
    wire N__25926;
    wire N__25925;
    wire N__25922;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25911;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25896;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25866;
    wire N__25857;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25808;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25800;
    wire N__25799;
    wire N__25798;
    wire N__25795;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25784;
    wire N__25781;
    wire N__25780;
    wire N__25777;
    wire N__25776;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25741;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25678;
    wire N__25675;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25632;
    wire N__25627;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25597;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25573;
    wire N__25572;
    wire N__25571;
    wire N__25570;
    wire N__25569;
    wire N__25568;
    wire N__25567;
    wire N__25564;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25520;
    wire N__25519;
    wire N__25518;
    wire N__25517;
    wire N__25514;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25502;
    wire N__25501;
    wire N__25498;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25469;
    wire N__25468;
    wire N__25465;
    wire N__25464;
    wire N__25463;
    wire N__25462;
    wire N__25461;
    wire N__25460;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25384;
    wire N__25383;
    wire N__25382;
    wire N__25381;
    wire N__25378;
    wire N__25375;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25302;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25281;
    wire N__25272;
    wire N__25269;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25258;
    wire N__25257;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25243;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25227;
    wire N__25222;
    wire N__25219;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25185;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25170;
    wire N__25165;
    wire N__25162;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25139;
    wire N__25136;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25013;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25005;
    wire N__25004;
    wire N__25003;
    wire N__25002;
    wire N__24999;
    wire N__24998;
    wire N__24997;
    wire N__24996;
    wire N__24995;
    wire N__24990;
    wire N__24987;
    wire N__24986;
    wire N__24985;
    wire N__24984;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24966;
    wire N__24965;
    wire N__24962;
    wire N__24961;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24949;
    wire N__24946;
    wire N__24937;
    wire N__24934;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24919;
    wire N__24916;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24875;
    wire N__24874;
    wire N__24871;
    wire N__24868;
    wire N__24865;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24851;
    wire N__24850;
    wire N__24849;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24831;
    wire N__24830;
    wire N__24827;
    wire N__24826;
    wire N__24825;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24811;
    wire N__24808;
    wire N__24807;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24793;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24740;
    wire N__24737;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24721;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24694;
    wire N__24691;
    wire N__24690;
    wire N__24689;
    wire N__24688;
    wire N__24683;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24599;
    wire N__24596;
    wire N__24595;
    wire N__24594;
    wire N__24593;
    wire N__24590;
    wire N__24589;
    wire N__24588;
    wire N__24587;
    wire N__24582;
    wire N__24577;
    wire N__24574;
    wire N__24569;
    wire N__24566;
    wire N__24561;
    wire N__24554;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24451;
    wire N__24450;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24433;
    wire N__24432;
    wire N__24431;
    wire N__24430;
    wire N__24429;
    wire N__24428;
    wire N__24427;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24404;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24390;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24345;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24333;
    wire N__24332;
    wire N__24325;
    wire N__24322;
    wire N__24319;
    wire N__24316;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24282;
    wire N__24281;
    wire N__24278;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24204;
    wire N__24201;
    wire N__24200;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24183;
    wire N__24182;
    wire N__24179;
    wire N__24178;
    wire N__24177;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24166;
    wire N__24165;
    wire N__24164;
    wire N__24163;
    wire N__24160;
    wire N__24159;
    wire N__24156;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24133;
    wire N__24132;
    wire N__24131;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24067;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24042;
    wire N__24039;
    wire N__24038;
    wire N__24035;
    wire N__24030;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23999;
    wire N__23996;
    wire N__23989;
    wire N__23986;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23951;
    wire N__23940;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23906;
    wire N__23905;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23893;
    wire N__23886;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23864;
    wire N__23863;
    wire N__23862;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23848;
    wire N__23845;
    wire N__23838;
    wire N__23835;
    wire N__23832;
    wire N__23829;
    wire N__23826;
    wire N__23825;
    wire N__23822;
    wire N__23821;
    wire N__23820;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23805;
    wire N__23802;
    wire N__23799;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23768;
    wire N__23767;
    wire N__23764;
    wire N__23763;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23730;
    wire N__23729;
    wire N__23728;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23712;
    wire N__23703;
    wire N__23702;
    wire N__23701;
    wire N__23698;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23677;
    wire N__23674;
    wire N__23673;
    wire N__23670;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23643;
    wire N__23642;
    wire N__23641;
    wire N__23638;
    wire N__23637;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23619;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23591;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23571;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23505;
    wire N__23504;
    wire N__23501;
    wire N__23496;
    wire N__23491;
    wire N__23484;
    wire N__23481;
    wire N__23478;
    wire N__23477;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23449;
    wire N__23448;
    wire N__23445;
    wire N__23442;
    wire N__23437;
    wire N__23434;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23413;
    wire N__23412;
    wire N__23409;
    wire N__23402;
    wire N__23399;
    wire N__23394;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23366;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23349;
    wire N__23346;
    wire N__23345;
    wire N__23344;
    wire N__23343;
    wire N__23340;
    wire N__23339;
    wire N__23338;
    wire N__23335;
    wire N__23334;
    wire N__23333;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23325;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23314;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23272;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23207;
    wire N__23204;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23181;
    wire N__23176;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23139;
    wire N__23138;
    wire N__23133;
    wire N__23130;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23118;
    wire N__23115;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23085;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22956;
    wire N__22949;
    wire N__22946;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22931;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22890;
    wire N__22887;
    wire N__22882;
    wire N__22875;
    wire N__22872;
    wire N__22871;
    wire N__22870;
    wire N__22867;
    wire N__22864;
    wire N__22863;
    wire N__22862;
    wire N__22861;
    wire N__22860;
    wire N__22859;
    wire N__22858;
    wire N__22855;
    wire N__22850;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22800;
    wire N__22799;
    wire N__22798;
    wire N__22795;
    wire N__22794;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22786;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22775;
    wire N__22774;
    wire N__22773;
    wire N__22772;
    wire N__22771;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22741;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22676;
    wire N__22673;
    wire N__22666;
    wire N__22663;
    wire N__22660;
    wire N__22653;
    wire N__22650;
    wire N__22645;
    wire N__22640;
    wire N__22637;
    wire N__22632;
    wire N__22627;
    wire N__22622;
    wire N__22619;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22607;
    wire N__22606;
    wire N__22605;
    wire N__22602;
    wire N__22597;
    wire N__22594;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22571;
    wire N__22570;
    wire N__22569;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22561;
    wire N__22560;
    wire N__22559;
    wire N__22558;
    wire N__22555;
    wire N__22554;
    wire N__22553;
    wire N__22552;
    wire N__22549;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22479;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22459;
    wire N__22454;
    wire N__22451;
    wire N__22446;
    wire N__22443;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22422;
    wire N__22419;
    wire N__22418;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22377;
    wire N__22374;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22356;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22334;
    wire N__22331;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22282;
    wire N__22281;
    wire N__22278;
    wire N__22275;
    wire N__22272;
    wire N__22271;
    wire N__22268;
    wire N__22267;
    wire N__22266;
    wire N__22265;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22246;
    wire N__22243;
    wire N__22242;
    wire N__22241;
    wire N__22238;
    wire N__22237;
    wire N__22232;
    wire N__22229;
    wire N__22228;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22185;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22134;
    wire N__22133;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22111;
    wire N__22108;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22090;
    wire N__22087;
    wire N__22082;
    wire N__22079;
    wire N__22072;
    wire N__22069;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22024;
    wire N__22023;
    wire N__22022;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22008;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__22000;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21972;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21955;
    wire N__21954;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21936;
    wire N__21933;
    wire N__21932;
    wire N__21931;
    wire N__21928;
    wire N__21927;
    wire N__21924;
    wire N__21919;
    wire N__21916;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21860;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21839;
    wire N__21838;
    wire N__21835;
    wire N__21830;
    wire N__21825;
    wire N__21820;
    wire N__21815;
    wire N__21812;
    wire N__21807;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21728;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21711;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21679;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21654;
    wire N__21651;
    wire N__21650;
    wire N__21649;
    wire N__21648;
    wire N__21643;
    wire N__21640;
    wire N__21639;
    wire N__21636;
    wire N__21635;
    wire N__21634;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21618;
    wire N__21613;
    wire N__21606;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21591;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21578;
    wire N__21577;
    wire N__21576;
    wire N__21573;
    wire N__21572;
    wire N__21571;
    wire N__21570;
    wire N__21567;
    wire N__21566;
    wire N__21565;
    wire N__21564;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21550;
    wire N__21549;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21538;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21477;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21434;
    wire N__21429;
    wire N__21428;
    wire N__21427;
    wire N__21424;
    wire N__21419;
    wire N__21414;
    wire N__21405;
    wire N__21402;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21352;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21338;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21318;
    wire N__21317;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21297;
    wire N__21296;
    wire N__21293;
    wire N__21292;
    wire N__21291;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21275;
    wire N__21272;
    wire N__21271;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21260;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21214;
    wire N__21213;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21186;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21029;
    wire N__21024;
    wire N__21023;
    wire N__21022;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21010;
    wire N__21007;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20993;
    wire N__20992;
    wire N__20991;
    wire N__20990;
    wire N__20989;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20936;
    wire N__20935;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20924;
    wire N__20921;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20904;
    wire N__20895;
    wire N__20894;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20886;
    wire N__20885;
    wire N__20882;
    wire N__20881;
    wire N__20878;
    wire N__20875;
    wire N__20866;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20842;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20802;
    wire N__20801;
    wire N__20800;
    wire N__20799;
    wire N__20796;
    wire N__20791;
    wire N__20782;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20621;
    wire N__20620;
    wire N__20613;
    wire N__20610;
    wire N__20609;
    wire N__20608;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20580;
    wire N__20579;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20556;
    wire N__20553;
    wire N__20552;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20523;
    wire N__20520;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20496;
    wire N__20493;
    wire N__20492;
    wire N__20489;
    wire N__20488;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20463;
    wire N__20460;
    wire N__20459;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20441;
    wire N__20436;
    wire N__20435;
    wire N__20434;
    wire N__20433;
    wire N__20430;
    wire N__20429;
    wire N__20426;
    wire N__20421;
    wire N__20420;
    wire N__20417;
    wire N__20416;
    wire N__20415;
    wire N__20414;
    wire N__20411;
    wire N__20410;
    wire N__20409;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20358;
    wire N__20355;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20343;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20335;
    wire N__20334;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20320;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20147;
    wire N__20146;
    wire N__20141;
    wire N__20138;
    wire N__20133;
    wire N__20132;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20115;
    wire N__20114;
    wire N__20111;
    wire N__20110;
    wire N__20109;
    wire N__20108;
    wire N__20105;
    wire N__20104;
    wire N__20103;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20092;
    wire N__20091;
    wire N__20090;
    wire N__20087;
    wire N__20082;
    wire N__20079;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20036;
    wire N__20031;
    wire N__20028;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20004;
    wire N__20001;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19976;
    wire N__19975;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19948;
    wire N__19945;
    wire N__19944;
    wire N__19939;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19884;
    wire N__19879;
    wire N__19872;
    wire N__19871;
    wire N__19866;
    wire N__19863;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19691;
    wire N__19690;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19678;
    wire N__19675;
    wire N__19668;
    wire N__19667;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19652;
    wire N__19651;
    wire N__19648;
    wire N__19647;
    wire N__19644;
    wire N__19643;
    wire N__19642;
    wire N__19641;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19585;
    wire N__19576;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19545;
    wire N__19544;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19527;
    wire N__19526;
    wire N__19523;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19437;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19413;
    wire N__19410;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19396;
    wire N__19395;
    wire N__19390;
    wire N__19385;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19361;
    wire N__19360;
    wire N__19357;
    wire N__19352;
    wire N__19347;
    wire N__19344;
    wire N__19343;
    wire N__19340;
    wire N__19339;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19326;
    wire N__19317;
    wire N__19314;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19302;
    wire N__19299;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19289;
    wire N__19288;
    wire N__19285;
    wire N__19284;
    wire N__19283;
    wire N__19278;
    wire N__19273;
    wire N__19270;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19253;
    wire N__19252;
    wire N__19251;
    wire N__19250;
    wire N__19249;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19220;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19190;
    wire N__19189;
    wire N__19186;
    wire N__19181;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19151;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19134;
    wire N__19133;
    wire N__19132;
    wire N__19131;
    wire N__19124;
    wire N__19123;
    wire N__19120;
    wire N__19119;
    wire N__19116;
    wire N__19115;
    wire N__19114;
    wire N__19113;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19102;
    wire N__19099;
    wire N__19090;
    wire N__19083;
    wire N__19080;
    wire N__19075;
    wire N__19072;
    wire N__19065;
    wire N__19064;
    wire N__19063;
    wire N__19062;
    wire N__19061;
    wire N__19060;
    wire N__19059;
    wire N__19058;
    wire N__19057;
    wire N__19056;
    wire N__19055;
    wire N__19054;
    wire N__19053;
    wire N__19048;
    wire N__19039;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19025;
    wire N__19020;
    wire N__19013;
    wire N__19010;
    wire N__19009;
    wire N__19008;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__19000;
    wire N__18999;
    wire N__18998;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18980;
    wire N__18975;
    wire N__18974;
    wire N__18969;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18948;
    wire N__18945;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18920;
    wire N__18919;
    wire N__18914;
    wire N__18911;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18884;
    wire N__18883;
    wire N__18880;
    wire N__18875;
    wire N__18872;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18862;
    wire N__18859;
    wire N__18858;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18840;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18832;
    wire N__18831;
    wire N__18824;
    wire N__18821;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18794;
    wire N__18789;
    wire N__18786;
    wire N__18785;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18777;
    wire N__18774;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18760;
    wire N__18759;
    wire N__18756;
    wire N__18751;
    wire N__18748;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18732;
    wire N__18731;
    wire N__18730;
    wire N__18729;
    wire N__18726;
    wire N__18719;
    wire N__18716;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18702;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18611;
    wire N__18610;
    wire N__18609;
    wire N__18606;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18588;
    wire N__18587;
    wire N__18586;
    wire N__18585;
    wire N__18580;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18569;
    wire N__18568;
    wire N__18567;
    wire N__18566;
    wire N__18565;
    wire N__18564;
    wire N__18561;
    wire N__18560;
    wire N__18559;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18539;
    wire N__18534;
    wire N__18525;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18484;
    wire N__18483;
    wire N__18478;
    wire N__18477;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18450;
    wire N__18449;
    wire N__18446;
    wire N__18445;
    wire N__18442;
    wire N__18439;
    wire N__18436;
    wire N__18429;
    wire N__18428;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18411;
    wire N__18408;
    wire N__18407;
    wire N__18404;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18387;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18366;
    wire N__18365;
    wire N__18364;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18346;
    wire N__18339;
    wire N__18338;
    wire N__18335;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18318;
    wire N__18315;
    wire N__18312;
    wire N__18309;
    wire N__18306;
    wire N__18305;
    wire N__18304;
    wire N__18303;
    wire N__18302;
    wire N__18299;
    wire N__18294;
    wire N__18289;
    wire N__18282;
    wire N__18281;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18261;
    wire N__18260;
    wire N__18257;
    wire N__18256;
    wire N__18255;
    wire N__18252;
    wire N__18251;
    wire N__18250;
    wire N__18249;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18241;
    wire N__18240;
    wire N__18239;
    wire N__18238;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18209;
    wire N__18206;
    wire N__18201;
    wire N__18196;
    wire N__18193;
    wire N__18188;
    wire N__18185;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18161;
    wire N__18156;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18137;
    wire N__18134;
    wire N__18133;
    wire N__18130;
    wire N__18125;
    wire N__18120;
    wire N__18117;
    wire N__18116;
    wire N__18115;
    wire N__18112;
    wire N__18107;
    wire N__18102;
    wire N__18099;
    wire N__18098;
    wire N__18097;
    wire N__18094;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18080;
    wire N__18075;
    wire N__18072;
    wire N__18071;
    wire N__18070;
    wire N__18067;
    wire N__18062;
    wire N__18057;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18020;
    wire N__18019;
    wire N__18016;
    wire N__18013;
    wire N__18012;
    wire N__18011;
    wire N__18010;
    wire N__18007;
    wire N__18006;
    wire N__18001;
    wire N__17998;
    wire N__17997;
    wire N__17996;
    wire N__17993;
    wire N__17992;
    wire N__17991;
    wire N__17990;
    wire N__17989;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17968;
    wire N__17965;
    wire N__17964;
    wire N__17963;
    wire N__17960;
    wire N__17959;
    wire N__17958;
    wire N__17957;
    wire N__17956;
    wire N__17953;
    wire N__17952;
    wire N__17949;
    wire N__17948;
    wire N__17947;
    wire N__17944;
    wire N__17943;
    wire N__17942;
    wire N__17935;
    wire N__17934;
    wire N__17927;
    wire N__17924;
    wire N__17923;
    wire N__17922;
    wire N__17919;
    wire N__17916;
    wire N__17913;
    wire N__17910;
    wire N__17907;
    wire N__17906;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17898;
    wire N__17897;
    wire N__17896;
    wire N__17895;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17884;
    wire N__17881;
    wire N__17878;
    wire N__17875;
    wire N__17872;
    wire N__17869;
    wire N__17866;
    wire N__17865;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17853;
    wire N__17850;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17838;
    wire N__17833;
    wire N__17830;
    wire N__17827;
    wire N__17824;
    wire N__17821;
    wire N__17818;
    wire N__17817;
    wire N__17814;
    wire N__17811;
    wire N__17810;
    wire N__17807;
    wire N__17806;
    wire N__17805;
    wire N__17804;
    wire N__17803;
    wire N__17800;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17782;
    wire N__17775;
    wire N__17772;
    wire N__17769;
    wire N__17768;
    wire N__17767;
    wire N__17766;
    wire N__17765;
    wire N__17756;
    wire N__17753;
    wire N__17752;
    wire N__17749;
    wire N__17740;
    wire N__17739;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17715;
    wire N__17714;
    wire N__17713;
    wire N__17710;
    wire N__17709;
    wire N__17706;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17692;
    wire N__17689;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17605;
    wire N__17604;
    wire N__17603;
    wire N__17602;
    wire N__17595;
    wire N__17592;
    wire N__17581;
    wire N__17578;
    wire N__17571;
    wire N__17566;
    wire N__17559;
    wire N__17558;
    wire N__17555;
    wire N__17554;
    wire N__17551;
    wire N__17550;
    wire N__17547;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17515;
    wire N__17502;
    wire N__17499;
    wire N__17496;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17457;
    wire N__17454;
    wire N__17453;
    wire N__17450;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17411;
    wire N__17408;
    wire N__17407;
    wire N__17406;
    wire N__17405;
    wire N__17402;
    wire N__17401;
    wire N__17400;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17392;
    wire N__17391;
    wire N__17388;
    wire N__17385;
    wire N__17384;
    wire N__17381;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17349;
    wire N__17348;
    wire N__17347;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17335;
    wire N__17332;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17304;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17277;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17245;
    wire N__17242;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17203;
    wire N__17200;
    wire N__17193;
    wire N__17190;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17178;
    wire N__17177;
    wire N__17176;
    wire N__17173;
    wire N__17172;
    wire N__17171;
    wire N__17170;
    wire N__17169;
    wire N__17168;
    wire N__17167;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17136;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17122;
    wire N__17121;
    wire N__17120;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17100;
    wire N__17095;
    wire N__17092;
    wire N__17087;
    wire N__17084;
    wire N__17073;
    wire N__17072;
    wire N__17069;
    wire N__17068;
    wire N__17067;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17057;
    wire N__17052;
    wire N__17051;
    wire N__17050;
    wire N__17049;
    wire N__17048;
    wire N__17047;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17031;
    wire N__17028;
    wire N__17025;
    wire N__17022;
    wire N__17021;
    wire N__17020;
    wire N__17019;
    wire N__17018;
    wire N__17017;
    wire N__17016;
    wire N__17011;
    wire N__17004;
    wire N__16999;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16983;
    wire N__16968;
    wire N__16965;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16946;
    wire N__16945;
    wire N__16942;
    wire N__16937;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16923;
    wire N__16920;
    wire N__16919;
    wire N__16918;
    wire N__16915;
    wire N__16910;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16898;
    wire N__16895;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16883;
    wire N__16878;
    wire N__16875;
    wire N__16872;
    wire N__16869;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16859;
    wire N__16858;
    wire N__16855;
    wire N__16850;
    wire N__16845;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16830;
    wire N__16827;
    wire N__16824;
    wire N__16821;
    wire N__16820;
    wire N__16819;
    wire N__16816;
    wire N__16811;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16797;
    wire N__16794;
    wire N__16791;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16778;
    wire N__16777;
    wire N__16776;
    wire N__16775;
    wire N__16772;
    wire N__16771;
    wire N__16768;
    wire N__16767;
    wire N__16766;
    wire N__16765;
    wire N__16764;
    wire N__16761;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16753;
    wire N__16744;
    wire N__16743;
    wire N__16742;
    wire N__16737;
    wire N__16736;
    wire N__16731;
    wire N__16728;
    wire N__16725;
    wire N__16722;
    wire N__16719;
    wire N__16716;
    wire N__16713;
    wire N__16712;
    wire N__16711;
    wire N__16708;
    wire N__16707;
    wire N__16704;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16692;
    wire N__16691;
    wire N__16690;
    wire N__16687;
    wire N__16686;
    wire N__16685;
    wire N__16682;
    wire N__16677;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16659;
    wire N__16656;
    wire N__16653;
    wire N__16648;
    wire N__16645;
    wire N__16640;
    wire N__16635;
    wire N__16630;
    wire N__16611;
    wire N__16610;
    wire N__16609;
    wire N__16608;
    wire N__16603;
    wire N__16602;
    wire N__16601;
    wire N__16600;
    wire N__16599;
    wire N__16598;
    wire N__16597;
    wire N__16596;
    wire N__16593;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16583;
    wire N__16578;
    wire N__16571;
    wire N__16568;
    wire N__16565;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16550;
    wire N__16549;
    wire N__16548;
    wire N__16535;
    wire N__16534;
    wire N__16531;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16506;
    wire N__16503;
    wire N__16502;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16490;
    wire N__16489;
    wire N__16488;
    wire N__16485;
    wire N__16484;
    wire N__16483;
    wire N__16482;
    wire N__16481;
    wire N__16480;
    wire N__16479;
    wire N__16478;
    wire N__16477;
    wire N__16476;
    wire N__16475;
    wire N__16474;
    wire N__16473;
    wire N__16470;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16459;
    wire N__16458;
    wire N__16457;
    wire N__16456;
    wire N__16455;
    wire N__16452;
    wire N__16451;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16437;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16427;
    wire N__16426;
    wire N__16425;
    wire N__16424;
    wire N__16415;
    wire N__16412;
    wire N__16405;
    wire N__16400;
    wire N__16395;
    wire N__16394;
    wire N__16389;
    wire N__16386;
    wire N__16385;
    wire N__16382;
    wire N__16377;
    wire N__16370;
    wire N__16367;
    wire N__16366;
    wire N__16357;
    wire N__16354;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16333;
    wire N__16324;
    wire N__16321;
    wire N__16312;
    wire N__16307;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16280;
    wire N__16279;
    wire N__16276;
    wire N__16271;
    wire N__16266;
    wire N__16265;
    wire N__16264;
    wire N__16263;
    wire N__16260;
    wire N__16259;
    wire N__16256;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16240;
    wire N__16233;
    wire N__16230;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16220;
    wire N__16217;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16137;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16098;
    wire N__16097;
    wire N__16096;
    wire N__16095;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16084;
    wire N__16083;
    wire N__16080;
    wire N__16077;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16062;
    wire N__16061;
    wire N__16058;
    wire N__16057;
    wire N__16056;
    wire N__16053;
    wire N__16050;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16027;
    wire N__16026;
    wire N__16023;
    wire N__16022;
    wire N__16019;
    wire N__16012;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__16000;
    wire N__15999;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15989;
    wire N__15984;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15949;
    wire N__15946;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15905;
    wire N__15902;
    wire N__15897;
    wire N__15896;
    wire N__15895;
    wire N__15892;
    wire N__15887;
    wire N__15882;
    wire N__15879;
    wire N__15876;
    wire N__15875;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15860;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15845;
    wire N__15840;
    wire N__15837;
    wire N__15834;
    wire N__15833;
    wire N__15832;
    wire N__15831;
    wire N__15822;
    wire N__15819;
    wire N__15818;
    wire N__15817;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15805;
    wire N__15804;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15791;
    wire N__15790;
    wire N__15787;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15765;
    wire N__15762;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15750;
    wire N__15747;
    wire N__15744;
    wire N__15741;
    wire N__15738;
    wire N__15735;
    wire N__15732;
    wire N__15729;
    wire N__15728;
    wire N__15727;
    wire N__15724;
    wire N__15719;
    wire N__15714;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15702;
    wire N__15701;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15657;
    wire N__15654;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15614;
    wire N__15611;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15597;
    wire N__15594;
    wire N__15591;
    wire N__15590;
    wire N__15589;
    wire N__15588;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15573;
    wire N__15570;
    wire N__15567;
    wire N__15562;
    wire N__15561;
    wire N__15560;
    wire N__15559;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15541;
    wire N__15538;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15489;
    wire N__15486;
    wire N__15485;
    wire N__15482;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15464;
    wire N__15463;
    wire N__15458;
    wire N__15457;
    wire N__15456;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15429;
    wire N__15426;
    wire N__15425;
    wire N__15422;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15405;
    wire N__15404;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15396;
    wire N__15395;
    wire N__15394;
    wire N__15393;
    wire N__15392;
    wire N__15391;
    wire N__15388;
    wire N__15387;
    wire N__15382;
    wire N__15379;
    wire N__15374;
    wire N__15371;
    wire N__15366;
    wire N__15365;
    wire N__15362;
    wire N__15361;
    wire N__15360;
    wire N__15357;
    wire N__15352;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15306;
    wire N__15303;
    wire N__15302;
    wire N__15299;
    wire N__15298;
    wire N__15297;
    wire N__15296;
    wire N__15295;
    wire N__15292;
    wire N__15291;
    wire N__15288;
    wire N__15283;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15275;
    wire N__15274;
    wire N__15273;
    wire N__15272;
    wire N__15271;
    wire N__15268;
    wire N__15267;
    wire N__15264;
    wire N__15263;
    wire N__15258;
    wire N__15255;
    wire N__15250;
    wire N__15247;
    wire N__15242;
    wire N__15241;
    wire N__15240;
    wire N__15237;
    wire N__15236;
    wire N__15235;
    wire N__15234;
    wire N__15231;
    wire N__15230;
    wire N__15227;
    wire N__15226;
    wire N__15225;
    wire N__15222;
    wire N__15217;
    wire N__15214;
    wire N__15205;
    wire N__15198;
    wire N__15197;
    wire N__15194;
    wire N__15185;
    wire N__15182;
    wire N__15177;
    wire N__15166;
    wire N__15163;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15128;
    wire N__15127;
    wire N__15126;
    wire N__15125;
    wire N__15122;
    wire N__15119;
    wire N__15118;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15108;
    wire N__15107;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15093;
    wire N__15092;
    wire N__15089;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15075;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15057;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15045;
    wire N__15042;
    wire N__15039;
    wire N__15038;
    wire N__15035;
    wire N__15030;
    wire N__15027;
    wire N__15024;
    wire N__15021;
    wire N__15018;
    wire N__15015;
    wire N__15012;
    wire N__15009;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14988;
    wire N__14985;
    wire N__14982;
    wire N__14979;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14943;
    wire N__14940;
    wire N__14937;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14913;
    wire N__14904;
    wire N__14901;
    wire N__14898;
    wire N__14895;
    wire N__14892;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14867;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14838;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14826;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14814;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14799;
    wire N__14796;
    wire N__14795;
    wire N__14792;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14774;
    wire N__14769;
    wire N__14768;
    wire N__14767;
    wire N__14766;
    wire N__14765;
    wire N__14764;
    wire N__14763;
    wire N__14762;
    wire N__14761;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14733;
    wire N__14732;
    wire N__14731;
    wire N__14730;
    wire N__14729;
    wire N__14728;
    wire N__14727;
    wire N__14726;
    wire N__14725;
    wire N__14724;
    wire N__14723;
    wire N__14720;
    wire N__14697;
    wire N__14694;
    wire N__14691;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14680;
    wire N__14679;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14671;
    wire N__14666;
    wire N__14665;
    wire N__14664;
    wire N__14663;
    wire N__14660;
    wire N__14655;
    wire N__14652;
    wire N__14649;
    wire N__14642;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14619;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14607;
    wire N__14606;
    wire N__14603;
    wire N__14602;
    wire N__14601;
    wire N__14598;
    wire N__14597;
    wire N__14596;
    wire N__14593;
    wire N__14592;
    wire N__14591;
    wire N__14588;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14559;
    wire N__14552;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14523;
    wire N__14520;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14508;
    wire N__14505;
    wire N__14502;
    wire N__14501;
    wire N__14500;
    wire N__14497;
    wire N__14496;
    wire N__14495;
    wire N__14494;
    wire N__14491;
    wire N__14490;
    wire N__14489;
    wire N__14488;
    wire N__14487;
    wire N__14484;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14470;
    wire N__14469;
    wire N__14466;
    wire N__14465;
    wire N__14464;
    wire N__14461;
    wire N__14460;
    wire N__14457;
    wire N__14454;
    wire N__14451;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14439;
    wire N__14436;
    wire N__14433;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14421;
    wire N__14418;
    wire N__14415;
    wire N__14412;
    wire N__14409;
    wire N__14406;
    wire N__14403;
    wire N__14400;
    wire N__14397;
    wire N__14394;
    wire N__14391;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14356;
    wire N__14351;
    wire N__14348;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14328;
    wire N__14325;
    wire N__14322;
    wire N__14319;
    wire N__14314;
    wire N__14309;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14291;
    wire N__14286;
    wire N__14277;
    wire N__14274;
    wire N__14271;
    wire N__14268;
    wire N__14265;
    wire N__14264;
    wire N__14259;
    wire N__14258;
    wire N__14255;
    wire N__14252;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14208;
    wire N__14205;
    wire N__14202;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14175;
    wire N__14174;
    wire N__14173;
    wire N__14172;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14164;
    wire N__14161;
    wire N__14160;
    wire N__14159;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14139;
    wire N__14134;
    wire N__14121;
    wire N__14120;
    wire N__14115;
    wire N__14112;
    wire N__14109;
    wire N__14106;
    wire N__14103;
    wire N__14102;
    wire N__14101;
    wire N__14100;
    wire N__14097;
    wire N__14094;
    wire N__14093;
    wire N__14090;
    wire N__14089;
    wire N__14088;
    wire N__14087;
    wire N__14084;
    wire N__14079;
    wire N__14074;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14064;
    wire N__14057;
    wire N__14054;
    wire N__14043;
    wire N__14042;
    wire N__14041;
    wire N__14040;
    wire N__14039;
    wire N__14038;
    wire N__14033;
    wire N__14028;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14001;
    wire N__14000;
    wire N__13999;
    wire N__13998;
    wire N__13995;
    wire N__13994;
    wire N__13991;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13971;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13949;
    wire N__13938;
    wire N__13937;
    wire N__13934;
    wire N__13933;
    wire N__13932;
    wire N__13931;
    wire N__13930;
    wire N__13929;
    wire N__13928;
    wire N__13927;
    wire N__13926;
    wire N__13925;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13913;
    wire N__13908;
    wire N__13895;
    wire N__13884;
    wire N__13883;
    wire N__13882;
    wire N__13881;
    wire N__13880;
    wire N__13879;
    wire N__13878;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13870;
    wire N__13869;
    wire N__13866;
    wire N__13861;
    wire N__13858;
    wire N__13849;
    wire N__13844;
    wire N__13833;
    wire N__13830;
    wire N__13829;
    wire N__13828;
    wire N__13827;
    wire N__13826;
    wire N__13825;
    wire N__13824;
    wire N__13821;
    wire N__13816;
    wire N__13811;
    wire N__13810;
    wire N__13809;
    wire N__13808;
    wire N__13807;
    wire N__13806;
    wire N__13805;
    wire N__13802;
    wire N__13799;
    wire N__13796;
    wire N__13793;
    wire N__13790;
    wire N__13783;
    wire N__13776;
    wire N__13761;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13746;
    wire N__13743;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13724;
    wire N__13721;
    wire N__13718;
    wire N__13717;
    wire N__13716;
    wire N__13715;
    wire N__13712;
    wire N__13711;
    wire N__13708;
    wire N__13705;
    wire N__13704;
    wire N__13701;
    wire N__13700;
    wire N__13697;
    wire N__13696;
    wire N__13695;
    wire N__13692;
    wire N__13689;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13671;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13647;
    wire N__13644;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13605;
    wire N__13602;
    wire N__13601;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13571;
    wire N__13566;
    wire N__13563;
    wire N__13558;
    wire N__13555;
    wire N__13552;
    wire N__13547;
    wire N__13544;
    wire N__13539;
    wire N__13536;
    wire N__13531;
    wire N__13526;
    wire N__13521;
    wire N__13518;
    wire N__13515;
    wire N__13508;
    wire N__13505;
    wire N__13500;
    wire N__13497;
    wire N__13494;
    wire N__13493;
    wire N__13492;
    wire N__13485;
    wire N__13482;
    wire N__13479;
    wire N__13476;
    wire N__13473;
    wire N__13470;
    wire N__13467;
    wire N__13466;
    wire N__13465;
    wire N__13464;
    wire N__13463;
    wire N__13460;
    wire N__13455;
    wire N__13450;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13434;
    wire N__13431;
    wire N__13428;
    wire N__13425;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13412;
    wire N__13407;
    wire N__13404;
    wire N__13401;
    wire N__13398;
    wire N__13395;
    wire N__13392;
    wire N__13389;
    wire N__13388;
    wire N__13387;
    wire N__13386;
    wire N__13385;
    wire N__13384;
    wire N__13383;
    wire N__13378;
    wire N__13377;
    wire N__13370;
    wire N__13369;
    wire N__13368;
    wire N__13367;
    wire N__13366;
    wire N__13365;
    wire N__13364;
    wire N__13363;
    wire N__13362;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13339;
    wire N__13332;
    wire N__13325;
    wire N__13308;
    wire N__13307;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13299;
    wire N__13298;
    wire N__13297;
    wire N__13296;
    wire N__13295;
    wire N__13294;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13277;
    wire N__13276;
    wire N__13275;
    wire N__13274;
    wire N__13271;
    wire N__13270;
    wire N__13269;
    wire N__13268;
    wire N__13265;
    wire N__13264;
    wire N__13261;
    wire N__13258;
    wire N__13251;
    wire N__13248;
    wire N__13245;
    wire N__13236;
    wire N__13227;
    wire N__13212;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13172;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13158;
    wire N__13155;
    wire N__13152;
    wire N__13149;
    wire N__13148;
    wire N__13147;
    wire N__13144;
    wire N__13139;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13121;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13088;
    wire N__13087;
    wire N__13082;
    wire N__13079;
    wire N__13076;
    wire N__13071;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13043;
    wire N__13040;
    wire N__13037;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13025;
    wire N__13022;
    wire N__13019;
    wire N__13014;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12993;
    wire N__12990;
    wire N__12987;
    wire N__12984;
    wire N__12981;
    wire N__12978;
    wire N__12975;
    wire N__12972;
    wire N__12969;
    wire N__12968;
    wire N__12967;
    wire N__12966;
    wire N__12965;
    wire N__12964;
    wire N__12963;
    wire N__12958;
    wire N__12955;
    wire N__12950;
    wire N__12949;
    wire N__12946;
    wire N__12945;
    wire N__12944;
    wire N__12943;
    wire N__12940;
    wire N__12939;
    wire N__12938;
    wire N__12937;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12921;
    wire N__12918;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12891;
    wire N__12882;
    wire N__12881;
    wire N__12880;
    wire N__12879;
    wire N__12876;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12862;
    wire N__12859;
    wire N__12856;
    wire N__12855;
    wire N__12854;
    wire N__12853;
    wire N__12852;
    wire N__12851;
    wire N__12850;
    wire N__12849;
    wire N__12846;
    wire N__12841;
    wire N__12838;
    wire N__12833;
    wire N__12826;
    wire N__12823;
    wire N__12816;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12782;
    wire N__12777;
    wire N__12776;
    wire N__12773;
    wire N__12772;
    wire N__12769;
    wire N__12768;
    wire N__12767;
    wire N__12764;
    wire N__12759;
    wire N__12754;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12725;
    wire N__12724;
    wire N__12721;
    wire N__12718;
    wire N__12717;
    wire N__12714;
    wire N__12713;
    wire N__12712;
    wire N__12711;
    wire N__12708;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12678;
    wire N__12675;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12653;
    wire N__12652;
    wire N__12651;
    wire N__12648;
    wire N__12647;
    wire N__12646;
    wire N__12645;
    wire N__12642;
    wire N__12637;
    wire N__12634;
    wire N__12631;
    wire N__12626;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12605;
    wire N__12604;
    wire N__12603;
    wire N__12598;
    wire N__12597;
    wire N__12594;
    wire N__12593;
    wire N__12590;
    wire N__12589;
    wire N__12586;
    wire N__12583;
    wire N__12582;
    wire N__12581;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12546;
    wire N__12543;
    wire N__12542;
    wire N__12541;
    wire N__12540;
    wire N__12539;
    wire N__12538;
    wire N__12537;
    wire N__12534;
    wire N__12529;
    wire N__12524;
    wire N__12519;
    wire N__12510;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12486;
    wire N__12483;
    wire N__12480;
    wire N__12477;
    wire N__12474;
    wire N__12471;
    wire N__12468;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12450;
    wire N__12447;
    wire N__12444;
    wire N__12441;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12414;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12374;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12363;
    wire N__12358;
    wire N__12355;
    wire N__12352;
    wire N__12349;
    wire N__12344;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12287;
    wire N__12284;
    wire N__12283;
    wire N__12282;
    wire N__12281;
    wire N__12280;
    wire N__12277;
    wire N__12272;
    wire N__12269;
    wire N__12264;
    wire N__12255;
    wire N__12252;
    wire N__12249;
    wire N__12246;
    wire N__12243;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12219;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12206;
    wire N__12205;
    wire N__12204;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12192;
    wire N__12189;
    wire N__12180;
    wire N__12179;
    wire N__12178;
    wire N__12177;
    wire N__12176;
    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12166;
    wire N__12165;
    wire N__12160;
    wire N__12157;
    wire N__12156;
    wire N__12147;
    wire N__12142;
    wire N__12139;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12120;
    wire N__12117;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12087;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12041;
    wire N__12040;
    wire N__12039;
    wire N__12034;
    wire N__12029;
    wire N__12024;
    wire N__12021;
    wire N__12020;
    wire N__12019;
    wire N__12016;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12004;
    wire N__11997;
    wire N__11994;
    wire N__11993;
    wire N__11992;
    wire N__11987;
    wire N__11984;
    wire N__11983;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11971;
    wire N__11964;
    wire N__11961;
    wire N__11958;
    wire N__11957;
    wire N__11956;
    wire N__11955;
    wire N__11954;
    wire N__11953;
    wire N__11952;
    wire N__11947;
    wire N__11944;
    wire N__11939;
    wire N__11934;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11918;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11873;
    wire N__11872;
    wire N__11871;
    wire N__11870;
    wire N__11867;
    wire N__11866;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11841;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11801;
    wire N__11800;
    wire N__11797;
    wire N__11792;
    wire N__11787;
    wire N__11786;
    wire N__11785;
    wire N__11782;
    wire N__11777;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11711;
    wire N__11708;
    wire N__11705;
    wire N__11702;
    wire N__11697;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11664;
    wire N__11661;
    wire N__11658;
    wire N__11655;
    wire N__11652;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11613;
    wire N__11610;
    wire N__11607;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11562;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11546;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11520;
    wire N__11517;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11403;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11393;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11319;
    wire N__11316;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11286;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11271;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11217;
    wire N__11214;
    wire N__11211;
    wire N__11208;
    wire N__11205;
    wire N__11202;
    wire N__11199;
    wire N__11196;
    wire N__11193;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11169;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11151;
    wire N__11148;
    wire N__11145;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11124;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire VCCG0;
    wire GNDG0;
    wire \this_vga_signals.N_692_0 ;
    wire port_clk_c;
    wire port_data_rw_0_i;
    wire port_nmib_0_i;
    wire this_vga_signals_vvisibility_i;
    wire rgb_c_0;
    wire rgb_c_1;
    wire M_this_vga_signals_address_2;
    wire M_this_vga_signals_address_6;
    wire M_this_vga_signals_address_4;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_0_cascade_ ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.g0_0_0_0_cascade_ ;
    wire \this_vga_signals.g1_1_1_cascade_ ;
    wire \this_vga_signals.g1_1_0 ;
    wire \this_vga_signals.N_4_0_0 ;
    wire \this_vga_signals.mult1_un47_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d_1 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d_1_cascade_ ;
    wire \this_vga_signals.g2_1_cascade_ ;
    wire \this_vga_signals.g2 ;
    wire \this_vga_signals.vsync_1_3_cascade_ ;
    wire this_vga_signals_vsync_1_i;
    wire \this_vga_signals.g0_2_0_cascade_ ;
    wire \this_vga_signals.N_43_1_cascade_ ;
    wire \this_vga_signals.un2_vsynclt8 ;
    wire \this_vga_signals.vsync_1_2 ;
    wire \this_vga_signals.g1_1 ;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire \this_vga_signals.g0_0_0 ;
    wire M_this_map_address_qZ0Z_0;
    wire bfn_9_23_0_;
    wire M_this_map_address_qZ0Z_1;
    wire un1_M_this_map_address_q_cry_0;
    wire M_this_map_address_qZ0Z_2;
    wire un1_M_this_map_address_q_cry_1;
    wire M_this_map_address_qZ0Z_3;
    wire un1_M_this_map_address_q_cry_2;
    wire M_this_map_address_qZ0Z_4;
    wire un1_M_this_map_address_q_cry_3;
    wire M_this_map_address_qZ0Z_5;
    wire un1_M_this_map_address_q_cry_4;
    wire M_this_map_address_qZ0Z_6;
    wire un1_M_this_map_address_q_cry_5;
    wire M_this_map_address_qZ0Z_7;
    wire un1_M_this_map_address_q_cry_6;
    wire un1_M_this_map_address_q_cry_7;
    wire M_this_map_address_qZ0Z_8;
    wire bfn_9_24_0_;
    wire un1_M_this_map_address_q_cry_8;
    wire M_this_map_address_qZ0Z_9;
    wire N_89_0;
    wire N_83_0;
    wire N_85_0;
    wire \this_vga_signals.vaddress_3_0_5_cascade_ ;
    wire \this_vga_signals.g0_6_0_0_0 ;
    wire \this_vga_signals.SUM_2_i_1_1_3_cascade_ ;
    wire \this_vga_signals.SUM_2_i_1_1_1_3 ;
    wire \this_vga_signals.N_1_3_1 ;
    wire \this_vga_signals.N_1_3_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_9 ;
    wire \this_vga_signals.vaddress_1_0_5_cascade_ ;
    wire \this_vga_signals.un6_vvisibilitylt8_cascade_ ;
    wire \this_vga_signals.vvisibility_1 ;
    wire \this_vga_signals.vaddress_0_5 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_3_cascade_ ;
    wire \this_vga_signals.g0_6_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d ;
    wire \this_vga_signals.i6_mux_0 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_ ;
    wire \this_vga_signals.g0_i_x4_0_a2_1 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_2 ;
    wire \this_vga_signals.SUM_3_1_tz ;
    wire this_vga_signals_hvisibility_i;
    wire M_stage_q_RNIC68K4_9;
    wire \this_vga_signals.vaddress_3_5 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_5_cascade_ ;
    wire \this_vga_signals.g0_6_0_0 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_0 ;
    wire \this_vga_signals.N_5_i_0_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.M_vcounter_q_8_repZ0Z1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_9_repZ0Z1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_0 ;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ;
    wire \this_vga_signals.vaddress_c2 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_cascade_ ;
    wire \this_vga_signals.g1_0_0_0 ;
    wire \this_vga_signals.vaddress_2_5 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_x0_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_5_repZ0Z1 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_1 ;
    wire \this_vga_signals.if_N_5_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z1 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_cascade_ ;
    wire \this_vga_signals.if_m8_0_a3_1_1_6 ;
    wire \this_vga_signals.N_5_i_0 ;
    wire \this_vga_signals.g1_2_1_0_0_cascade_ ;
    wire \this_vga_signals.g1_0_4_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_c3_2_0 ;
    wire \this_vga_signals.g1_0_4 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_4 ;
    wire \this_vga_signals.g1_0 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0_cascade_ ;
    wire \this_vga_signals.g0_1_0_0_0 ;
    wire \this_vga_signals.g2_1_0_1_cascade_ ;
    wire \this_vga_signals.g3_0_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_0_0 ;
    wire \this_vga_signals.M_hcounter_d7lt7_0_cascade_ ;
    wire \this_vga_signals.if_m2_0_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_c3_0_1_cascade_ ;
    wire \this_vga_signals.haddress_1_0_cascade_ ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.M_hcounter_d7lto7_1 ;
    wire \this_vga_signals.un2_hsynclto3_0 ;
    wire \this_vga_signals.un2_hsynclto3_0_cascade_ ;
    wire \this_vga_signals.un2_hsynclto6_0_cascade_ ;
    wire rgb_c_4;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire bfn_11_23_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_11_24_0_;
    wire \this_vga_signals.N_692_1 ;
    wire \this_vga_signals.M_vcounter_q_379_0 ;
    wire \this_vga_signals.g0_3_x0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_0 ;
    wire \this_vga_signals.g1_0_1_cascade_ ;
    wire \this_vga_signals.g0_i_x4_0_0 ;
    wire \this_vga_signals.g1 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d_0_1 ;
    wire \this_vga_signals.g0_1_0_0 ;
    wire \this_vga_signals.g1_2_1_cascade_ ;
    wire \this_vga_signals.g0_0_0_0_0 ;
    wire \this_vga_signals.g0_2_0_a2_1 ;
    wire \this_vga_signals.g0_2_0_a2_1_cascade_ ;
    wire \this_vga_signals.g0_3_x1 ;
    wire \this_vga_signals.g0_13_x0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb1_1 ;
    wire \this_vga_signals.mult1_un47_sum_c3_1 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d_2 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d_2_cascade_ ;
    wire \this_vga_signals.g0_13_x1 ;
    wire \this_vga_signals.mult1_un47_sum_c3 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_x0 ;
    wire \this_vga_signals.mult1_un61_sum_c3_cascade_ ;
    wire \this_vga_signals.vaddress_5 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_x1 ;
    wire \this_vga_signals.g1_2_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_d_0_0 ;
    wire \this_vga_signals.M_vcounter_q_RNITVMCUZ0Z_3_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_RNIANU4QZ0Z_3 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_2 ;
    wire \this_vga_signals.g2_0_0_cascade_ ;
    wire \this_vga_signals.g0_0_0_a3_0 ;
    wire \this_vga_signals.vaddress_c3_0 ;
    wire \this_vga_signals.SUM_2_i_1_1_3 ;
    wire \this_vga_signals.SUM_2_i_1_2_3 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i_0_cascade_ ;
    wire \this_vga_signals.g0_i_x4_0 ;
    wire \this_vga_signals.g0_i_x4_4_1_cascade_ ;
    wire \this_vga_signals.g0_i_x4_4 ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0 ;
    wire \this_vga_signals.g2_0 ;
    wire \this_vga_signals.g0_2_0_a2 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_ns ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_571 ;
    wire \this_vga_signals.mult1_un61_sum_c3 ;
    wire \this_vga_signals.N_4_0_0_1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_cascade_ ;
    wire M_this_vga_signals_address_3;
    wire \this_vga_signals.if_m2_0 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_c3_0 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3 ;
    wire M_this_vga_signals_address_1;
    wire \this_vga_signals.mult1_un75_sum_axb1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb2_1 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire M_this_vga_signals_address_5;
    wire \this_vga_signals.SUM_3 ;
    wire \this_vga_signals.SUM_3_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0 ;
    wire \this_vga_signals.N_6_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_0_0_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.un4_hsynclt4_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire N_91_0;
    wire N_93_0;
    wire M_this_map_ram_read_data_3;
    wire M_this_ppu_sprites_addr_9;
    wire M_this_map_ram_read_data_0;
    wire M_this_ppu_sprites_addr_6;
    wire bfn_13_17_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire bfn_13_18_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.N_692_0_g ;
    wire \this_vga_signals.N_988_g ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.un4_hsynclt8_0 ;
    wire \this_vga_signals.un2_hsynclt8_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire this_vga_signals_hsync_1_i;
    wire rgb_c_3;
    wire N_95_0;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire M_this_map_ram_read_data_2;
    wire M_this_ppu_sprites_addr_8;
    wire \this_vga_ramdac.N_24_mux ;
    wire \this_vga_ramdac.N_2862_reto ;
    wire this_pixel_clk_M_counter_q_i_1;
    wire rgb_c_2;
    wire \this_vga_ramdac.m6 ;
    wire \this_vga_ramdac.N_2863_reto ;
    wire \this_vga_ramdac.i2_mux_0 ;
    wire \this_vga_ramdac.m19 ;
    wire \this_vga_ramdac.N_2866_reto ;
    wire \this_vga_signals.M_this_vga_signals_pixel_clk_0_0 ;
    wire M_this_vga_ramdac_en_0;
    wire M_pcounter_q_ret_2_RNIH7PG8_cascade_;
    wire \this_vga_ramdac.i2_mux ;
    wire \this_vga_ramdac.N_2864_reto ;
    wire dma_0_i;
    wire \this_vga_signals.M_pcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_pcounter_q_3_0 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_pcounter_q_3_1 ;
    wire \this_vga_signals.N_3_0 ;
    wire \this_vga_signals.N_3_0_cascade_ ;
    wire \this_vga_signals.M_pcounter_q_i_3_1 ;
    wire \this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ;
    wire \this_vga_ramdac.N_2867_reto ;
    wire rgb_c_5;
    wire \this_vga_signals.N_2_0 ;
    wire \this_vga_signals.M_pcounter_q_i_3_0 ;
    wire bfn_14_25_0_;
    wire M_this_data_count_q_cry_0;
    wire M_this_data_count_q_cry_1;
    wire M_this_data_count_q_cry_2;
    wire M_this_data_count_q_cry_3;
    wire M_this_data_count_q_cry_4;
    wire M_this_data_count_q_cry_5;
    wire M_this_data_count_q_cry_6;
    wire M_this_data_count_q_cry_7;
    wire bfn_14_26_0_;
    wire M_this_data_count_q_cry_8;
    wire M_this_data_count_q_s_10;
    wire M_this_data_count_q_cry_9;
    wire M_this_data_count_q_cry_10;
    wire M_this_data_count_q_cry_11;
    wire M_this_data_count_q_cry_12;
    wire M_this_data_count_q_s_13;
    wire N_87_0;
    wire N_81_0;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_vcounter_d7lt8_0 ;
    wire \this_vga_signals.M_vcounter_d7lto8_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_d8_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ;
    wire this_pixel_clk_M_counter_q_0;
    wire M_pcounter_q_ret_2_RNIH7PG8;
    wire \this_vga_ramdac.N_2865_reto ;
    wire dma_ac0_5_0_cascade_;
    wire M_this_state_q_RNIOE1SZ0Z_11;
    wire un20_i_a2_x_3;
    wire M_this_state_q_RNIG01LZ0Z_12;
    wire \this_vga_signals.N_419_i_i_0Z0Z_1_cascade_ ;
    wire M_this_data_count_q_s_6;
    wire M_this_data_count_qZ0Z_6;
    wire M_this_data_count_q_cry_3_THRU_CO;
    wire M_this_data_count_qZ0Z_4;
    wire M_this_data_count_q_cry_4_THRU_CO;
    wire M_this_data_count_qZ0Z_5;
    wire M_this_data_count_q_cry_6_THRU_CO;
    wire M_this_data_count_qZ0Z_7;
    wire M_this_data_count_q_cry_2_THRU_CO;
    wire M_this_data_count_q_cry_10_THRU_CO;
    wire M_this_data_count_q_cry_11_THRU_CO;
    wire M_this_data_count_qZ0Z_12;
    wire M_this_data_count_qZ0Z_13;
    wire M_this_data_count_q_cry_7_THRU_CO;
    wire M_this_data_count_qZ0Z_8;
    wire M_this_data_count_q_cry_1_THRU_CO;
    wire M_this_data_count_q_cry_8_THRU_CO;
    wire M_this_data_count_qZ0Z_9;
    wire M_this_map_ram_read_data_1;
    wire M_this_ppu_sprites_addr_7;
    wire \this_ppu.M_count_d_0_sqmuxa_1_7_cascade_ ;
    wire \this_vga_signals.un4_lvisibility_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire bfn_16_19_0_;
    wire \this_ppu.un1_M_count_q_1_cry_0_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_1_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_2_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_3_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_4_s1 ;
    wire CONSTANT_ONE_NET;
    wire \this_ppu.un1_M_count_q_1_cry_5_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_6_s1 ;
    wire \this_ppu.M_count_q_RNO_0Z0Z_7 ;
    wire \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ;
    wire \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ;
    wire \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ;
    wire \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_5 ;
    wire \this_ppu.M_count_qZ0Z_4 ;
    wire \this_ppu.M_count_qZ0Z_6 ;
    wire \this_ppu.M_count_qZ0Z_2 ;
    wire \this_ppu.M_count_d_1_sqmuxa_1_i_a2_4 ;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire \this_vga_signals.un20_i_a2_sxZ0Z_3_cascade_ ;
    wire \this_vga_signals.N_322_cascade_ ;
    wire this_vga_signals_M_this_state_q_ns_i_o3_0_10;
    wire M_this_state_qZ0Z_10;
    wire N_212;
    wire N_160_0;
    wire M_this_state_qc_3_1;
    wire \this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_4_cascade_ ;
    wire N_465_0;
    wire N_610_0_i;
    wire M_this_data_count_q_cry_0_THRU_CO;
    wire M_this_data_count_qe_0_i;
    wire M_this_data_count_qZ0Z_3;
    wire M_this_data_count_qZ0Z_2;
    wire M_this_data_count_qZ0Z_1;
    wire M_this_data_count_qZ0Z_10;
    wire M_this_data_count_qZ0Z_11;
    wire M_this_data_count_qZ0Z_0;
    wire \this_vga_signals.M_this_state_d55Z0Z_9 ;
    wire \this_vga_signals.M_this_state_d55Z0Z_8 ;
    wire \this_vga_signals.M_this_state_d55Z0Z_7_cascade_ ;
    wire \this_vga_signals.M_this_state_d55Z0Z_6 ;
    wire M_this_vram_read_data_2;
    wire M_this_vram_read_data_1;
    wire M_this_vram_read_data_3;
    wire M_this_vram_read_data_0;
    wire \this_vga_ramdac.m16 ;
    wire \this_reset_cond.M_stage_qZ0Z_5 ;
    wire \this_reset_cond.M_stage_qZ0Z_8 ;
    wire \this_reset_cond.M_stage_qZ0Z_6 ;
    wire \this_reset_cond.M_stage_qZ0Z_7 ;
    wire \this_ppu.M_count_qZ0Z_7 ;
    wire \this_ppu.M_count_d_1_sqmuxa_1_i_a2_3 ;
    wire \this_ppu.N_132_0_cascade_ ;
    wire \this_ppu.M_count_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_d8 ;
    wire \this_vga_signals.un1_M_hcounter_d7_1_0_cascade_ ;
    wire \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_1 ;
    wire \this_vga_signals.M_hcounter_d7_0 ;
    wire \this_vga_signals.GZ0Z_330 ;
    wire \this_vga_signals.un1_M_hcounter_d7_1_0 ;
    wire \this_vga_signals.CO0_cascade_ ;
    wire \this_ppu.N_1157_0_1 ;
    wire \this_ppu.un16_0 ;
    wire \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ;
    wire \this_ppu.un16_0_cascade_ ;
    wire \this_ppu.N_1157_0 ;
    wire \this_ppu.M_count_qZ0Z_3 ;
    wire N_459_0_cascade_;
    wire N_458_0_cascade_;
    wire this_vga_signals_N_419_i_i_0_a3_1_0;
    wire N_496_0_cascade_;
    wire N_278;
    wire M_this_state_qsr_0_cascade_;
    wire N_462_0;
    wire M_this_state_qsr_2_cascade_;
    wire N_484_0;
    wire \this_vga_signals.N_159_0_cascade_ ;
    wire M_this_state_qZ0Z_9;
    wire N_168_0;
    wire N_168_0_cascade_;
    wire \this_vga_signals.M_this_external_address_d_0_sqmuxa_1Z0Z_2 ;
    wire M_this_state_qZ0Z_11;
    wire N_456_0_1;
    wire N_500;
    wire M_this_sprites_ram_write_data_0;
    wire M_this_state_d_2_sqmuxa;
    wire M_this_substate_qZ0;
    wire this_vga_signals_M_this_state_q_ns_0_a3_0_0_1;
    wire \this_sprites_ram.mem_out_bus7_0 ;
    wire \this_sprites_ram.mem_out_bus3_0 ;
    wire \this_sprites_ram.mem_out_bus6_0 ;
    wire \this_sprites_ram.mem_out_bus2_0 ;
    wire \this_sprites_ram.mem_out_bus5_0 ;
    wire \this_sprites_ram.mem_out_bus1_0 ;
    wire \this_sprites_ram.mem_out_bus4_0 ;
    wire \this_sprites_ram.mem_out_bus0_0 ;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_ ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_ ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire \this_reset_cond.M_stage_qZ0Z_3 ;
    wire \this_reset_cond.M_stage_qZ0Z_4 ;
    wire \this_sprites_ram.mem_out_bus4_2 ;
    wire \this_sprites_ram.mem_out_bus0_2 ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ;
    wire M_this_map_ram_read_data_7;
    wire \this_sprites_ram.mem_out_bus7_2 ;
    wire \this_sprites_ram.mem_out_bus3_2 ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ;
    wire \this_vga_signals.M_lcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_lcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire \this_vga_signals.line_clk_1 ;
    wire M_this_sprites_ram_write_data_3;
    wire \this_vga_signals.N_169_0 ;
    wire N_210_cascade_;
    wire \this_vga_signals.N_159_0 ;
    wire \this_vga_signals.N_167_0_cascade_ ;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_5_cascade_ ;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_6 ;
    wire M_this_state_d55;
    wire this_vga_signals_M_this_state_q_ns_i_o3_0_7_cascade_;
    wire \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3Z0Z_0 ;
    wire \this_vga_signals.N_279 ;
    wire M_this_state_qZ0Z_6;
    wire N_210;
    wire M_this_state_qZ0Z_5;
    wire \this_vga_signals.N_166 ;
    wire M_this_state_qZ0Z_3;
    wire \this_sprites_ram.mem_out_bus5_1 ;
    wire \this_sprites_ram.mem_out_bus1_1 ;
    wire M_this_map_ram_read_data_5;
    wire M_this_ppu_vram_data_3;
    wire M_this_ppu_vram_data_2;
    wire M_this_ppu_vram_data_3_cascade_;
    wire M_this_ppu_vram_data_0;
    wire \this_ppu.N_156_cascade_ ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3 ;
    wire \this_sprites_ram.mem_out_bus5_2 ;
    wire \this_sprites_ram.mem_out_bus1_2 ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ;
    wire \this_ppu.un1_M_haddress_q_3_c2_cascade_ ;
    wire \this_ppu.un1_M_haddress_q_3_c5 ;
    wire \this_sprites_ram.mem_out_bus6_3 ;
    wire \this_sprites_ram.mem_out_bus2_3 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus7_3 ;
    wire \this_sprites_ram.mem_out_bus3_3 ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire this_start_data_delay_M_last_q;
    wire port_enb_c;
    wire M_this_delay_clk_out_0;
    wire N_156_0_cascade_;
    wire N_35_0;
    wire port_rw_in;
    wire led_c_1;
    wire N_459_0;
    wire un1_M_this_state_q_12_0;
    wire bfn_19_22_0_;
    wire un1_M_this_sprites_address_q_cry_0;
    wire un1_M_this_sprites_address_q_cry_1;
    wire un1_M_this_sprites_address_q_cry_2;
    wire un1_M_this_sprites_address_q_cry_3;
    wire M_this_sprites_address_qZ0Z_5;
    wire un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0;
    wire un1_M_this_sprites_address_q_cry_4;
    wire M_this_sprites_address_qZ0Z_6;
    wire un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0;
    wire un1_M_this_sprites_address_q_cry_5;
    wire un1_M_this_sprites_address_q_cry_6;
    wire un1_M_this_sprites_address_q_cry_7;
    wire bfn_19_23_0_;
    wire un1_M_this_sprites_address_q_cry_8;
    wire un1_M_this_sprites_address_q_cry_9;
    wire un1_M_this_sprites_address_q_cry_10;
    wire un1_M_this_sprites_address_q_cry_11;
    wire un1_M_this_sprites_address_q_cry_12;
    wire M_this_state_d25;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_9_cascade_ ;
    wire un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0;
    wire M_this_sprites_address_qZ0Z_9;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_2_cascade_ ;
    wire un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0;
    wire M_this_sprites_address_qZ0Z_2;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3_cascade_ ;
    wire un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_ ;
    wire un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0;
    wire M_this_sprites_address_qZ0Z_7;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_7 ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ;
    wire M_this_ppu_vram_data_1;
    wire \this_sprites_ram.mem_WE_14 ;
    wire \this_sprites_ram.mem_out_bus7_1 ;
    wire \this_sprites_ram.mem_out_bus3_1 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus4_3 ;
    wire \this_sprites_ram.mem_out_bus0_3 ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ;
    wire this_vga_signals_vvisibility;
    wire dma_0;
    wire \this_ppu.N_150_cascade_ ;
    wire M_this_reset_cond_out_0;
    wire M_this_ppu_sprites_addr_2;
    wire M_this_ppu_vram_en_0;
    wire \this_ppu.N_156 ;
    wire \this_ppu.un2_hscroll_axb_0_cascade_ ;
    wire M_this_ppu_sprites_addr_0;
    wire \this_ppu.un1_M_haddress_q_3_c2 ;
    wire \this_ppu.M_state_q_RNIGL6V4Z0Z_0 ;
    wire \this_sprites_ram.mem_WE_8 ;
    wire \this_ppu.N_1046_0_cascade_ ;
    wire \this_ppu.M_state_qZ0Z_5 ;
    wire \this_ppu.un1_M_oam_idx_q_1_c1_cascade_ ;
    wire \this_ppu.un1_M_oam_idx_q_1_c3 ;
    wire M_this_ppu_oam_addr_2;
    wire M_this_ppu_oam_addr_0;
    wire \this_ppu.M_oam_idx_qZ0Z_4 ;
    wire \this_ppu.N_144_4_cascade_ ;
    wire \this_ppu.M_state_qZ0Z_4 ;
    wire \this_ppu.N_1046_0 ;
    wire \this_ppu.un1_M_oam_idx_q_1_c1 ;
    wire M_this_ppu_oam_addr_1;
    wire M_this_ppu_oam_addr_3;
    wire \this_ppu.N_144_4 ;
    wire \this_ppu.N_144 ;
    wire M_this_state_qZ0Z_8;
    wire M_this_state_qZ0Z_7;
    wire M_this_sprites_ram_write_data_2;
    wire \this_sprites_ram.mem_WE_6 ;
    wire un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13 ;
    wire un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12 ;
    wire un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0 ;
    wire M_this_sprites_address_q_RNIQ61C7Z0Z_0;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_0 ;
    wire M_this_sprites_address_qZ0Z_0;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_11 ;
    wire M_this_substate_q_RNOZ0Z_1;
    wire M_this_substate_q_s_1;
    wire this_vga_signals_M_this_state_d_2_sqmuxa_0;
    wire N_17_0;
    wire M_this_sprites_address_qZ0Z_3;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_3 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_12 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_13 ;
    wire M_this_state_qZ0Z_2;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_10_cascade_ ;
    wire un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0;
    wire M_this_sprites_address_qZ0Z_10;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10 ;
    wire M_this_substate_q_RNOZ0Z_3;
    wire \this_sprites_ram.mem_out_bus0_1 ;
    wire \this_sprites_ram.mem_out_bus4_1 ;
    wire \this_sprites_ram.mem_radregZ0Z_11 ;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_ ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1 ;
    wire \this_sprites_ram.mem_out_bus6_1 ;
    wire \this_sprites_ram.mem_out_bus2_1 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ;
    wire \this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ;
    wire bfn_21_16_0_;
    wire \this_ppu.un2_hscroll_cry_0 ;
    wire \this_ppu.un2_hscroll_cry_1 ;
    wire \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0 ;
    wire \this_sprites_ram.mem_WE_12 ;
    wire \this_sprites_ram.mem_out_bus6_2 ;
    wire \this_sprites_ram.mem_out_bus2_2 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ;
    wire M_this_oam_ram_read_data_i_9;
    wire \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0 ;
    wire M_this_ppu_sprites_addr_1;
    wire M_this_ppu_vram_addr_0;
    wire bfn_21_18_0_;
    wire M_this_ppu_vram_addr_1;
    wire \this_ppu.un1_M_haddress_q_2_cry_0 ;
    wire M_this_ppu_vram_addr_2;
    wire \this_ppu.un1_M_haddress_q_2_cry_1 ;
    wire M_this_oam_ram_read_data_i_11;
    wire M_this_ppu_map_addr_0;
    wire \this_ppu.un1_M_haddress_q_2_cry_2 ;
    wire \this_ppu.un1_M_haddress_q_2_4 ;
    wire M_this_ppu_map_addr_1;
    wire \this_ppu.un1_M_haddress_q_2_cry_3 ;
    wire M_this_ppu_map_addr_2;
    wire \this_ppu.un1_M_haddress_q_2_cry_4 ;
    wire M_this_ppu_map_addr_3;
    wire \this_ppu.un1_M_haddress_q_2_cry_5 ;
    wire M_this_ppu_map_addr_4;
    wire \this_ppu.un1_M_haddress_q_2_cry_6 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_7 ;
    wire bfn_21_19_0_;
    wire \this_ppu.vscroll8 ;
    wire \this_ppu.M_state_qZ0Z_2 ;
    wire N_48_0;
    wire M_this_oam_ram_write_data_28;
    wire \this_ppu.M_state_qZ0Z_3 ;
    wire \this_ppu.M_state_qZ0Z_1 ;
    wire \this_ppu.M_count_d_0_sqmuxa_1_7 ;
    wire \this_ppu.N_148 ;
    wire M_this_data_tmp_qZ0Z_20;
    wire \this_sprites_ram.mem_WE_4 ;
    wire M_this_state_d22;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11 ;
    wire port_address_in_0;
    wire \this_vga_signals.M_this_state_d21Z0Z_6 ;
    wire \this_vga_signals.M_this_state_dZ0Z24 ;
    wire \this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_8 ;
    wire un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0;
    wire M_this_sprites_address_qZ0Z_8;
    wire M_this_state_qZ0Z_1;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_1_cascade_ ;
    wire un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0;
    wire M_this_sprites_address_qZ0Z_1;
    wire \this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4 ;
    wire \this_vga_signals.un1_M_this_state_q_14_0 ;
    wire \this_vga_signals.M_this_sprites_address_q_mZ0Z_4 ;
    wire un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0;
    wire M_this_sprites_address_qZ0Z_4;
    wire \this_vga_signals.M_this_state_q_ns_8 ;
    wire \this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ;
    wire M_this_sprites_ram_write_data_1;
    wire M_this_map_ram_read_data_4;
    wire M_this_ppu_sprites_addr_10;
    wire M_this_ppu_sprites_addr_4;
    wire \this_ppu.un1_M_vaddress_q_2_c5 ;
    wire bfn_22_17_0_;
    wire \this_ppu.un1_M_vaddress_q_3_cry_0 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_1 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_2 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_3 ;
    wire M_this_ppu_map_addr_7;
    wire \this_ppu.un1_M_vaddress_q_3_cry_4 ;
    wire M_this_ppu_map_addr_8;
    wire \this_ppu.un1_M_vaddress_q_3_cry_5 ;
    wire M_this_ppu_map_addr_9;
    wire \this_ppu.un1_M_vaddress_q_3_cry_6 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_7 ;
    wire bfn_22_18_0_;
    wire \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO ;
    wire \this_ppu.un1_M_haddress_q_2_5 ;
    wire un1_M_this_oam_address_q_c3_cascade_;
    wire M_this_data_tmp_qZ0Z_7;
    wire N_65_0;
    wire \this_ppu.M_this_ppu_vram_addr_i_0 ;
    wire M_this_oam_ram_read_data_8;
    wire bfn_22_19_0_;
    wire \this_ppu.M_this_ppu_vram_addr_i_1 ;
    wire M_this_oam_ram_read_data_9;
    wire \this_ppu.un1_M_haddress_q_cry_0 ;
    wire \this_ppu.M_this_ppu_vram_addr_i_2 ;
    wire M_this_oam_ram_read_data_10;
    wire \this_ppu.un1_M_haddress_q_cry_1 ;
    wire \this_ppu.M_this_ppu_map_addr_i_0 ;
    wire \this_ppu.un1_M_haddress_q_cry_2 ;
    wire \this_ppu.M_this_ppu_map_addr_i_1 ;
    wire \this_ppu.un1_M_haddress_q_cry_3 ;
    wire \this_ppu.M_this_ppu_map_addr_i_2 ;
    wire \this_ppu.un1_M_haddress_q_cry_4 ;
    wire \this_ppu.M_this_ppu_map_addr_i_3 ;
    wire \this_ppu.un1_M_haddress_q_cry_5 ;
    wire \this_ppu.M_this_ppu_map_addr_i_4 ;
    wire \this_ppu.un1_M_haddress_q_cry_6 ;
    wire \this_ppu.un1_M_haddress_q_cry_7 ;
    wire bfn_22_20_0_;
    wire \this_ppu.vscroll8_1 ;
    wire port_address_in_5;
    wire port_address_in_6;
    wire port_address_in_7;
    wire M_this_state_qZ0Z_12;
    wire N_56_0;
    wire M_this_data_tmp_qZ0Z_13;
    wire M_this_state_d21_1;
    wire port_address_in_4;
    wire port_address_in_2;
    wire M_this_state_d21_6_x;
    wire M_this_substate_q_RNOZ0Z_2;
    wire port_address_in_3;
    wire port_address_in_1;
    wire \this_vga_signals.M_this_state_d24Z0Z_1 ;
    wire \this_sprites_ram.mem_WE_0 ;
    wire M_this_data_tmp_qZ0Z_15;
    wire M_this_oam_ram_write_data_15;
    wire \this_ppu.M_this_oam_ram_read_data_i_16 ;
    wire bfn_23_16_0_;
    wire \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0 ;
    wire \this_ppu.un2_vscroll_cry_0 ;
    wire \this_ppu.un2_vscroll_cry_1 ;
    wire M_this_map_ram_read_data_6;
    wire \this_sprites_ram.mem_radregZ0Z_12 ;
    wire \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0 ;
    wire M_this_ppu_sprites_addr_5;
    wire \this_ppu.M_vaddress_qZ0Z_1 ;
    wire \this_ppu.N_132_0 ;
    wire \this_ppu.M_state_qZ0Z_6 ;
    wire \this_ppu.un2_vscroll_axb_0_cascade_ ;
    wire \this_ppu.M_state_qZ0Z_7 ;
    wire M_this_ppu_sprites_addr_3;
    wire \this_ppu.M_vaddress_qZ0Z_2 ;
    wire \this_ppu.un1_M_vaddress_q_2_c2 ;
    wire M_this_ppu_map_addr_5;
    wire M_this_ppu_map_addr_6;
    wire \this_ppu.M_state_qZ0Z_0 ;
    wire \this_ppu.M_last_q ;
    wire M_this_vga_signals_line_clk_0;
    wire M_this_ppu_vram_addr_7;
    wire \this_ppu.M_state_q_RNI42KTAZ0Z_0 ;
    wire M_this_data_tmp_qZ0Z_4;
    wire N_71_0;
    wire \this_ppu.M_this_ppu_vram_addr_i_7 ;
    wire M_this_oam_ram_read_data_16;
    wire bfn_23_19_0_;
    wire \this_ppu.M_vaddress_q_i_1 ;
    wire \this_ppu.un1_M_vaddress_q_cry_0 ;
    wire \this_ppu.M_vaddress_q_i_2 ;
    wire M_this_oam_ram_read_data_18;
    wire \this_ppu.un1_M_vaddress_q_cry_1 ;
    wire \this_ppu.M_this_ppu_map_addr_i_5 ;
    wire \this_ppu.un1_M_vaddress_q_cry_2 ;
    wire \this_ppu.M_this_ppu_map_addr_i_6 ;
    wire \this_ppu.un1_M_vaddress_q_cry_3 ;
    wire \this_ppu.M_this_ppu_map_addr_i_7 ;
    wire \this_ppu.un1_M_vaddress_q_cry_4 ;
    wire \this_ppu.M_this_ppu_map_addr_i_8 ;
    wire \this_ppu.un1_M_vaddress_q_cry_5 ;
    wire \this_ppu.M_this_ppu_map_addr_i_9 ;
    wire \this_ppu.un1_M_vaddress_q_cry_6 ;
    wire \this_ppu.un1_M_vaddress_q_cry_7 ;
    wire bfn_23_20_0_;
    wire \this_ppu.un1_M_vaddress_q_cry_7_THRU_CO ;
    wire N_61_0;
    wire M_this_data_tmp_qZ0Z_3;
    wire N_73_0;
    wire M_this_oam_address_qZ0Z_4;
    wire M_this_oam_address_qZ0Z_5;
    wire N_1152_0;
    wire M_this_oam_address_qZ0Z_3;
    wire M_this_oam_address_qZ0Z_2;
    wire un1_M_this_oam_address_q_c2;
    wire un1_M_this_oam_address_q_c4;
    wire N_50_0;
    wire N_46_0;
    wire M_this_data_tmp_qZ0Z_21;
    wire M_this_data_tmp_qZ0Z_10;
    wire \this_sprites_ram.mem_out_bus5_3 ;
    wire \this_sprites_ram.mem_out_bus1_3 ;
    wire \this_sprites_ram.mem_radregZ0Z_13 ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ;
    wire \this_sprites_ram.mem_WE_10 ;
    wire M_this_oam_ram_read_data_17;
    wire M_this_oam_ram_read_data_i_17;
    wire M_this_oam_ram_read_data_2;
    wire M_this_oam_ram_read_data_1;
    wire M_this_oam_ram_read_data_0;
    wire M_this_oam_ram_read_data_3;
    wire \this_ppu.un9lto7Z0Z_5 ;
    wire \this_ppu.un1_M_haddress_q_2_6 ;
    wire M_this_oam_ram_read_data_4;
    wire M_this_oam_ram_read_data_6;
    wire M_this_oam_ram_read_data_7;
    wire M_this_oam_ram_read_data_5;
    wire \this_ppu.un9lto7Z0Z_4 ;
    wire \this_ppu.un1_M_vaddress_q_3_4 ;
    wire M_this_oam_ram_read_data_11;
    wire M_this_oam_ram_read_data_12;
    wire M_this_oam_ram_read_data_15;
    wire M_this_oam_ram_read_data_14;
    wire \this_ppu.un1_oam_data_1_c2_cascade_ ;
    wire M_this_oam_ram_read_data_13;
    wire \this_ppu.un1_M_haddress_q_2_7 ;
    wire M_this_data_tmp_qZ0Z_6;
    wire N_67_0;
    wire M_this_oam_ram_read_data_23;
    wire \this_ppu.un1_oam_data_c2_cascade_ ;
    wire \this_ppu.un1_M_vaddress_q_3_7 ;
    wire M_this_oam_ram_write_data_22;
    wire M_this_oam_ram_read_data_22;
    wire \this_ppu.un1_M_vaddress_q_3_6 ;
    wire M_this_oam_ram_write_data_31;
    wire N_52_0;
    wire M_this_oam_ram_write_data_16;
    wire N_158_0;
    wire M_this_oam_ram_read_data_21;
    wire M_this_oam_ram_read_data_20;
    wire \this_ppu.un1_M_vaddress_q_3_5 ;
    wire M_this_oam_ram_read_data_19;
    wire M_this_oam_ram_read_data_i_19;
    wire M_this_data_tmp_qZ0Z_16;
    wire M_this_data_tmp_qZ0Z_19;
    wire M_this_data_tmp_qZ0Z_18;
    wire M_this_data_tmp_qZ0Z_22;
    wire M_this_data_tmp_qZ0Z_17;
    wire N_54_0;
    wire N_1126_0;
    wire M_this_oam_ram_write_data_30;
    wire bfn_24_22_0_;
    wire un1_M_this_external_address_q_cry_0;
    wire un1_M_this_external_address_q_cry_1;
    wire un1_M_this_external_address_q_cry_2;
    wire un1_M_this_external_address_q_cry_3;
    wire un1_M_this_external_address_q_cry_4;
    wire un1_M_this_external_address_q_cry_5;
    wire un1_M_this_external_address_q_cry_6;
    wire un1_M_this_external_address_q_cry_7;
    wire bfn_24_23_0_;
    wire M_this_external_address_qZ0Z_9;
    wire un1_M_this_external_address_q_cry_8_c_RNI09PBZ0;
    wire un1_M_this_external_address_q_cry_8;
    wire un1_M_this_external_address_q_cry_9;
    wire un1_M_this_external_address_q_cry_10;
    wire un1_M_this_external_address_q_cry_11;
    wire un1_M_this_external_address_q_cry_12;
    wire un1_M_this_external_address_q_cry_13;
    wire un1_M_this_external_address_q_cry_14;
    wire M_this_sprites_address_qZ0Z_12;
    wire M_this_sprites_address_qZ0Z_11;
    wire M_this_sprites_address_qZ0Z_13;
    wire M_this_sprites_ram_write_en_0_0;
    wire \this_sprites_ram.mem_WE_2 ;
    wire M_this_oam_ram_write_data_8;
    wire M_this_data_tmp_qZ0Z_8;
    wire N_79_0;
    wire M_this_data_tmp_qZ0Z_0;
    wire N_43_0;
    wire N_77_0;
    wire M_this_data_tmp_qZ0Z_1;
    wire N_58_0;
    wire M_this_oam_ram_write_data_14;
    wire N_63_0;
    wire N_75_0;
    wire M_this_oam_ram_write_data_11;
    wire M_this_data_tmp_qZ0Z_11;
    wire M_this_data_tmp_qZ0Z_12;
    wire M_this_data_tmp_qZ0Z_9;
    wire M_this_data_tmp_qZ0Z_14;
    wire N_1134_0;
    wire N_39_0;
    wire M_this_oam_ram_write_data_27;
    wire M_this_data_tmp_qZ0Z_23;
    wire M_this_oam_ram_write_data_23;
    wire port_data_c_1;
    wire N_41_0;
    wire M_this_data_tmp_qZ0Z_2;
    wire un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0;
    wire port_data_c_3;
    wire M_this_external_address_qZ0Z_11;
    wire un1_M_this_external_address_q_cry_6_THRU_CO;
    wire M_this_external_address_qZ0Z_7;
    wire un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0;
    wire port_data_c_4;
    wire M_this_external_address_qZ0Z_12;
    wire un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0;
    wire M_this_external_address_qZ0Z_13;
    wire un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0;
    wire port_data_c_6;
    wire M_this_external_address_qZ0Z_14;
    wire un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0;
    wire port_data_c_0;
    wire M_this_external_address_qZ0Z_8;
    wire port_data_c_7;
    wire un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0;
    wire M_this_external_address_qZ0Z_15;
    wire un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0;
    wire port_data_c_2;
    wire M_this_external_address_qZ0Z_10;
    wire un1_M_this_state_q_11_0_i;
    wire M_this_external_address_qZ0Z_0;
    wire un1_M_this_external_address_q_cry_0_THRU_CO;
    wire M_this_external_address_qZ0Z_1;
    wire un1_M_this_external_address_q_cry_1_THRU_CO;
    wire M_this_external_address_qZ0Z_2;
    wire un1_M_this_external_address_q_cry_2_THRU_CO;
    wire M_this_external_address_qZ0Z_3;
    wire un1_M_this_external_address_q_cry_3_THRU_CO;
    wire M_this_external_address_qZ0Z_4;
    wire un1_M_this_external_address_q_cry_4_THRU_CO;
    wire M_this_external_address_qZ0Z_5;
    wire N_458_0;
    wire M_this_state_qZ0Z_4;
    wire un1_M_this_external_address_q_cry_5_THRU_CO;
    wire M_this_external_address_qZ0Z_6;
    wire M_this_oam_address_qZ0Z_1;
    wire N_156_0;
    wire M_this_oam_address_qZ0Z_0;
    wire N_69_0;
    wire port_data_c_5;
    wire M_this_data_tmp_qZ0Z_5;
    wire _gnd_net_;
    wire clk_0_c_g;
    wire N_1142_0;
    wire M_this_reset_cond_out_g_0;

    defparam \this_map_ram.mem_mem_0_0_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_0_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,M_this_map_ram_read_data_3,dangling_wire_2,dangling_wire_3,dangling_wire_4,M_this_map_ram_read_data_2,dangling_wire_5,dangling_wire_6,dangling_wire_7,M_this_map_ram_read_data_1,dangling_wire_8,dangling_wire_9,dangling_wire_10,M_this_map_ram_read_data_0,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__27777,N__27825,N__27870,N__29529,N__29577,N__25155,N__25212,N__25272,N__25335,N__25416}),
            .WADDR({dangling_wire_13,N__11496,N__11529,N__11559,N__11589,N__11268,N__11298,N__11328,N__11358,N__11388,N__11415}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__11469,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__13761,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__13752,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__15501,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__34586),
            .RE(N__17947),
            .WCLKE(N__18250),
            .WCLK(N__34587),
            .WE(N__17943));
    defparam \this_map_ram.mem_mem_0_1_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_1_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_42,dangling_wire_43,M_this_map_ram_read_data_7,dangling_wire_44,dangling_wire_45,dangling_wire_46,M_this_map_ram_read_data_6,dangling_wire_47,dangling_wire_48,dangling_wire_49,M_this_map_ram_read_data_5,dangling_wire_50,dangling_wire_51,dangling_wire_52,M_this_map_ram_read_data_4,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__27771,N__27819,N__27864,N__29523,N__29571,N__25149,N__25206,N__25265,N__25325,N__25409}),
            .WADDR({dangling_wire_55,N__11490,N__11523,N__11553,N__11583,N__11262,N__11292,N__11322,N__11352,N__11382,N__11409}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__16158,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__11463,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__11457,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__16170,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__34590),
            .RE(N__17948),
            .WCLKE(N__18261),
            .WCLK(N__34591),
            .WE(N__17989));
    defparam \this_oam_ram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_0_physical  (
            .RDATA({M_this_oam_ram_read_data_15,M_this_oam_ram_read_data_14,M_this_oam_ram_read_data_13,M_this_oam_ram_read_data_12,M_this_oam_ram_read_data_11,M_this_oam_ram_read_data_10,M_this_oam_ram_read_data_9,M_this_oam_ram_read_data_8,M_this_oam_ram_read_data_7,M_this_oam_ram_read_data_6,M_this_oam_ram_read_data_5,M_this_oam_ram_read_data_4,M_this_oam_ram_read_data_3,M_this_oam_ram_read_data_2,M_this_oam_ram_read_data_1,M_this_oam_ram_read_data_0}),
            .RADDR({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,N__23838,N__23469,N__23874,N__23427}),
            .WADDR({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,N__30717,N__30198,N__30639,N__30597}),
            .MASK({dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113}),
            .WDATA({N__29064,N__32052,N__28605,N__32058,N__32235,N__30234,N__32247,N__32115,N__28056,N__30723,N__34782,N__29226,N__30210,N__32241,N__32073,N__32100}),
            .RCLKE(),
            .RCLK(N__34546),
            .RE(N__17738),
            .WCLKE(N__31314),
            .WCLK(N__34547),
            .WE(N__17923));
    defparam \this_oam_ram.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,M_this_oam_ram_read_data_23,M_this_oam_ram_read_data_22,M_this_oam_ram_read_data_21,M_this_oam_ram_read_data_20,M_this_oam_ram_read_data_19,M_this_oam_ram_read_data_18,M_this_oam_ram_read_data_17,M_this_oam_ram_read_data_16}),
            .RADDR({dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__23832,N__23463,N__23868,N__23421}),
            .WADDR({dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,N__30711,N__30192,N__30631,N__30591}),
            .MASK({dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151}),
            .WDATA({N__31332,N__31578,N__20772,N__25965,N__32121,N__32127,N__32865,N__32085,N__32994,N__31380,N__30522,N__25980,N__30531,N__31326,N__31455,N__31320}),
            .RCLKE(),
            .RCLK(N__34564),
            .RE(N__17898),
            .WCLKE(N__31310),
            .WCLK(N__34565),
            .WE(N__17905));
    defparam \this_sprites_ram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,\this_sprites_ram.mem_out_bus0_1 ,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,\this_sprites_ram.mem_out_bus0_0 ,dangling_wire_163,dangling_wire_164,dangling_wire_165}),
            .RADDR({N__27154,N__13724,N__15127,N__17412,N__14489,N__28948,N__26996,N__29869,N__22800,N__25812,N__23346}),
            .WADDR({N__24879,N__22558,N__26613,N__21982,N__21360,N__21565,N__27633,N__24163,N__22265,N__26223,N__24468}),
            .MASK({dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181}),
            .WDATA({dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,N__27321,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,N__19652,dangling_wire_193,dangling_wire_194,dangling_wire_195}),
            .RCLKE(),
            .RCLK(N__34467),
            .RE(N__17992),
            .WCLKE(N__23085),
            .WCLK(N__34468),
            .WE(N__17922));
    defparam \this_sprites_ram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,\this_sprites_ram.mem_out_bus0_3 ,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,\this_sprites_ram.mem_out_bus0_2 ,dangling_wire_207,dangling_wire_208,dangling_wire_209}),
            .RADDR({N__27204,N__13717,N__15088,N__17407,N__14502,N__28878,N__26986,N__29862,N__22740,N__25808,N__23339}),
            .WADDR({N__24875,N__22559,N__26609,N__22008,N__21359,N__21564,N__27629,N__24164,N__22293,N__26222,N__24467}),
            .MASK({dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225}),
            .WDATA({dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,N__19980,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,N__23643,dangling_wire_237,dangling_wire_238,dangling_wire_239}),
            .RCLKE(),
            .RCLK(N__34469),
            .RE(N__17849),
            .WCLKE(N__23084),
            .WCLK(N__34470),
            .WE(N__17964));
    defparam \this_sprites_ram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,\this_sprites_ram.mem_out_bus1_1 ,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,\this_sprites_ram.mem_out_bus1_0 ,dangling_wire_251,dangling_wire_252,dangling_wire_253}),
            .RADDR({N__27196,N__13704,N__15132,N__17347,N__14496,N__28937,N__26985,N__29847,N__22794,N__25800,N__23338}),
            .WADDR({N__24874,N__22560,N__26608,N__22007,N__21352,N__21563,N__27622,N__24165,N__22289,N__26215,N__24460}),
            .MASK({dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269}),
            .WDATA({dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,N__27317,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,N__19653,dangling_wire_281,dangling_wire_282,dangling_wire_283}),
            .RCLKE(),
            .RCLK(N__34471),
            .RE(N__17959),
            .WCLKE(N__25092),
            .WCLK(N__34472),
            .WE(N__17963));
    defparam \this_sprites_ram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,\this_sprites_ram.mem_out_bus1_3 ,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,\this_sprites_ram.mem_out_bus1_2 ,dangling_wire_295,dangling_wire_296,dangling_wire_297}),
            .RADDR({N__27175,N__13695,N__15128,N__17392,N__14470,N__28920,N__26960,N__29814,N__22793,N__25784,N__23314}),
            .WADDR({N__24864,N__22561,N__26598,N__22024,N__21351,N__21566,N__27612,N__24166,N__22282,N__26214,N__24427}),
            .MASK({dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313}),
            .WDATA({dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,N__19976,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,N__23637,dangling_wire_325,dangling_wire_326,dangling_wire_327}),
            .RCLKE(),
            .RCLK(N__34481),
            .RE(N__17752),
            .WCLKE(N__25088),
            .WCLK(N__34480),
            .WE(N__17906));
    defparam \this_sprites_ram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,\this_sprites_ram.mem_out_bus2_1 ,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,\this_sprites_ram.mem_out_bus2_0 ,dangling_wire_339,dangling_wire_340,dangling_wire_341}),
            .RADDR({N__27144,N__13678,N__15118,N__17391,N__14495,N__28896,N__26946,N__29815,N__22775,N__25715,N__23313}),
            .WADDR({N__24825,N__22568,N__26584,N__22023,N__21338,N__21538,N__27599,N__24182,N__22253,N__26201,N__24450}),
            .MASK({dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,dangling_wire_357}),
            .WDATA({dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,N__27309,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,N__19651,dangling_wire_369,dangling_wire_370,dangling_wire_371}),
            .RCLKE(),
            .RCLK(N__34495),
            .RE(N__18019),
            .WCLKE(N__30357),
            .WCLK(N__34496),
            .WE(N__18010));
    defparam \this_sprites_ram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,\this_sprites_ram.mem_out_bus2_3 ,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,\this_sprites_ram.mem_out_bus2_2 ,dangling_wire_383,dangling_wire_384,dangling_wire_385}),
            .RADDR({N__27131,N__13601,N__15117,N__17358,N__14494,N__28850,N__26907,N__29798,N__22774,N__25757,N__23272}),
            .WADDR({N__24851,N__22571,N__26563,N__22032,N__21337,N__21537,N__27584,N__24178,N__22271,N__26200,N__24449}),
            .MASK({dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,dangling_wire_401}),
            .WDATA({dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,N__19938,dangling_wire_406,dangling_wire_407,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,N__23636,dangling_wire_413,dangling_wire_414,dangling_wire_415}),
            .RCLKE(),
            .RCLK(N__34511),
            .RE(N__17739),
            .WCLKE(N__30356),
            .WCLK(N__34512),
            .WE(N__18006));
    defparam \this_sprites_ram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,\this_sprites_ram.mem_out_bus3_1 ,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,\this_sprites_ram.mem_out_bus3_0 ,dangling_wire_427,dangling_wire_428,dangling_wire_429}),
            .RADDR({N__27080,N__13688,N__15093,N__17277,N__14460,N__28841,N__26859,N__29777,N__22741,N__25722,N__23271}),
            .WADDR({N__24850,N__22572,N__26535,N__22031,N__21318,N__21578,N__27568,N__24183,N__22228,N__26178,N__24433}),
            .MASK({dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,dangling_wire_445}),
            .WDATA({dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,N__27295,dangling_wire_450,dangling_wire_451,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,N__19643,dangling_wire_457,dangling_wire_458,dangling_wire_459}),
            .RCLKE(),
            .RCLK(N__34531),
            .RE(N__17957),
            .WCLKE(N__23114),
            .WCLK(N__34532),
            .WE(N__17934));
    defparam \this_sprites_ram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,\this_sprites_ram.mem_out_bus3_3 ,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,\this_sprites_ram.mem_out_bus3_2 ,dangling_wire_471,dangling_wire_472,dangling_wire_473}),
            .RADDR({N__27119,N__13631,N__15056,N__17348,N__14487,N__28930,N__26897,N__29870,N__22770,N__25794,N__23332}),
            .WADDR({N__24830,N__22569,N__26597,N__21972,N__21317,N__21572,N__27611,N__24176,N__22237,N__26199,N__24430}),
            .MASK({dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,dangling_wire_489}),
            .WDATA({dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,N__19974,dangling_wire_494,dangling_wire_495,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,N__23642,dangling_wire_501,dangling_wire_502,dangling_wire_503}),
            .RCLKE(),
            .RCLK(N__34522),
            .RE(N__17991),
            .WCLKE(N__23118),
            .WCLK(N__34523),
            .WE(N__17956));
    defparam \this_sprites_ram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,\this_sprites_ram.mem_out_bus4_1 ,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,dangling_wire_514,\this_sprites_ram.mem_out_bus4_0 ,dangling_wire_515,dangling_wire_516,dangling_wire_517}),
            .RADDR({N__27182,N__13671,N__15057,N__17384,N__14488,N__28944,N__26970,N__29883,N__22771,N__25807,N__23333}),
            .WADDR({N__24849,N__22552,N__26580,N__22000,N__21292,N__21576,N__27580,N__24159,N__22281,N__26198,N__24429}),
            .MASK({dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,dangling_wire_526,dangling_wire_527,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,dangling_wire_533}),
            .WDATA({dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,N__27316,dangling_wire_538,dangling_wire_539,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,N__19647,dangling_wire_545,dangling_wire_546,dangling_wire_547}),
            .RCLKE(),
            .RCLK(N__34553),
            .RE(N__17768),
            .WCLKE(N__23571),
            .WCLK(N__34554),
            .WE(N__17884));
    defparam \this_sprites_ram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,\this_sprites_ram.mem_out_bus4_3 ,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,dangling_wire_558,\this_sprites_ram.mem_out_bus4_2 ,dangling_wire_559,dangling_wire_560,dangling_wire_561}),
            .RADDR({N__27200,N__13700,N__15075,N__17405,N__14483,N__28949,N__26990,N__29875,N__22772,N__25780,N__23334}),
            .WADDR({N__24826,N__22553,N__26579,N__22022,N__21260,N__21577,N__27561,N__24177,N__22267,N__26197,N__24390}),
            .MASK({dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,dangling_wire_570,dangling_wire_571,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,dangling_wire_577}),
            .WDATA({dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,N__19967,dangling_wire_582,dangling_wire_583,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,N__23641,dangling_wire_589,dangling_wire_590,dangling_wire_591}),
            .RCLKE(),
            .RCLK(N__34571),
            .RE(N__17864),
            .WCLKE(N__23570),
            .WCLK(N__34572),
            .WE(N__17894));
    defparam \this_sprites_ram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,\this_sprites_ram.mem_out_bus5_1 ,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,dangling_wire_602,\this_sprites_ram.mem_out_bus5_0 ,dangling_wire_603,dangling_wire_604,dangling_wire_605}),
            .RADDR({N__27201,N__13716,N__15092,N__17406,N__14500,N__28950,N__26991,N__29882,N__22773,N__25799,N__23345}),
            .WADDR({N__24793,N__22478,N__26578,N__22021,N__21291,N__21579,N__27538,N__24130,N__22227,N__26196,N__24428}),
            .MASK({dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,dangling_wire_614,dangling_wire_615,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,dangling_wire_621}),
            .WDATA({dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,N__27305,dangling_wire_626,dangling_wire_627,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,N__19641,dangling_wire_633,dangling_wire_634,dangling_wire_635}),
            .RCLKE(),
            .RCLK(N__34578),
            .RE(N__17865),
            .WCLKE(N__26793),
            .WCLK(N__34579),
            .WE(N__17942));
    defparam \this_sprites_ram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,\this_sprites_ram.mem_out_bus5_3 ,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646,\this_sprites_ram.mem_out_bus5_2 ,dangling_wire_647,dangling_wire_648,dangling_wire_649}),
            .RADDR({N__27165,N__13711,N__15038,N__17399,N__14469,N__28851,N__26947,N__29808,N__22757,N__25740,N__23288}),
            .WADDR({N__24811,N__22570,N__26527,N__21955,N__21214,N__21550,N__27529,N__24133,N__22246,N__26147,N__24333}),
            .MASK({dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,dangling_wire_658,dangling_wire_659,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,dangling_wire_665}),
            .WDATA({dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,N__19948,dangling_wire_670,dangling_wire_671,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,N__23618,dangling_wire_677,dangling_wire_678,dangling_wire_679}),
            .RCLKE(),
            .RCLK(N__34573),
            .RE(N__17765),
            .WCLKE(N__26786),
            .WCLK(N__34574),
            .WE(N__17968));
    defparam \this_sprites_ram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,\this_sprites_ram.mem_out_bus6_1 ,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,\this_sprites_ram.mem_out_bus6_0 ,dangling_wire_691,dangling_wire_692,dangling_wire_693}),
            .RADDR({N__27189,N__13696,N__15106,N__17400,N__14501,N__28888,N__26977,N__29822,N__22785,N__25741,N__23324}),
            .WADDR({N__24740,N__22442,N__26491,N__21931,N__21270,N__21570,N__27493,N__24098,N__22185,N__26139,N__24403}),
            .MASK({dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,dangling_wire_702,dangling_wire_703,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,dangling_wire_709}),
            .WDATA({dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713,N__27263,dangling_wire_714,dangling_wire_715,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,N__19640,dangling_wire_721,dangling_wire_722,dangling_wire_723}),
            .RCLKE(),
            .RCLK(N__34582),
            .RE(N__17958),
            .WCLKE(N__31592),
            .WCLK(N__34583),
            .WE(N__17996));
    defparam \this_sprites_ram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_724,dangling_wire_725,dangling_wire_726,dangling_wire_727,\this_sprites_ram.mem_out_bus6_3 ,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,\this_sprites_ram.mem_out_bus6_2 ,dangling_wire_735,dangling_wire_736,dangling_wire_737}),
            .RADDR({N__27202,N__13670,N__15107,N__17401,N__14464,N__28889,N__26978,N__29858,N__22786,N__25775,N__23325}),
            .WADDR({N__24806,N__22554,N__26528,N__21927,N__21271,N__21571,N__27522,N__24132,N__22241,N__26140,N__24404}),
            .MASK({dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741,dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,dangling_wire_753}),
            .WDATA({dangling_wire_754,dangling_wire_755,dangling_wire_756,dangling_wire_757,N__19944,dangling_wire_758,dangling_wire_759,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,N__23619,dangling_wire_765,dangling_wire_766,dangling_wire_767}),
            .RCLKE(),
            .RCLK(N__34588),
            .RE(N__17766),
            .WCLKE(N__31593),
            .WCLK(N__34589),
            .WE(N__17997));
    defparam \this_sprites_ram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_768,dangling_wire_769,dangling_wire_770,dangling_wire_771,\this_sprites_ram.mem_out_bus7_1 ,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,dangling_wire_778,\this_sprites_ram.mem_out_bus7_0 ,dangling_wire_779,dangling_wire_780,dangling_wire_781}),
            .RADDR({N__27164,N__13715,N__15125,N__17380,N__14465,N__28918,N__26992,N__29851,N__22798,N__25776,N__23343}),
            .WADDR({N__24807,N__22520,N__26561,N__21932,N__21296,N__21548,N__27548,N__24131,N__22242,N__26176,N__24431}),
            .MASK({dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785,dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,dangling_wire_797}),
            .WDATA({dangling_wire_798,dangling_wire_799,dangling_wire_800,dangling_wire_801,N__27264,dangling_wire_802,dangling_wire_803,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,N__19642,dangling_wire_809,dangling_wire_810,dangling_wire_811}),
            .RCLKE(),
            .RCLK(N__34593),
            .RE(N__18012),
            .WCLKE(N__28313),
            .WCLK(N__34594),
            .WE(N__18020));
    defparam \this_sprites_ram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_812,dangling_wire_813,dangling_wire_814,dangling_wire_815,\this_sprites_ram.mem_out_bus7_3 ,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,dangling_wire_822,\this_sprites_ram.mem_out_bus7_2 ,dangling_wire_823,dangling_wire_824,dangling_wire_825}),
            .RADDR({N__27203,N__13725,N__15126,N__17411,N__14490,N__28919,N__26997,N__29874,N__22799,N__25798,N__23344}),
            .WADDR({N__24831,N__22548,N__26562,N__21954,N__21297,N__21549,N__27549,N__24155,N__22266,N__26177,N__24432}),
            .MASK({dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829,dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,dangling_wire_834,dangling_wire_835,dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,dangling_wire_840,dangling_wire_841}),
            .WDATA({dangling_wire_842,dangling_wire_843,dangling_wire_844,dangling_wire_845,N__19975,dangling_wire_846,dangling_wire_847,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,N__23629,dangling_wire_853,dangling_wire_854,dangling_wire_855}),
            .RCLKE(),
            .RCLK(N__34595),
            .RE(N__17767),
            .WCLKE(N__28314),
            .WCLK(N__34596),
            .WE(N__18021));
    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_856,dangling_wire_857,dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,dangling_wire_867,M_this_vram_read_data_3,M_this_vram_read_data_2,M_this_vram_read_data_1,M_this_vram_read_data_0}),
            .RADDR({dangling_wire_868,dangling_wire_869,dangling_wire_870,N__11079,N__11106,N__13428,N__11094,N__13194,N__11115,N__13104,N__12225}),
            .WADDR({dangling_wire_871,dangling_wire_872,dangling_wire_873,N__29337,N__25202,N__25268,N__25334,N__25412,N__25476,N__25533,N__25590}),
            .MASK({dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,dangling_wire_884,dangling_wire_885,dangling_wire_886,dangling_wire_887,dangling_wire_888,dangling_wire_889}),
            .WDATA({dangling_wire_890,dangling_wire_891,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,dangling_wire_899,dangling_wire_900,dangling_wire_901,N__20739,N__20721,N__21786,N__20694}),
            .RCLKE(),
            .RCLK(N__34539),
            .RE(N__17803),
            .WCLKE(N__22614),
            .WCLK(N__34540),
            .WE(N__17952));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__36349),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__36351),
            .DIN(N__36350),
            .DOUT(N__36349),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__36351),
            .PADOUT(N__36350),
            .PADIN(N__36349),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__36340),
            .DIN(N__36339),
            .DOUT(N__36338),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__36340),
            .PADOUT(N__36339),
            .PADIN(N__36338),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__36331),
            .DIN(N__36330),
            .DOUT(N__36329),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__36331),
            .PADOUT(N__36330),
            .PADIN(N__36329),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__36322),
            .DIN(N__36321),
            .DOUT(N__36320),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__36322),
            .PADOUT(N__36321),
            .PADIN(N__36320),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11760),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__36313),
            .DIN(N__36312),
            .DOUT(N__36311),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__36313),
            .PADOUT(N__36312),
            .PADIN(N__36311),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14541),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_0_iopad (
            .OE(N__36304),
            .DIN(N__36303),
            .DOUT(N__36302),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__36304),
            .PADOUT(N__36303),
            .PADIN(N__36302),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__18011),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_1_iopad (
            .OE(N__36295),
            .DIN(N__36294),
            .DOUT(N__36293),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__36295),
            .PADOUT(N__36294),
            .PADIN(N__36293),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21699),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_2_iopad (
            .OE(N__36286),
            .DIN(N__36285),
            .DOUT(N__36284),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__36286),
            .PADOUT(N__36285),
            .PADIN(N__36284),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_3_iopad (
            .OE(N__36277),
            .DIN(N__36276),
            .DOUT(N__36275),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__36277),
            .PADOUT(N__36276),
            .PADIN(N__36275),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_4_iopad (
            .OE(N__36268),
            .DIN(N__36267),
            .DOUT(N__36266),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__36268),
            .PADOUT(N__36267),
            .PADIN(N__36266),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_5_iopad (
            .OE(N__36259),
            .DIN(N__36258),
            .DOUT(N__36257),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__36259),
            .PADOUT(N__36258),
            .PADIN(N__36257),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_6_iopad (
            .OE(N__36250),
            .DIN(N__36249),
            .DOUT(N__36248),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__36250),
            .PADOUT(N__36249),
            .PADIN(N__36248),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_7_iopad (
            .OE(N__36241),
            .DIN(N__36240),
            .DOUT(N__36239),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__36241),
            .PADOUT(N__36240),
            .PADIN(N__36239),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__36232),
            .DIN(N__36231),
            .DOUT(N__36230),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__36232),
            .PADOUT(N__36231),
            .PADIN(N__36230),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__33279),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16000));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__36223),
            .DIN(N__36222),
            .DOUT(N__36221),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__36223),
            .PADOUT(N__36222),
            .PADIN(N__36221),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__33221),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15989));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__36214),
            .DIN(N__36213),
            .DOUT(N__36212),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__36214),
            .PADOUT(N__36213),
            .PADIN(N__36212),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__33180),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16056));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__36205),
            .DIN(N__36204),
            .DOUT(N__36203),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__36205),
            .PADOUT(N__36204),
            .PADIN(N__36203),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__33132),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16096));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__36196),
            .DIN(N__36195),
            .DOUT(N__36194),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__36196),
            .PADOUT(N__36195),
            .PADIN(N__36194),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__33083),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16083));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__36187),
            .DIN(N__36186),
            .DOUT(N__36185),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__36187),
            .PADOUT(N__36186),
            .PADIN(N__36185),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__33042),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16061));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__36178),
            .DIN(N__36177),
            .DOUT(N__36176),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__36178),
            .PADOUT(N__36177),
            .PADIN(N__36176),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__35526),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16097));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__36169),
            .DIN(N__36168),
            .DOUT(N__36167),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__36169),
            .PADOUT(N__36168),
            .PADIN(N__36167),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__32652),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16094));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__36160),
            .DIN(N__36159),
            .DOUT(N__36158),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__36160),
            .PADOUT(N__36159),
            .PADIN(N__36158),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__33330),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16027));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__36151),
            .DIN(N__36150),
            .DOUT(N__36149),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__36151),
            .PADOUT(N__36150),
            .PADIN(N__36149),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__32691),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16095));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__36142),
            .DIN(N__36141),
            .DOUT(N__36140),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__36142),
            .PADOUT(N__36141),
            .PADIN(N__36140),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__32481),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16084));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__36133),
            .DIN(N__36132),
            .DOUT(N__36131),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__36133),
            .PADOUT(N__36132),
            .PADIN(N__36131),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__32445),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16062));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__36124),
            .DIN(N__36123),
            .DOUT(N__36122),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__36124),
            .PADOUT(N__36123),
            .PADIN(N__36122),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__32277),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16098));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__36115),
            .DIN(N__36114),
            .DOUT(N__36113),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__36115),
            .PADOUT(N__36114),
            .PADIN(N__36113),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__33534),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16022));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__36106),
            .DIN(N__36105),
            .DOUT(N__36104),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__36106),
            .PADOUT(N__36105),
            .PADIN(N__36104),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__33696),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15999));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__36097),
            .DIN(N__36096),
            .DOUT(N__36095),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__36097),
            .PADOUT(N__36096),
            .PADIN(N__36095),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__32043),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16057));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__36088),
            .DIN(N__36087),
            .DOUT(N__36086),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__36088),
            .PADOUT(N__36087),
            .PADIN(N__36086),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__36079),
            .DIN(N__36078),
            .DOUT(N__36077),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__36079),
            .PADOUT(N__36078),
            .PADIN(N__36077),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__36070),
            .DIN(N__36069),
            .DOUT(N__36068),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__36070),
            .PADOUT(N__36069),
            .PADIN(N__36068),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__36061),
            .DIN(N__36060),
            .DOUT(N__36059),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__36061),
            .PADOUT(N__36060),
            .PADIN(N__36059),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__36052),
            .DIN(N__36051),
            .DOUT(N__36050),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__36052),
            .PADOUT(N__36051),
            .PADIN(N__36050),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__36043),
            .DIN(N__36042),
            .DOUT(N__36041),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__36043),
            .PADOUT(N__36042),
            .PADIN(N__36041),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__36034),
            .DIN(N__36033),
            .DOUT(N__36032),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__36034),
            .PADOUT(N__36033),
            .PADIN(N__36032),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__36025),
            .DIN(N__36024),
            .DOUT(N__36023),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__36025),
            .PADOUT(N__36024),
            .PADIN(N__36023),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_7_iopad (
            .OE(N__36016),
            .DIN(N__36015),
            .DOUT(N__36014),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_7_preio (
            .PADOEN(N__36016),
            .PADOUT(N__36015),
            .PADIN(N__36014),
            .CLOCKENABLE(),
            .DIN0(port_data_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__36007),
            .DIN(N__36006),
            .DOUT(N__36005),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__36007),
            .PADOUT(N__36006),
            .PADIN(N__36005),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11058),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__35998),
            .DIN(N__35997),
            .DOUT(N__35996),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__35998),
            .PADOUT(N__35997),
            .PADIN(N__35996),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22941),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__35989),
            .DIN(N__35988),
            .DOUT(N__35987),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__35989),
            .PADOUT(N__35988),
            .PADIN(N__35987),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__35980),
            .DIN(N__35979),
            .DOUT(N__35978),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__35980),
            .PADOUT(N__35979),
            .PADIN(N__35978),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11052),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__35971),
            .DIN(N__35970),
            .DOUT(N__35969),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__35971),
            .PADOUT(N__35970),
            .PADIN(N__35969),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__17990),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__16026));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__35962),
            .DIN(N__35961),
            .DOUT(N__35960),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__35962),
            .PADOUT(N__35961),
            .PADIN(N__35960),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11139),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__35953),
            .DIN(N__35952),
            .DOUT(N__35951),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__35953),
            .PADOUT(N__35952),
            .PADIN(N__35951),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11124),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__35944),
            .DIN(N__35943),
            .DOUT(N__35942),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__35944),
            .PADOUT(N__35943),
            .PADIN(N__35942),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__15693),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__35935),
            .DIN(N__35934),
            .DOUT(N__35933),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__35935),
            .PADOUT(N__35934),
            .PADIN(N__35933),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__15522),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__35926),
            .DIN(N__35925),
            .DOUT(N__35924),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__35926),
            .PADOUT(N__35925),
            .PADIN(N__35924),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12309),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__35917),
            .DIN(N__35916),
            .DOUT(N__35915),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__35917),
            .PADOUT(N__35916),
            .PADIN(N__35915),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__15750),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__35908),
            .DIN(N__35907),
            .DOUT(N__35906),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__35908),
            .PADOUT(N__35907),
            .PADIN(N__35906),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__35899),
            .DIN(N__35898),
            .DOUT(N__35897),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__35899),
            .PADOUT(N__35898),
            .PADIN(N__35897),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11037),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__35890),
            .DIN(N__35889),
            .DOUT(N__35888),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__35890),
            .PADOUT(N__35889),
            .PADIN(N__35888),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11235),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__9096 (
            .O(N__35871),
            .I(N__35868));
    InMux I__9095 (
            .O(N__35868),
            .I(N__35847));
    InMux I__9094 (
            .O(N__35867),
            .I(N__35829));
    InMux I__9093 (
            .O(N__35866),
            .I(N__35829));
    InMux I__9092 (
            .O(N__35865),
            .I(N__35829));
    InMux I__9091 (
            .O(N__35864),
            .I(N__35829));
    InMux I__9090 (
            .O(N__35863),
            .I(N__35829));
    InMux I__9089 (
            .O(N__35862),
            .I(N__35829));
    InMux I__9088 (
            .O(N__35861),
            .I(N__35829));
    InMux I__9087 (
            .O(N__35860),
            .I(N__35829));
    InMux I__9086 (
            .O(N__35859),
            .I(N__35814));
    InMux I__9085 (
            .O(N__35858),
            .I(N__35814));
    InMux I__9084 (
            .O(N__35857),
            .I(N__35814));
    InMux I__9083 (
            .O(N__35856),
            .I(N__35814));
    InMux I__9082 (
            .O(N__35855),
            .I(N__35814));
    InMux I__9081 (
            .O(N__35854),
            .I(N__35814));
    InMux I__9080 (
            .O(N__35853),
            .I(N__35814));
    InMux I__9079 (
            .O(N__35852),
            .I(N__35806));
    InMux I__9078 (
            .O(N__35851),
            .I(N__35803));
    InMux I__9077 (
            .O(N__35850),
            .I(N__35800));
    LocalMux I__9076 (
            .O(N__35847),
            .I(N__35797));
    InMux I__9075 (
            .O(N__35846),
            .I(N__35794));
    LocalMux I__9074 (
            .O(N__35829),
            .I(N__35788));
    LocalMux I__9073 (
            .O(N__35814),
            .I(N__35788));
    InMux I__9072 (
            .O(N__35813),
            .I(N__35775));
    InMux I__9071 (
            .O(N__35812),
            .I(N__35766));
    InMux I__9070 (
            .O(N__35811),
            .I(N__35766));
    InMux I__9069 (
            .O(N__35810),
            .I(N__35766));
    InMux I__9068 (
            .O(N__35809),
            .I(N__35766));
    LocalMux I__9067 (
            .O(N__35806),
            .I(N__35756));
    LocalMux I__9066 (
            .O(N__35803),
            .I(N__35756));
    LocalMux I__9065 (
            .O(N__35800),
            .I(N__35756));
    Span4Mux_v I__9064 (
            .O(N__35797),
            .I(N__35750));
    LocalMux I__9063 (
            .O(N__35794),
            .I(N__35750));
    InMux I__9062 (
            .O(N__35793),
            .I(N__35747));
    Span4Mux_v I__9061 (
            .O(N__35788),
            .I(N__35744));
    InMux I__9060 (
            .O(N__35787),
            .I(N__35741));
    InMux I__9059 (
            .O(N__35786),
            .I(N__35738));
    InMux I__9058 (
            .O(N__35785),
            .I(N__35731));
    InMux I__9057 (
            .O(N__35784),
            .I(N__35731));
    InMux I__9056 (
            .O(N__35783),
            .I(N__35731));
    InMux I__9055 (
            .O(N__35782),
            .I(N__35728));
    InMux I__9054 (
            .O(N__35781),
            .I(N__35725));
    InMux I__9053 (
            .O(N__35780),
            .I(N__35718));
    InMux I__9052 (
            .O(N__35779),
            .I(N__35718));
    InMux I__9051 (
            .O(N__35778),
            .I(N__35718));
    LocalMux I__9050 (
            .O(N__35775),
            .I(N__35708));
    LocalMux I__9049 (
            .O(N__35766),
            .I(N__35708));
    InMux I__9048 (
            .O(N__35765),
            .I(N__35701));
    InMux I__9047 (
            .O(N__35764),
            .I(N__35701));
    InMux I__9046 (
            .O(N__35763),
            .I(N__35701));
    Span4Mux_v I__9045 (
            .O(N__35756),
            .I(N__35698));
    InMux I__9044 (
            .O(N__35755),
            .I(N__35695));
    Span4Mux_h I__9043 (
            .O(N__35750),
            .I(N__35692));
    LocalMux I__9042 (
            .O(N__35747),
            .I(N__35689));
    Sp12to4 I__9041 (
            .O(N__35744),
            .I(N__35680));
    LocalMux I__9040 (
            .O(N__35741),
            .I(N__35680));
    LocalMux I__9039 (
            .O(N__35738),
            .I(N__35680));
    LocalMux I__9038 (
            .O(N__35731),
            .I(N__35680));
    LocalMux I__9037 (
            .O(N__35728),
            .I(N__35673));
    LocalMux I__9036 (
            .O(N__35725),
            .I(N__35673));
    LocalMux I__9035 (
            .O(N__35718),
            .I(N__35673));
    InMux I__9034 (
            .O(N__35717),
            .I(N__35666));
    InMux I__9033 (
            .O(N__35716),
            .I(N__35666));
    InMux I__9032 (
            .O(N__35715),
            .I(N__35666));
    InMux I__9031 (
            .O(N__35714),
            .I(N__35661));
    InMux I__9030 (
            .O(N__35713),
            .I(N__35661));
    Odrv4 I__9029 (
            .O(N__35708),
            .I(N_458_0));
    LocalMux I__9028 (
            .O(N__35701),
            .I(N_458_0));
    Odrv4 I__9027 (
            .O(N__35698),
            .I(N_458_0));
    LocalMux I__9026 (
            .O(N__35695),
            .I(N_458_0));
    Odrv4 I__9025 (
            .O(N__35692),
            .I(N_458_0));
    Odrv4 I__9024 (
            .O(N__35689),
            .I(N_458_0));
    Odrv12 I__9023 (
            .O(N__35680),
            .I(N_458_0));
    Odrv4 I__9022 (
            .O(N__35673),
            .I(N_458_0));
    LocalMux I__9021 (
            .O(N__35666),
            .I(N_458_0));
    LocalMux I__9020 (
            .O(N__35661),
            .I(N_458_0));
    InMux I__9019 (
            .O(N__35640),
            .I(N__35619));
    InMux I__9018 (
            .O(N__35639),
            .I(N__35619));
    InMux I__9017 (
            .O(N__35638),
            .I(N__35619));
    InMux I__9016 (
            .O(N__35637),
            .I(N__35619));
    InMux I__9015 (
            .O(N__35636),
            .I(N__35619));
    InMux I__9014 (
            .O(N__35635),
            .I(N__35619));
    InMux I__9013 (
            .O(N__35634),
            .I(N__35619));
    LocalMux I__9012 (
            .O(N__35619),
            .I(N__35606));
    InMux I__9011 (
            .O(N__35618),
            .I(N__35589));
    InMux I__9010 (
            .O(N__35617),
            .I(N__35589));
    InMux I__9009 (
            .O(N__35616),
            .I(N__35589));
    InMux I__9008 (
            .O(N__35615),
            .I(N__35589));
    InMux I__9007 (
            .O(N__35614),
            .I(N__35589));
    InMux I__9006 (
            .O(N__35613),
            .I(N__35589));
    InMux I__9005 (
            .O(N__35612),
            .I(N__35589));
    InMux I__9004 (
            .O(N__35611),
            .I(N__35589));
    InMux I__9003 (
            .O(N__35610),
            .I(N__35586));
    CascadeMux I__9002 (
            .O(N__35609),
            .I(N__35583));
    Span4Mux_v I__9001 (
            .O(N__35606),
            .I(N__35580));
    LocalMux I__9000 (
            .O(N__35589),
            .I(N__35573));
    LocalMux I__8999 (
            .O(N__35586),
            .I(N__35573));
    InMux I__8998 (
            .O(N__35583),
            .I(N__35570));
    Span4Mux_h I__8997 (
            .O(N__35580),
            .I(N__35567));
    InMux I__8996 (
            .O(N__35579),
            .I(N__35564));
    InMux I__8995 (
            .O(N__35578),
            .I(N__35561));
    Span12Mux_h I__8994 (
            .O(N__35573),
            .I(N__35558));
    LocalMux I__8993 (
            .O(N__35570),
            .I(N__35555));
    Span4Mux_h I__8992 (
            .O(N__35567),
            .I(N__35552));
    LocalMux I__8991 (
            .O(N__35564),
            .I(N__35549));
    LocalMux I__8990 (
            .O(N__35561),
            .I(M_this_state_qZ0Z_4));
    Odrv12 I__8989 (
            .O(N__35558),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__8988 (
            .O(N__35555),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__8987 (
            .O(N__35552),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__8986 (
            .O(N__35549),
            .I(M_this_state_qZ0Z_4));
    InMux I__8985 (
            .O(N__35538),
            .I(N__35535));
    LocalMux I__8984 (
            .O(N__35535),
            .I(N__35532));
    Span4Mux_h I__8983 (
            .O(N__35532),
            .I(N__35529));
    Odrv4 I__8982 (
            .O(N__35529),
            .I(un1_M_this_external_address_q_cry_5_THRU_CO));
    IoInMux I__8981 (
            .O(N__35526),
            .I(N__35523));
    LocalMux I__8980 (
            .O(N__35523),
            .I(N__35520));
    IoSpan4Mux I__8979 (
            .O(N__35520),
            .I(N__35516));
    InMux I__8978 (
            .O(N__35519),
            .I(N__35512));
    IoSpan4Mux I__8977 (
            .O(N__35516),
            .I(N__35509));
    CascadeMux I__8976 (
            .O(N__35515),
            .I(N__35506));
    LocalMux I__8975 (
            .O(N__35512),
            .I(N__35503));
    Span4Mux_s3_h I__8974 (
            .O(N__35509),
            .I(N__35500));
    InMux I__8973 (
            .O(N__35506),
            .I(N__35497));
    Span4Mux_h I__8972 (
            .O(N__35503),
            .I(N__35494));
    Odrv4 I__8971 (
            .O(N__35500),
            .I(M_this_external_address_qZ0Z_6));
    LocalMux I__8970 (
            .O(N__35497),
            .I(M_this_external_address_qZ0Z_6));
    Odrv4 I__8969 (
            .O(N__35494),
            .I(M_this_external_address_qZ0Z_6));
    InMux I__8968 (
            .O(N__35487),
            .I(N__35470));
    InMux I__8967 (
            .O(N__35486),
            .I(N__35470));
    InMux I__8966 (
            .O(N__35485),
            .I(N__35470));
    InMux I__8965 (
            .O(N__35484),
            .I(N__35470));
    InMux I__8964 (
            .O(N__35483),
            .I(N__35463));
    InMux I__8963 (
            .O(N__35482),
            .I(N__35460));
    InMux I__8962 (
            .O(N__35481),
            .I(N__35453));
    InMux I__8961 (
            .O(N__35480),
            .I(N__35453));
    InMux I__8960 (
            .O(N__35479),
            .I(N__35453));
    LocalMux I__8959 (
            .O(N__35470),
            .I(N__35449));
    CascadeMux I__8958 (
            .O(N__35469),
            .I(N__35446));
    InMux I__8957 (
            .O(N__35468),
            .I(N__35436));
    CascadeMux I__8956 (
            .O(N__35467),
            .I(N__35432));
    InMux I__8955 (
            .O(N__35466),
            .I(N__35424));
    LocalMux I__8954 (
            .O(N__35463),
            .I(N__35415));
    LocalMux I__8953 (
            .O(N__35460),
            .I(N__35410));
    LocalMux I__8952 (
            .O(N__35453),
            .I(N__35410));
    InMux I__8951 (
            .O(N__35452),
            .I(N__35407));
    Span4Mux_h I__8950 (
            .O(N__35449),
            .I(N__35404));
    InMux I__8949 (
            .O(N__35446),
            .I(N__35401));
    InMux I__8948 (
            .O(N__35445),
            .I(N__35392));
    InMux I__8947 (
            .O(N__35444),
            .I(N__35392));
    InMux I__8946 (
            .O(N__35443),
            .I(N__35383));
    InMux I__8945 (
            .O(N__35442),
            .I(N__35383));
    InMux I__8944 (
            .O(N__35441),
            .I(N__35383));
    InMux I__8943 (
            .O(N__35440),
            .I(N__35383));
    InMux I__8942 (
            .O(N__35439),
            .I(N__35380));
    LocalMux I__8941 (
            .O(N__35436),
            .I(N__35377));
    InMux I__8940 (
            .O(N__35435),
            .I(N__35372));
    InMux I__8939 (
            .O(N__35432),
            .I(N__35372));
    InMux I__8938 (
            .O(N__35431),
            .I(N__35369));
    InMux I__8937 (
            .O(N__35430),
            .I(N__35366));
    InMux I__8936 (
            .O(N__35429),
            .I(N__35359));
    InMux I__8935 (
            .O(N__35428),
            .I(N__35359));
    InMux I__8934 (
            .O(N__35427),
            .I(N__35359));
    LocalMux I__8933 (
            .O(N__35424),
            .I(N__35356));
    InMux I__8932 (
            .O(N__35423),
            .I(N__35345));
    InMux I__8931 (
            .O(N__35422),
            .I(N__35345));
    InMux I__8930 (
            .O(N__35421),
            .I(N__35345));
    InMux I__8929 (
            .O(N__35420),
            .I(N__35345));
    InMux I__8928 (
            .O(N__35419),
            .I(N__35345));
    CascadeMux I__8927 (
            .O(N__35418),
            .I(N__35342));
    Span4Mux_h I__8926 (
            .O(N__35415),
            .I(N__35337));
    Span4Mux_h I__8925 (
            .O(N__35410),
            .I(N__35334));
    LocalMux I__8924 (
            .O(N__35407),
            .I(N__35327));
    Span4Mux_v I__8923 (
            .O(N__35404),
            .I(N__35327));
    LocalMux I__8922 (
            .O(N__35401),
            .I(N__35327));
    InMux I__8921 (
            .O(N__35400),
            .I(N__35324));
    InMux I__8920 (
            .O(N__35399),
            .I(N__35321));
    InMux I__8919 (
            .O(N__35398),
            .I(N__35316));
    InMux I__8918 (
            .O(N__35397),
            .I(N__35316));
    LocalMux I__8917 (
            .O(N__35392),
            .I(N__35313));
    LocalMux I__8916 (
            .O(N__35383),
            .I(N__35306));
    LocalMux I__8915 (
            .O(N__35380),
            .I(N__35306));
    Span4Mux_v I__8914 (
            .O(N__35377),
            .I(N__35306));
    LocalMux I__8913 (
            .O(N__35372),
            .I(N__35303));
    LocalMux I__8912 (
            .O(N__35369),
            .I(N__35292));
    LocalMux I__8911 (
            .O(N__35366),
            .I(N__35292));
    LocalMux I__8910 (
            .O(N__35359),
            .I(N__35292));
    Span4Mux_v I__8909 (
            .O(N__35356),
            .I(N__35292));
    LocalMux I__8908 (
            .O(N__35345),
            .I(N__35292));
    InMux I__8907 (
            .O(N__35342),
            .I(N__35289));
    InMux I__8906 (
            .O(N__35341),
            .I(N__35284));
    InMux I__8905 (
            .O(N__35340),
            .I(N__35284));
    Span4Mux_h I__8904 (
            .O(N__35337),
            .I(N__35279));
    Span4Mux_h I__8903 (
            .O(N__35334),
            .I(N__35279));
    Span4Mux_h I__8902 (
            .O(N__35327),
            .I(N__35274));
    LocalMux I__8901 (
            .O(N__35324),
            .I(N__35274));
    LocalMux I__8900 (
            .O(N__35321),
            .I(N__35261));
    LocalMux I__8899 (
            .O(N__35316),
            .I(N__35261));
    Span4Mux_v I__8898 (
            .O(N__35313),
            .I(N__35261));
    Span4Mux_h I__8897 (
            .O(N__35306),
            .I(N__35261));
    Span4Mux_v I__8896 (
            .O(N__35303),
            .I(N__35261));
    Span4Mux_v I__8895 (
            .O(N__35292),
            .I(N__35261));
    LocalMux I__8894 (
            .O(N__35289),
            .I(M_this_oam_address_qZ0Z_1));
    LocalMux I__8893 (
            .O(N__35284),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__8892 (
            .O(N__35279),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__8891 (
            .O(N__35274),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__8890 (
            .O(N__35261),
            .I(M_this_oam_address_qZ0Z_1));
    CascadeMux I__8889 (
            .O(N__35250),
            .I(N__35243));
    CascadeMux I__8888 (
            .O(N__35249),
            .I(N__35240));
    CascadeMux I__8887 (
            .O(N__35248),
            .I(N__35225));
    InMux I__8886 (
            .O(N__35247),
            .I(N__35222));
    InMux I__8885 (
            .O(N__35246),
            .I(N__35213));
    InMux I__8884 (
            .O(N__35243),
            .I(N__35213));
    InMux I__8883 (
            .O(N__35240),
            .I(N__35213));
    InMux I__8882 (
            .O(N__35239),
            .I(N__35213));
    InMux I__8881 (
            .O(N__35238),
            .I(N__35210));
    InMux I__8880 (
            .O(N__35237),
            .I(N__35201));
    InMux I__8879 (
            .O(N__35236),
            .I(N__35201));
    InMux I__8878 (
            .O(N__35235),
            .I(N__35201));
    InMux I__8877 (
            .O(N__35234),
            .I(N__35201));
    CascadeMux I__8876 (
            .O(N__35233),
            .I(N__35197));
    CascadeMux I__8875 (
            .O(N__35232),
            .I(N__35194));
    CascadeMux I__8874 (
            .O(N__35231),
            .I(N__35191));
    InMux I__8873 (
            .O(N__35230),
            .I(N__35180));
    CascadeMux I__8872 (
            .O(N__35229),
            .I(N__35177));
    CascadeMux I__8871 (
            .O(N__35228),
            .I(N__35171));
    InMux I__8870 (
            .O(N__35225),
            .I(N__35166));
    LocalMux I__8869 (
            .O(N__35222),
            .I(N__35159));
    LocalMux I__8868 (
            .O(N__35213),
            .I(N__35159));
    LocalMux I__8867 (
            .O(N__35210),
            .I(N__35156));
    LocalMux I__8866 (
            .O(N__35201),
            .I(N__35153));
    InMux I__8865 (
            .O(N__35200),
            .I(N__35142));
    InMux I__8864 (
            .O(N__35197),
            .I(N__35142));
    InMux I__8863 (
            .O(N__35194),
            .I(N__35142));
    InMux I__8862 (
            .O(N__35191),
            .I(N__35142));
    InMux I__8861 (
            .O(N__35190),
            .I(N__35142));
    InMux I__8860 (
            .O(N__35189),
            .I(N__35139));
    InMux I__8859 (
            .O(N__35188),
            .I(N__35136));
    InMux I__8858 (
            .O(N__35187),
            .I(N__35129));
    InMux I__8857 (
            .O(N__35186),
            .I(N__35129));
    InMux I__8856 (
            .O(N__35185),
            .I(N__35129));
    InMux I__8855 (
            .O(N__35184),
            .I(N__35126));
    CascadeMux I__8854 (
            .O(N__35183),
            .I(N__35123));
    LocalMux I__8853 (
            .O(N__35180),
            .I(N__35116));
    InMux I__8852 (
            .O(N__35177),
            .I(N__35111));
    InMux I__8851 (
            .O(N__35176),
            .I(N__35111));
    InMux I__8850 (
            .O(N__35175),
            .I(N__35106));
    InMux I__8849 (
            .O(N__35174),
            .I(N__35106));
    InMux I__8848 (
            .O(N__35171),
            .I(N__35099));
    InMux I__8847 (
            .O(N__35170),
            .I(N__35099));
    InMux I__8846 (
            .O(N__35169),
            .I(N__35099));
    LocalMux I__8845 (
            .O(N__35166),
            .I(N__35095));
    InMux I__8844 (
            .O(N__35165),
            .I(N__35090));
    InMux I__8843 (
            .O(N__35164),
            .I(N__35090));
    Span4Mux_v I__8842 (
            .O(N__35159),
            .I(N__35081));
    Span4Mux_h I__8841 (
            .O(N__35156),
            .I(N__35081));
    Span4Mux_v I__8840 (
            .O(N__35153),
            .I(N__35081));
    LocalMux I__8839 (
            .O(N__35142),
            .I(N__35081));
    LocalMux I__8838 (
            .O(N__35139),
            .I(N__35071));
    LocalMux I__8837 (
            .O(N__35136),
            .I(N__35071));
    LocalMux I__8836 (
            .O(N__35129),
            .I(N__35071));
    LocalMux I__8835 (
            .O(N__35126),
            .I(N__35071));
    InMux I__8834 (
            .O(N__35123),
            .I(N__35064));
    InMux I__8833 (
            .O(N__35122),
            .I(N__35064));
    InMux I__8832 (
            .O(N__35121),
            .I(N__35064));
    InMux I__8831 (
            .O(N__35120),
            .I(N__35061));
    InMux I__8830 (
            .O(N__35119),
            .I(N__35058));
    Span4Mux_v I__8829 (
            .O(N__35116),
            .I(N__35049));
    LocalMux I__8828 (
            .O(N__35111),
            .I(N__35049));
    LocalMux I__8827 (
            .O(N__35106),
            .I(N__35049));
    LocalMux I__8826 (
            .O(N__35099),
            .I(N__35049));
    InMux I__8825 (
            .O(N__35098),
            .I(N__35046));
    Span4Mux_h I__8824 (
            .O(N__35095),
            .I(N__35043));
    LocalMux I__8823 (
            .O(N__35090),
            .I(N__35038));
    Span4Mux_h I__8822 (
            .O(N__35081),
            .I(N__35038));
    InMux I__8821 (
            .O(N__35080),
            .I(N__35035));
    Span12Mux_h I__8820 (
            .O(N__35071),
            .I(N__35032));
    LocalMux I__8819 (
            .O(N__35064),
            .I(N__35027));
    LocalMux I__8818 (
            .O(N__35061),
            .I(N__35027));
    LocalMux I__8817 (
            .O(N__35058),
            .I(N__35020));
    Span4Mux_v I__8816 (
            .O(N__35049),
            .I(N__35020));
    LocalMux I__8815 (
            .O(N__35046),
            .I(N__35020));
    Span4Mux_h I__8814 (
            .O(N__35043),
            .I(N__35015));
    Span4Mux_h I__8813 (
            .O(N__35038),
            .I(N__35015));
    LocalMux I__8812 (
            .O(N__35035),
            .I(N_156_0));
    Odrv12 I__8811 (
            .O(N__35032),
            .I(N_156_0));
    Odrv12 I__8810 (
            .O(N__35027),
            .I(N_156_0));
    Odrv4 I__8809 (
            .O(N__35020),
            .I(N_156_0));
    Odrv4 I__8808 (
            .O(N__35015),
            .I(N_156_0));
    CascadeMux I__8807 (
            .O(N__35004),
            .I(N__34991));
    CascadeMux I__8806 (
            .O(N__35003),
            .I(N__34983));
    InMux I__8805 (
            .O(N__35002),
            .I(N__34975));
    InMux I__8804 (
            .O(N__35001),
            .I(N__34966));
    InMux I__8803 (
            .O(N__35000),
            .I(N__34966));
    InMux I__8802 (
            .O(N__34999),
            .I(N__34966));
    InMux I__8801 (
            .O(N__34998),
            .I(N__34966));
    InMux I__8800 (
            .O(N__34997),
            .I(N__34963));
    CascadeMux I__8799 (
            .O(N__34996),
            .I(N__34959));
    InMux I__8798 (
            .O(N__34995),
            .I(N__34954));
    InMux I__8797 (
            .O(N__34994),
            .I(N__34954));
    InMux I__8796 (
            .O(N__34991),
            .I(N__34947));
    InMux I__8795 (
            .O(N__34990),
            .I(N__34940));
    InMux I__8794 (
            .O(N__34989),
            .I(N__34940));
    InMux I__8793 (
            .O(N__34988),
            .I(N__34940));
    InMux I__8792 (
            .O(N__34987),
            .I(N__34930));
    InMux I__8791 (
            .O(N__34986),
            .I(N__34930));
    InMux I__8790 (
            .O(N__34983),
            .I(N__34927));
    InMux I__8789 (
            .O(N__34982),
            .I(N__34924));
    InMux I__8788 (
            .O(N__34981),
            .I(N__34911));
    InMux I__8787 (
            .O(N__34980),
            .I(N__34911));
    InMux I__8786 (
            .O(N__34979),
            .I(N__34911));
    InMux I__8785 (
            .O(N__34978),
            .I(N__34911));
    LocalMux I__8784 (
            .O(N__34975),
            .I(N__34908));
    LocalMux I__8783 (
            .O(N__34966),
            .I(N__34903));
    LocalMux I__8782 (
            .O(N__34963),
            .I(N__34903));
    InMux I__8781 (
            .O(N__34962),
            .I(N__34900));
    InMux I__8780 (
            .O(N__34959),
            .I(N__34897));
    LocalMux I__8779 (
            .O(N__34954),
            .I(N__34894));
    InMux I__8778 (
            .O(N__34953),
            .I(N__34882));
    InMux I__8777 (
            .O(N__34952),
            .I(N__34882));
    InMux I__8776 (
            .O(N__34951),
            .I(N__34882));
    InMux I__8775 (
            .O(N__34950),
            .I(N__34879));
    LocalMux I__8774 (
            .O(N__34947),
            .I(N__34874));
    LocalMux I__8773 (
            .O(N__34940),
            .I(N__34874));
    InMux I__8772 (
            .O(N__34939),
            .I(N__34867));
    InMux I__8771 (
            .O(N__34938),
            .I(N__34867));
    InMux I__8770 (
            .O(N__34937),
            .I(N__34867));
    InMux I__8769 (
            .O(N__34936),
            .I(N__34862));
    InMux I__8768 (
            .O(N__34935),
            .I(N__34862));
    LocalMux I__8767 (
            .O(N__34930),
            .I(N__34857));
    LocalMux I__8766 (
            .O(N__34927),
            .I(N__34857));
    LocalMux I__8765 (
            .O(N__34924),
            .I(N__34854));
    InMux I__8764 (
            .O(N__34923),
            .I(N__34851));
    InMux I__8763 (
            .O(N__34922),
            .I(N__34848));
    InMux I__8762 (
            .O(N__34921),
            .I(N__34843));
    InMux I__8761 (
            .O(N__34920),
            .I(N__34843));
    LocalMux I__8760 (
            .O(N__34911),
            .I(N__34836));
    Span4Mux_v I__8759 (
            .O(N__34908),
            .I(N__34836));
    Span4Mux_v I__8758 (
            .O(N__34903),
            .I(N__34836));
    LocalMux I__8757 (
            .O(N__34900),
            .I(N__34833));
    LocalMux I__8756 (
            .O(N__34897),
            .I(N__34828));
    Span4Mux_v I__8755 (
            .O(N__34894),
            .I(N__34828));
    InMux I__8754 (
            .O(N__34893),
            .I(N__34817));
    InMux I__8753 (
            .O(N__34892),
            .I(N__34817));
    InMux I__8752 (
            .O(N__34891),
            .I(N__34817));
    InMux I__8751 (
            .O(N__34890),
            .I(N__34817));
    InMux I__8750 (
            .O(N__34889),
            .I(N__34817));
    LocalMux I__8749 (
            .O(N__34882),
            .I(N__34814));
    LocalMux I__8748 (
            .O(N__34879),
            .I(N__34803));
    Span4Mux_h I__8747 (
            .O(N__34874),
            .I(N__34803));
    LocalMux I__8746 (
            .O(N__34867),
            .I(N__34803));
    LocalMux I__8745 (
            .O(N__34862),
            .I(N__34803));
    Span4Mux_h I__8744 (
            .O(N__34857),
            .I(N__34803));
    Odrv12 I__8743 (
            .O(N__34854),
            .I(M_this_oam_address_qZ0Z_0));
    LocalMux I__8742 (
            .O(N__34851),
            .I(M_this_oam_address_qZ0Z_0));
    LocalMux I__8741 (
            .O(N__34848),
            .I(M_this_oam_address_qZ0Z_0));
    LocalMux I__8740 (
            .O(N__34843),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__8739 (
            .O(N__34836),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__8738 (
            .O(N__34833),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__8737 (
            .O(N__34828),
            .I(M_this_oam_address_qZ0Z_0));
    LocalMux I__8736 (
            .O(N__34817),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__8735 (
            .O(N__34814),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__8734 (
            .O(N__34803),
            .I(M_this_oam_address_qZ0Z_0));
    InMux I__8733 (
            .O(N__34782),
            .I(N__34779));
    LocalMux I__8732 (
            .O(N__34779),
            .I(N__34776));
    Span4Mux_v I__8731 (
            .O(N__34776),
            .I(N__34773));
    Odrv4 I__8730 (
            .O(N__34773),
            .I(N_69_0));
    CascadeMux I__8729 (
            .O(N__34770),
            .I(N__34767));
    InMux I__8728 (
            .O(N__34767),
            .I(N__34763));
    InMux I__8727 (
            .O(N__34766),
            .I(N__34758));
    LocalMux I__8726 (
            .O(N__34763),
            .I(N__34754));
    CascadeMux I__8725 (
            .O(N__34762),
            .I(N__34751));
    CascadeMux I__8724 (
            .O(N__34761),
            .I(N__34747));
    LocalMux I__8723 (
            .O(N__34758),
            .I(N__34744));
    InMux I__8722 (
            .O(N__34757),
            .I(N__34741));
    Span4Mux_v I__8721 (
            .O(N__34754),
            .I(N__34736));
    InMux I__8720 (
            .O(N__34751),
            .I(N__34733));
    InMux I__8719 (
            .O(N__34750),
            .I(N__34730));
    InMux I__8718 (
            .O(N__34747),
            .I(N__34727));
    Span4Mux_h I__8717 (
            .O(N__34744),
            .I(N__34722));
    LocalMux I__8716 (
            .O(N__34741),
            .I(N__34722));
    InMux I__8715 (
            .O(N__34740),
            .I(N__34719));
    CascadeMux I__8714 (
            .O(N__34739),
            .I(N__34716));
    Span4Mux_h I__8713 (
            .O(N__34736),
            .I(N__34707));
    LocalMux I__8712 (
            .O(N__34733),
            .I(N__34707));
    LocalMux I__8711 (
            .O(N__34730),
            .I(N__34707));
    LocalMux I__8710 (
            .O(N__34727),
            .I(N__34707));
    Span4Mux_v I__8709 (
            .O(N__34722),
            .I(N__34702));
    LocalMux I__8708 (
            .O(N__34719),
            .I(N__34699));
    InMux I__8707 (
            .O(N__34716),
            .I(N__34696));
    Span4Mux_v I__8706 (
            .O(N__34707),
            .I(N__34691));
    InMux I__8705 (
            .O(N__34706),
            .I(N__34688));
    CascadeMux I__8704 (
            .O(N__34705),
            .I(N__34685));
    Span4Mux_h I__8703 (
            .O(N__34702),
            .I(N__34679));
    Span4Mux_v I__8702 (
            .O(N__34699),
            .I(N__34679));
    LocalMux I__8701 (
            .O(N__34696),
            .I(N__34676));
    InMux I__8700 (
            .O(N__34695),
            .I(N__34673));
    CascadeMux I__8699 (
            .O(N__34694),
            .I(N__34670));
    Span4Mux_h I__8698 (
            .O(N__34691),
            .I(N__34665));
    LocalMux I__8697 (
            .O(N__34688),
            .I(N__34665));
    InMux I__8696 (
            .O(N__34685),
            .I(N__34659));
    InMux I__8695 (
            .O(N__34684),
            .I(N__34659));
    Span4Mux_h I__8694 (
            .O(N__34679),
            .I(N__34652));
    Span4Mux_v I__8693 (
            .O(N__34676),
            .I(N__34652));
    LocalMux I__8692 (
            .O(N__34673),
            .I(N__34652));
    InMux I__8691 (
            .O(N__34670),
            .I(N__34649));
    Span4Mux_v I__8690 (
            .O(N__34665),
            .I(N__34646));
    InMux I__8689 (
            .O(N__34664),
            .I(N__34643));
    LocalMux I__8688 (
            .O(N__34659),
            .I(N__34640));
    Span4Mux_h I__8687 (
            .O(N__34652),
            .I(N__34635));
    LocalMux I__8686 (
            .O(N__34649),
            .I(N__34635));
    Span4Mux_h I__8685 (
            .O(N__34646),
            .I(N__34630));
    LocalMux I__8684 (
            .O(N__34643),
            .I(N__34630));
    Span12Mux_v I__8683 (
            .O(N__34640),
            .I(N__34627));
    Span4Mux_h I__8682 (
            .O(N__34635),
            .I(N__34624));
    Span4Mux_v I__8681 (
            .O(N__34630),
            .I(N__34621));
    Span12Mux_h I__8680 (
            .O(N__34627),
            .I(N__34618));
    IoSpan4Mux I__8679 (
            .O(N__34624),
            .I(N__34615));
    Span4Mux_h I__8678 (
            .O(N__34621),
            .I(N__34612));
    Odrv12 I__8677 (
            .O(N__34618),
            .I(port_data_c_5));
    Odrv4 I__8676 (
            .O(N__34615),
            .I(port_data_c_5));
    Odrv4 I__8675 (
            .O(N__34612),
            .I(port_data_c_5));
    CascadeMux I__8674 (
            .O(N__34605),
            .I(N__34602));
    InMux I__8673 (
            .O(N__34602),
            .I(N__34599));
    LocalMux I__8672 (
            .O(N__34599),
            .I(M_this_data_tmp_qZ0Z_5));
    ClkMux I__8671 (
            .O(N__34596),
            .I(N__34206));
    ClkMux I__8670 (
            .O(N__34595),
            .I(N__34206));
    ClkMux I__8669 (
            .O(N__34594),
            .I(N__34206));
    ClkMux I__8668 (
            .O(N__34593),
            .I(N__34206));
    ClkMux I__8667 (
            .O(N__34592),
            .I(N__34206));
    ClkMux I__8666 (
            .O(N__34591),
            .I(N__34206));
    ClkMux I__8665 (
            .O(N__34590),
            .I(N__34206));
    ClkMux I__8664 (
            .O(N__34589),
            .I(N__34206));
    ClkMux I__8663 (
            .O(N__34588),
            .I(N__34206));
    ClkMux I__8662 (
            .O(N__34587),
            .I(N__34206));
    ClkMux I__8661 (
            .O(N__34586),
            .I(N__34206));
    ClkMux I__8660 (
            .O(N__34585),
            .I(N__34206));
    ClkMux I__8659 (
            .O(N__34584),
            .I(N__34206));
    ClkMux I__8658 (
            .O(N__34583),
            .I(N__34206));
    ClkMux I__8657 (
            .O(N__34582),
            .I(N__34206));
    ClkMux I__8656 (
            .O(N__34581),
            .I(N__34206));
    ClkMux I__8655 (
            .O(N__34580),
            .I(N__34206));
    ClkMux I__8654 (
            .O(N__34579),
            .I(N__34206));
    ClkMux I__8653 (
            .O(N__34578),
            .I(N__34206));
    ClkMux I__8652 (
            .O(N__34577),
            .I(N__34206));
    ClkMux I__8651 (
            .O(N__34576),
            .I(N__34206));
    ClkMux I__8650 (
            .O(N__34575),
            .I(N__34206));
    ClkMux I__8649 (
            .O(N__34574),
            .I(N__34206));
    ClkMux I__8648 (
            .O(N__34573),
            .I(N__34206));
    ClkMux I__8647 (
            .O(N__34572),
            .I(N__34206));
    ClkMux I__8646 (
            .O(N__34571),
            .I(N__34206));
    ClkMux I__8645 (
            .O(N__34570),
            .I(N__34206));
    ClkMux I__8644 (
            .O(N__34569),
            .I(N__34206));
    ClkMux I__8643 (
            .O(N__34568),
            .I(N__34206));
    ClkMux I__8642 (
            .O(N__34567),
            .I(N__34206));
    ClkMux I__8641 (
            .O(N__34566),
            .I(N__34206));
    ClkMux I__8640 (
            .O(N__34565),
            .I(N__34206));
    ClkMux I__8639 (
            .O(N__34564),
            .I(N__34206));
    ClkMux I__8638 (
            .O(N__34563),
            .I(N__34206));
    ClkMux I__8637 (
            .O(N__34562),
            .I(N__34206));
    ClkMux I__8636 (
            .O(N__34561),
            .I(N__34206));
    ClkMux I__8635 (
            .O(N__34560),
            .I(N__34206));
    ClkMux I__8634 (
            .O(N__34559),
            .I(N__34206));
    ClkMux I__8633 (
            .O(N__34558),
            .I(N__34206));
    ClkMux I__8632 (
            .O(N__34557),
            .I(N__34206));
    ClkMux I__8631 (
            .O(N__34556),
            .I(N__34206));
    ClkMux I__8630 (
            .O(N__34555),
            .I(N__34206));
    ClkMux I__8629 (
            .O(N__34554),
            .I(N__34206));
    ClkMux I__8628 (
            .O(N__34553),
            .I(N__34206));
    ClkMux I__8627 (
            .O(N__34552),
            .I(N__34206));
    ClkMux I__8626 (
            .O(N__34551),
            .I(N__34206));
    ClkMux I__8625 (
            .O(N__34550),
            .I(N__34206));
    ClkMux I__8624 (
            .O(N__34549),
            .I(N__34206));
    ClkMux I__8623 (
            .O(N__34548),
            .I(N__34206));
    ClkMux I__8622 (
            .O(N__34547),
            .I(N__34206));
    ClkMux I__8621 (
            .O(N__34546),
            .I(N__34206));
    ClkMux I__8620 (
            .O(N__34545),
            .I(N__34206));
    ClkMux I__8619 (
            .O(N__34544),
            .I(N__34206));
    ClkMux I__8618 (
            .O(N__34543),
            .I(N__34206));
    ClkMux I__8617 (
            .O(N__34542),
            .I(N__34206));
    ClkMux I__8616 (
            .O(N__34541),
            .I(N__34206));
    ClkMux I__8615 (
            .O(N__34540),
            .I(N__34206));
    ClkMux I__8614 (
            .O(N__34539),
            .I(N__34206));
    ClkMux I__8613 (
            .O(N__34538),
            .I(N__34206));
    ClkMux I__8612 (
            .O(N__34537),
            .I(N__34206));
    ClkMux I__8611 (
            .O(N__34536),
            .I(N__34206));
    ClkMux I__8610 (
            .O(N__34535),
            .I(N__34206));
    ClkMux I__8609 (
            .O(N__34534),
            .I(N__34206));
    ClkMux I__8608 (
            .O(N__34533),
            .I(N__34206));
    ClkMux I__8607 (
            .O(N__34532),
            .I(N__34206));
    ClkMux I__8606 (
            .O(N__34531),
            .I(N__34206));
    ClkMux I__8605 (
            .O(N__34530),
            .I(N__34206));
    ClkMux I__8604 (
            .O(N__34529),
            .I(N__34206));
    ClkMux I__8603 (
            .O(N__34528),
            .I(N__34206));
    ClkMux I__8602 (
            .O(N__34527),
            .I(N__34206));
    ClkMux I__8601 (
            .O(N__34526),
            .I(N__34206));
    ClkMux I__8600 (
            .O(N__34525),
            .I(N__34206));
    ClkMux I__8599 (
            .O(N__34524),
            .I(N__34206));
    ClkMux I__8598 (
            .O(N__34523),
            .I(N__34206));
    ClkMux I__8597 (
            .O(N__34522),
            .I(N__34206));
    ClkMux I__8596 (
            .O(N__34521),
            .I(N__34206));
    ClkMux I__8595 (
            .O(N__34520),
            .I(N__34206));
    ClkMux I__8594 (
            .O(N__34519),
            .I(N__34206));
    ClkMux I__8593 (
            .O(N__34518),
            .I(N__34206));
    ClkMux I__8592 (
            .O(N__34517),
            .I(N__34206));
    ClkMux I__8591 (
            .O(N__34516),
            .I(N__34206));
    ClkMux I__8590 (
            .O(N__34515),
            .I(N__34206));
    ClkMux I__8589 (
            .O(N__34514),
            .I(N__34206));
    ClkMux I__8588 (
            .O(N__34513),
            .I(N__34206));
    ClkMux I__8587 (
            .O(N__34512),
            .I(N__34206));
    ClkMux I__8586 (
            .O(N__34511),
            .I(N__34206));
    ClkMux I__8585 (
            .O(N__34510),
            .I(N__34206));
    ClkMux I__8584 (
            .O(N__34509),
            .I(N__34206));
    ClkMux I__8583 (
            .O(N__34508),
            .I(N__34206));
    ClkMux I__8582 (
            .O(N__34507),
            .I(N__34206));
    ClkMux I__8581 (
            .O(N__34506),
            .I(N__34206));
    ClkMux I__8580 (
            .O(N__34505),
            .I(N__34206));
    ClkMux I__8579 (
            .O(N__34504),
            .I(N__34206));
    ClkMux I__8578 (
            .O(N__34503),
            .I(N__34206));
    ClkMux I__8577 (
            .O(N__34502),
            .I(N__34206));
    ClkMux I__8576 (
            .O(N__34501),
            .I(N__34206));
    ClkMux I__8575 (
            .O(N__34500),
            .I(N__34206));
    ClkMux I__8574 (
            .O(N__34499),
            .I(N__34206));
    ClkMux I__8573 (
            .O(N__34498),
            .I(N__34206));
    ClkMux I__8572 (
            .O(N__34497),
            .I(N__34206));
    ClkMux I__8571 (
            .O(N__34496),
            .I(N__34206));
    ClkMux I__8570 (
            .O(N__34495),
            .I(N__34206));
    ClkMux I__8569 (
            .O(N__34494),
            .I(N__34206));
    ClkMux I__8568 (
            .O(N__34493),
            .I(N__34206));
    ClkMux I__8567 (
            .O(N__34492),
            .I(N__34206));
    ClkMux I__8566 (
            .O(N__34491),
            .I(N__34206));
    ClkMux I__8565 (
            .O(N__34490),
            .I(N__34206));
    ClkMux I__8564 (
            .O(N__34489),
            .I(N__34206));
    ClkMux I__8563 (
            .O(N__34488),
            .I(N__34206));
    ClkMux I__8562 (
            .O(N__34487),
            .I(N__34206));
    ClkMux I__8561 (
            .O(N__34486),
            .I(N__34206));
    ClkMux I__8560 (
            .O(N__34485),
            .I(N__34206));
    ClkMux I__8559 (
            .O(N__34484),
            .I(N__34206));
    ClkMux I__8558 (
            .O(N__34483),
            .I(N__34206));
    ClkMux I__8557 (
            .O(N__34482),
            .I(N__34206));
    ClkMux I__8556 (
            .O(N__34481),
            .I(N__34206));
    ClkMux I__8555 (
            .O(N__34480),
            .I(N__34206));
    ClkMux I__8554 (
            .O(N__34479),
            .I(N__34206));
    ClkMux I__8553 (
            .O(N__34478),
            .I(N__34206));
    ClkMux I__8552 (
            .O(N__34477),
            .I(N__34206));
    ClkMux I__8551 (
            .O(N__34476),
            .I(N__34206));
    ClkMux I__8550 (
            .O(N__34475),
            .I(N__34206));
    ClkMux I__8549 (
            .O(N__34474),
            .I(N__34206));
    ClkMux I__8548 (
            .O(N__34473),
            .I(N__34206));
    ClkMux I__8547 (
            .O(N__34472),
            .I(N__34206));
    ClkMux I__8546 (
            .O(N__34471),
            .I(N__34206));
    ClkMux I__8545 (
            .O(N__34470),
            .I(N__34206));
    ClkMux I__8544 (
            .O(N__34469),
            .I(N__34206));
    ClkMux I__8543 (
            .O(N__34468),
            .I(N__34206));
    ClkMux I__8542 (
            .O(N__34467),
            .I(N__34206));
    GlobalMux I__8541 (
            .O(N__34206),
            .I(N__34203));
    gio2CtrlBuf I__8540 (
            .O(N__34203),
            .I(clk_0_c_g));
    CEMux I__8539 (
            .O(N__34200),
            .I(N__34195));
    CEMux I__8538 (
            .O(N__34199),
            .I(N__34192));
    CEMux I__8537 (
            .O(N__34198),
            .I(N__34189));
    LocalMux I__8536 (
            .O(N__34195),
            .I(N__34184));
    LocalMux I__8535 (
            .O(N__34192),
            .I(N__34179));
    LocalMux I__8534 (
            .O(N__34189),
            .I(N__34179));
    CEMux I__8533 (
            .O(N__34188),
            .I(N__34176));
    CEMux I__8532 (
            .O(N__34187),
            .I(N__34173));
    Span4Mux_v I__8531 (
            .O(N__34184),
            .I(N__34170));
    Span4Mux_v I__8530 (
            .O(N__34179),
            .I(N__34167));
    LocalMux I__8529 (
            .O(N__34176),
            .I(N__34164));
    LocalMux I__8528 (
            .O(N__34173),
            .I(N__34159));
    Span4Mux_h I__8527 (
            .O(N__34170),
            .I(N__34152));
    Span4Mux_v I__8526 (
            .O(N__34167),
            .I(N__34152));
    Span4Mux_h I__8525 (
            .O(N__34164),
            .I(N__34152));
    CEMux I__8524 (
            .O(N__34163),
            .I(N__34149));
    CEMux I__8523 (
            .O(N__34162),
            .I(N__34146));
    Span4Mux_v I__8522 (
            .O(N__34159),
            .I(N__34143));
    Span4Mux_h I__8521 (
            .O(N__34152),
            .I(N__34138));
    LocalMux I__8520 (
            .O(N__34149),
            .I(N__34138));
    LocalMux I__8519 (
            .O(N__34146),
            .I(N__34135));
    Span4Mux_h I__8518 (
            .O(N__34143),
            .I(N__34130));
    Span4Mux_h I__8517 (
            .O(N__34138),
            .I(N__34130));
    Odrv12 I__8516 (
            .O(N__34135),
            .I(N_1142_0));
    Odrv4 I__8515 (
            .O(N__34130),
            .I(N_1142_0));
    InMux I__8514 (
            .O(N__34125),
            .I(N__34101));
    InMux I__8513 (
            .O(N__34124),
            .I(N__34098));
    InMux I__8512 (
            .O(N__34123),
            .I(N__34095));
    InMux I__8511 (
            .O(N__34122),
            .I(N__34092));
    InMux I__8510 (
            .O(N__34121),
            .I(N__34085));
    InMux I__8509 (
            .O(N__34120),
            .I(N__34085));
    InMux I__8508 (
            .O(N__34119),
            .I(N__34085));
    InMux I__8507 (
            .O(N__34118),
            .I(N__34082));
    InMux I__8506 (
            .O(N__34117),
            .I(N__34079));
    InMux I__8505 (
            .O(N__34116),
            .I(N__34076));
    InMux I__8504 (
            .O(N__34115),
            .I(N__34073));
    InMux I__8503 (
            .O(N__34114),
            .I(N__34070));
    InMux I__8502 (
            .O(N__34113),
            .I(N__34067));
    InMux I__8501 (
            .O(N__34112),
            .I(N__34064));
    InMux I__8500 (
            .O(N__34111),
            .I(N__34061));
    InMux I__8499 (
            .O(N__34110),
            .I(N__34058));
    InMux I__8498 (
            .O(N__34109),
            .I(N__34055));
    InMux I__8497 (
            .O(N__34108),
            .I(N__34052));
    InMux I__8496 (
            .O(N__34107),
            .I(N__34049));
    InMux I__8495 (
            .O(N__34106),
            .I(N__34046));
    InMux I__8494 (
            .O(N__34105),
            .I(N__34041));
    InMux I__8493 (
            .O(N__34104),
            .I(N__34041));
    LocalMux I__8492 (
            .O(N__34101),
            .I(N__34007));
    LocalMux I__8491 (
            .O(N__34098),
            .I(N__34004));
    LocalMux I__8490 (
            .O(N__34095),
            .I(N__34001));
    LocalMux I__8489 (
            .O(N__34092),
            .I(N__33998));
    LocalMux I__8488 (
            .O(N__34085),
            .I(N__33995));
    LocalMux I__8487 (
            .O(N__34082),
            .I(N__33992));
    LocalMux I__8486 (
            .O(N__34079),
            .I(N__33989));
    LocalMux I__8485 (
            .O(N__34076),
            .I(N__33986));
    LocalMux I__8484 (
            .O(N__34073),
            .I(N__33983));
    LocalMux I__8483 (
            .O(N__34070),
            .I(N__33980));
    LocalMux I__8482 (
            .O(N__34067),
            .I(N__33977));
    LocalMux I__8481 (
            .O(N__34064),
            .I(N__33974));
    LocalMux I__8480 (
            .O(N__34061),
            .I(N__33971));
    LocalMux I__8479 (
            .O(N__34058),
            .I(N__33968));
    LocalMux I__8478 (
            .O(N__34055),
            .I(N__33965));
    LocalMux I__8477 (
            .O(N__34052),
            .I(N__33962));
    LocalMux I__8476 (
            .O(N__34049),
            .I(N__33959));
    LocalMux I__8475 (
            .O(N__34046),
            .I(N__33956));
    LocalMux I__8474 (
            .O(N__34041),
            .I(N__33953));
    SRMux I__8473 (
            .O(N__34040),
            .I(N__33852));
    SRMux I__8472 (
            .O(N__34039),
            .I(N__33852));
    SRMux I__8471 (
            .O(N__34038),
            .I(N__33852));
    SRMux I__8470 (
            .O(N__34037),
            .I(N__33852));
    SRMux I__8469 (
            .O(N__34036),
            .I(N__33852));
    SRMux I__8468 (
            .O(N__34035),
            .I(N__33852));
    SRMux I__8467 (
            .O(N__34034),
            .I(N__33852));
    SRMux I__8466 (
            .O(N__34033),
            .I(N__33852));
    SRMux I__8465 (
            .O(N__34032),
            .I(N__33852));
    SRMux I__8464 (
            .O(N__34031),
            .I(N__33852));
    SRMux I__8463 (
            .O(N__34030),
            .I(N__33852));
    SRMux I__8462 (
            .O(N__34029),
            .I(N__33852));
    SRMux I__8461 (
            .O(N__34028),
            .I(N__33852));
    SRMux I__8460 (
            .O(N__34027),
            .I(N__33852));
    SRMux I__8459 (
            .O(N__34026),
            .I(N__33852));
    SRMux I__8458 (
            .O(N__34025),
            .I(N__33852));
    SRMux I__8457 (
            .O(N__34024),
            .I(N__33852));
    SRMux I__8456 (
            .O(N__34023),
            .I(N__33852));
    SRMux I__8455 (
            .O(N__34022),
            .I(N__33852));
    SRMux I__8454 (
            .O(N__34021),
            .I(N__33852));
    SRMux I__8453 (
            .O(N__34020),
            .I(N__33852));
    SRMux I__8452 (
            .O(N__34019),
            .I(N__33852));
    SRMux I__8451 (
            .O(N__34018),
            .I(N__33852));
    SRMux I__8450 (
            .O(N__34017),
            .I(N__33852));
    SRMux I__8449 (
            .O(N__34016),
            .I(N__33852));
    SRMux I__8448 (
            .O(N__34015),
            .I(N__33852));
    SRMux I__8447 (
            .O(N__34014),
            .I(N__33852));
    SRMux I__8446 (
            .O(N__34013),
            .I(N__33852));
    SRMux I__8445 (
            .O(N__34012),
            .I(N__33852));
    SRMux I__8444 (
            .O(N__34011),
            .I(N__33852));
    SRMux I__8443 (
            .O(N__34010),
            .I(N__33852));
    Glb2LocalMux I__8442 (
            .O(N__34007),
            .I(N__33852));
    Glb2LocalMux I__8441 (
            .O(N__34004),
            .I(N__33852));
    Glb2LocalMux I__8440 (
            .O(N__34001),
            .I(N__33852));
    Glb2LocalMux I__8439 (
            .O(N__33998),
            .I(N__33852));
    Glb2LocalMux I__8438 (
            .O(N__33995),
            .I(N__33852));
    Glb2LocalMux I__8437 (
            .O(N__33992),
            .I(N__33852));
    Glb2LocalMux I__8436 (
            .O(N__33989),
            .I(N__33852));
    Glb2LocalMux I__8435 (
            .O(N__33986),
            .I(N__33852));
    Glb2LocalMux I__8434 (
            .O(N__33983),
            .I(N__33852));
    Glb2LocalMux I__8433 (
            .O(N__33980),
            .I(N__33852));
    Glb2LocalMux I__8432 (
            .O(N__33977),
            .I(N__33852));
    Glb2LocalMux I__8431 (
            .O(N__33974),
            .I(N__33852));
    Glb2LocalMux I__8430 (
            .O(N__33971),
            .I(N__33852));
    Glb2LocalMux I__8429 (
            .O(N__33968),
            .I(N__33852));
    Glb2LocalMux I__8428 (
            .O(N__33965),
            .I(N__33852));
    Glb2LocalMux I__8427 (
            .O(N__33962),
            .I(N__33852));
    Glb2LocalMux I__8426 (
            .O(N__33959),
            .I(N__33852));
    Glb2LocalMux I__8425 (
            .O(N__33956),
            .I(N__33852));
    Glb2LocalMux I__8424 (
            .O(N__33953),
            .I(N__33852));
    GlobalMux I__8423 (
            .O(N__33852),
            .I(N__33849));
    gio2CtrlBuf I__8422 (
            .O(N__33849),
            .I(M_this_reset_cond_out_g_0));
    InMux I__8421 (
            .O(N__33846),
            .I(N__33843));
    LocalMux I__8420 (
            .O(N__33843),
            .I(N__33840));
    Span4Mux_v I__8419 (
            .O(N__33840),
            .I(N__33837));
    Odrv4 I__8418 (
            .O(N__33837),
            .I(un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0));
    CascadeMux I__8417 (
            .O(N__33834),
            .I(N__33830));
    CascadeMux I__8416 (
            .O(N__33833),
            .I(N__33827));
    InMux I__8415 (
            .O(N__33830),
            .I(N__33822));
    InMux I__8414 (
            .O(N__33827),
            .I(N__33819));
    InMux I__8413 (
            .O(N__33826),
            .I(N__33815));
    InMux I__8412 (
            .O(N__33825),
            .I(N__33810));
    LocalMux I__8411 (
            .O(N__33822),
            .I(N__33807));
    LocalMux I__8410 (
            .O(N__33819),
            .I(N__33804));
    CascadeMux I__8409 (
            .O(N__33818),
            .I(N__33801));
    LocalMux I__8408 (
            .O(N__33815),
            .I(N__33796));
    InMux I__8407 (
            .O(N__33814),
            .I(N__33791));
    InMux I__8406 (
            .O(N__33813),
            .I(N__33791));
    LocalMux I__8405 (
            .O(N__33810),
            .I(N__33788));
    Span4Mux_v I__8404 (
            .O(N__33807),
            .I(N__33785));
    Span4Mux_h I__8403 (
            .O(N__33804),
            .I(N__33782));
    InMux I__8402 (
            .O(N__33801),
            .I(N__33779));
    InMux I__8401 (
            .O(N__33800),
            .I(N__33776));
    InMux I__8400 (
            .O(N__33799),
            .I(N__33773));
    Span4Mux_v I__8399 (
            .O(N__33796),
            .I(N__33770));
    LocalMux I__8398 (
            .O(N__33791),
            .I(N__33767));
    Span4Mux_v I__8397 (
            .O(N__33788),
            .I(N__33764));
    Span4Mux_h I__8396 (
            .O(N__33785),
            .I(N__33757));
    Span4Mux_v I__8395 (
            .O(N__33782),
            .I(N__33757));
    LocalMux I__8394 (
            .O(N__33779),
            .I(N__33757));
    LocalMux I__8393 (
            .O(N__33776),
            .I(N__33754));
    LocalMux I__8392 (
            .O(N__33773),
            .I(N__33751));
    Sp12to4 I__8391 (
            .O(N__33770),
            .I(N__33745));
    Span12Mux_v I__8390 (
            .O(N__33767),
            .I(N__33745));
    Span4Mux_v I__8389 (
            .O(N__33764),
            .I(N__33742));
    Span4Mux_h I__8388 (
            .O(N__33757),
            .I(N__33739));
    Span4Mux_v I__8387 (
            .O(N__33754),
            .I(N__33734));
    Span4Mux_v I__8386 (
            .O(N__33751),
            .I(N__33734));
    InMux I__8385 (
            .O(N__33750),
            .I(N__33731));
    Span12Mux_h I__8384 (
            .O(N__33745),
            .I(N__33728));
    Sp12to4 I__8383 (
            .O(N__33742),
            .I(N__33725));
    Span4Mux_v I__8382 (
            .O(N__33739),
            .I(N__33722));
    Span4Mux_h I__8381 (
            .O(N__33734),
            .I(N__33717));
    LocalMux I__8380 (
            .O(N__33731),
            .I(N__33717));
    Span12Mux_v I__8379 (
            .O(N__33728),
            .I(N__33714));
    Span12Mux_h I__8378 (
            .O(N__33725),
            .I(N__33711));
    Span4Mux_h I__8377 (
            .O(N__33722),
            .I(N__33708));
    Sp12to4 I__8376 (
            .O(N__33717),
            .I(N__33705));
    Odrv12 I__8375 (
            .O(N__33714),
            .I(port_data_c_0));
    Odrv12 I__8374 (
            .O(N__33711),
            .I(port_data_c_0));
    Odrv4 I__8373 (
            .O(N__33708),
            .I(port_data_c_0));
    Odrv12 I__8372 (
            .O(N__33705),
            .I(port_data_c_0));
    IoInMux I__8371 (
            .O(N__33696),
            .I(N__33692));
    InMux I__8370 (
            .O(N__33695),
            .I(N__33689));
    LocalMux I__8369 (
            .O(N__33692),
            .I(N__33686));
    LocalMux I__8368 (
            .O(N__33689),
            .I(N__33683));
    Span12Mux_s10_v I__8367 (
            .O(N__33686),
            .I(N__33680));
    Span4Mux_h I__8366 (
            .O(N__33683),
            .I(N__33677));
    Odrv12 I__8365 (
            .O(N__33680),
            .I(M_this_external_address_qZ0Z_8));
    Odrv4 I__8364 (
            .O(N__33677),
            .I(M_this_external_address_qZ0Z_8));
    InMux I__8363 (
            .O(N__33672),
            .I(N__33665));
    InMux I__8362 (
            .O(N__33671),
            .I(N__33662));
    InMux I__8361 (
            .O(N__33670),
            .I(N__33659));
    InMux I__8360 (
            .O(N__33669),
            .I(N__33654));
    InMux I__8359 (
            .O(N__33668),
            .I(N__33651));
    LocalMux I__8358 (
            .O(N__33665),
            .I(N__33644));
    LocalMux I__8357 (
            .O(N__33662),
            .I(N__33644));
    LocalMux I__8356 (
            .O(N__33659),
            .I(N__33644));
    CascadeMux I__8355 (
            .O(N__33658),
            .I(N__33641));
    InMux I__8354 (
            .O(N__33657),
            .I(N__33638));
    LocalMux I__8353 (
            .O(N__33654),
            .I(N__33634));
    LocalMux I__8352 (
            .O(N__33651),
            .I(N__33631));
    Span4Mux_v I__8351 (
            .O(N__33644),
            .I(N__33626));
    InMux I__8350 (
            .O(N__33641),
            .I(N__33623));
    LocalMux I__8349 (
            .O(N__33638),
            .I(N__33620));
    CascadeMux I__8348 (
            .O(N__33637),
            .I(N__33617));
    Span4Mux_v I__8347 (
            .O(N__33634),
            .I(N__33614));
    Span4Mux_v I__8346 (
            .O(N__33631),
            .I(N__33611));
    InMux I__8345 (
            .O(N__33630),
            .I(N__33608));
    InMux I__8344 (
            .O(N__33629),
            .I(N__33605));
    Sp12to4 I__8343 (
            .O(N__33626),
            .I(N__33600));
    LocalMux I__8342 (
            .O(N__33623),
            .I(N__33600));
    Span12Mux_s10_v I__8341 (
            .O(N__33620),
            .I(N__33597));
    InMux I__8340 (
            .O(N__33617),
            .I(N__33594));
    Span4Mux_h I__8339 (
            .O(N__33614),
            .I(N__33589));
    Span4Mux_h I__8338 (
            .O(N__33611),
            .I(N__33589));
    LocalMux I__8337 (
            .O(N__33608),
            .I(N__33584));
    LocalMux I__8336 (
            .O(N__33605),
            .I(N__33584));
    Span12Mux_v I__8335 (
            .O(N__33600),
            .I(N__33581));
    Span12Mux_v I__8334 (
            .O(N__33597),
            .I(N__33578));
    LocalMux I__8333 (
            .O(N__33594),
            .I(N__33575));
    IoSpan4Mux I__8332 (
            .O(N__33589),
            .I(N__33572));
    Span4Mux_v I__8331 (
            .O(N__33584),
            .I(N__33569));
    Span12Mux_h I__8330 (
            .O(N__33581),
            .I(N__33566));
    Span12Mux_h I__8329 (
            .O(N__33578),
            .I(N__33561));
    Span12Mux_v I__8328 (
            .O(N__33575),
            .I(N__33561));
    IoSpan4Mux I__8327 (
            .O(N__33572),
            .I(N__33558));
    Sp12to4 I__8326 (
            .O(N__33569),
            .I(N__33555));
    Odrv12 I__8325 (
            .O(N__33566),
            .I(port_data_c_7));
    Odrv12 I__8324 (
            .O(N__33561),
            .I(port_data_c_7));
    Odrv4 I__8323 (
            .O(N__33558),
            .I(port_data_c_7));
    Odrv12 I__8322 (
            .O(N__33555),
            .I(port_data_c_7));
    InMux I__8321 (
            .O(N__33546),
            .I(N__33543));
    LocalMux I__8320 (
            .O(N__33543),
            .I(N__33540));
    Span4Mux_h I__8319 (
            .O(N__33540),
            .I(N__33537));
    Odrv4 I__8318 (
            .O(N__33537),
            .I(un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0));
    IoInMux I__8317 (
            .O(N__33534),
            .I(N__33531));
    LocalMux I__8316 (
            .O(N__33531),
            .I(N__33528));
    Span4Mux_s2_h I__8315 (
            .O(N__33528),
            .I(N__33525));
    Span4Mux_h I__8314 (
            .O(N__33525),
            .I(N__33521));
    InMux I__8313 (
            .O(N__33524),
            .I(N__33518));
    Sp12to4 I__8312 (
            .O(N__33521),
            .I(N__33515));
    LocalMux I__8311 (
            .O(N__33518),
            .I(N__33512));
    Span12Mux_v I__8310 (
            .O(N__33515),
            .I(N__33509));
    Span4Mux_h I__8309 (
            .O(N__33512),
            .I(N__33506));
    Odrv12 I__8308 (
            .O(N__33509),
            .I(M_this_external_address_qZ0Z_15));
    Odrv4 I__8307 (
            .O(N__33506),
            .I(M_this_external_address_qZ0Z_15));
    InMux I__8306 (
            .O(N__33501),
            .I(N__33498));
    LocalMux I__8305 (
            .O(N__33498),
            .I(N__33495));
    Odrv4 I__8304 (
            .O(N__33495),
            .I(un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0));
    InMux I__8303 (
            .O(N__33492),
            .I(N__33488));
    CascadeMux I__8302 (
            .O(N__33491),
            .I(N__33484));
    LocalMux I__8301 (
            .O(N__33488),
            .I(N__33479));
    InMux I__8300 (
            .O(N__33487),
            .I(N__33476));
    InMux I__8299 (
            .O(N__33484),
            .I(N__33473));
    CascadeMux I__8298 (
            .O(N__33483),
            .I(N__33468));
    CascadeMux I__8297 (
            .O(N__33482),
            .I(N__33465));
    Span4Mux_h I__8296 (
            .O(N__33479),
            .I(N__33458));
    LocalMux I__8295 (
            .O(N__33476),
            .I(N__33458));
    LocalMux I__8294 (
            .O(N__33473),
            .I(N__33458));
    InMux I__8293 (
            .O(N__33472),
            .I(N__33455));
    InMux I__8292 (
            .O(N__33471),
            .I(N__33451));
    InMux I__8291 (
            .O(N__33468),
            .I(N__33448));
    InMux I__8290 (
            .O(N__33465),
            .I(N__33445));
    Span4Mux_h I__8289 (
            .O(N__33458),
            .I(N__33440));
    LocalMux I__8288 (
            .O(N__33455),
            .I(N__33437));
    InMux I__8287 (
            .O(N__33454),
            .I(N__33434));
    LocalMux I__8286 (
            .O(N__33451),
            .I(N__33431));
    LocalMux I__8285 (
            .O(N__33448),
            .I(N__33428));
    LocalMux I__8284 (
            .O(N__33445),
            .I(N__33425));
    InMux I__8283 (
            .O(N__33444),
            .I(N__33422));
    InMux I__8282 (
            .O(N__33443),
            .I(N__33417));
    Span4Mux_h I__8281 (
            .O(N__33440),
            .I(N__33414));
    Span4Mux_h I__8280 (
            .O(N__33437),
            .I(N__33411));
    LocalMux I__8279 (
            .O(N__33434),
            .I(N__33408));
    Span4Mux_v I__8278 (
            .O(N__33431),
            .I(N__33401));
    Span4Mux_h I__8277 (
            .O(N__33428),
            .I(N__33401));
    Span4Mux_v I__8276 (
            .O(N__33425),
            .I(N__33401));
    LocalMux I__8275 (
            .O(N__33422),
            .I(N__33398));
    CascadeMux I__8274 (
            .O(N__33421),
            .I(N__33395));
    CascadeMux I__8273 (
            .O(N__33420),
            .I(N__33391));
    LocalMux I__8272 (
            .O(N__33417),
            .I(N__33388));
    Span4Mux_h I__8271 (
            .O(N__33414),
            .I(N__33383));
    Span4Mux_v I__8270 (
            .O(N__33411),
            .I(N__33383));
    Span4Mux_h I__8269 (
            .O(N__33408),
            .I(N__33380));
    Span4Mux_h I__8268 (
            .O(N__33401),
            .I(N__33375));
    Span4Mux_v I__8267 (
            .O(N__33398),
            .I(N__33375));
    InMux I__8266 (
            .O(N__33395),
            .I(N__33372));
    InMux I__8265 (
            .O(N__33394),
            .I(N__33369));
    InMux I__8264 (
            .O(N__33391),
            .I(N__33366));
    Span12Mux_h I__8263 (
            .O(N__33388),
            .I(N__33363));
    Span4Mux_v I__8262 (
            .O(N__33383),
            .I(N__33360));
    Span4Mux_h I__8261 (
            .O(N__33380),
            .I(N__33357));
    Span4Mux_h I__8260 (
            .O(N__33375),
            .I(N__33348));
    LocalMux I__8259 (
            .O(N__33372),
            .I(N__33348));
    LocalMux I__8258 (
            .O(N__33369),
            .I(N__33348));
    LocalMux I__8257 (
            .O(N__33366),
            .I(N__33348));
    Span12Mux_h I__8256 (
            .O(N__33363),
            .I(N__33345));
    Span4Mux_v I__8255 (
            .O(N__33360),
            .I(N__33342));
    Sp12to4 I__8254 (
            .O(N__33357),
            .I(N__33337));
    Sp12to4 I__8253 (
            .O(N__33348),
            .I(N__33337));
    Odrv12 I__8252 (
            .O(N__33345),
            .I(port_data_c_2));
    Odrv4 I__8251 (
            .O(N__33342),
            .I(port_data_c_2));
    Odrv12 I__8250 (
            .O(N__33337),
            .I(port_data_c_2));
    IoInMux I__8249 (
            .O(N__33330),
            .I(N__33327));
    LocalMux I__8248 (
            .O(N__33327),
            .I(N__33324));
    IoSpan4Mux I__8247 (
            .O(N__33324),
            .I(N__33321));
    Span4Mux_s1_v I__8246 (
            .O(N__33321),
            .I(N__33318));
    Span4Mux_v I__8245 (
            .O(N__33318),
            .I(N__33314));
    InMux I__8244 (
            .O(N__33317),
            .I(N__33311));
    Span4Mux_v I__8243 (
            .O(N__33314),
            .I(N__33306));
    LocalMux I__8242 (
            .O(N__33311),
            .I(N__33306));
    Odrv4 I__8241 (
            .O(N__33306),
            .I(M_this_external_address_qZ0Z_10));
    InMux I__8240 (
            .O(N__33303),
            .I(N__33300));
    LocalMux I__8239 (
            .O(N__33300),
            .I(N__33297));
    Span4Mux_v I__8238 (
            .O(N__33297),
            .I(N__33293));
    InMux I__8237 (
            .O(N__33296),
            .I(N__33290));
    Sp12to4 I__8236 (
            .O(N__33293),
            .I(N__33285));
    LocalMux I__8235 (
            .O(N__33290),
            .I(N__33285));
    Span12Mux_s11_h I__8234 (
            .O(N__33285),
            .I(N__33282));
    Odrv12 I__8233 (
            .O(N__33282),
            .I(un1_M_this_state_q_11_0_i));
    IoInMux I__8232 (
            .O(N__33279),
            .I(N__33276));
    LocalMux I__8231 (
            .O(N__33276),
            .I(N__33273));
    IoSpan4Mux I__8230 (
            .O(N__33273),
            .I(N__33269));
    CascadeMux I__8229 (
            .O(N__33272),
            .I(N__33266));
    IoSpan4Mux I__8228 (
            .O(N__33269),
            .I(N__33263));
    InMux I__8227 (
            .O(N__33266),
            .I(N__33259));
    IoSpan4Mux I__8226 (
            .O(N__33263),
            .I(N__33256));
    CascadeMux I__8225 (
            .O(N__33262),
            .I(N__33253));
    LocalMux I__8224 (
            .O(N__33259),
            .I(N__33250));
    Sp12to4 I__8223 (
            .O(N__33256),
            .I(N__33247));
    InMux I__8222 (
            .O(N__33253),
            .I(N__33244));
    Span4Mux_v I__8221 (
            .O(N__33250),
            .I(N__33241));
    Odrv12 I__8220 (
            .O(N__33247),
            .I(M_this_external_address_qZ0Z_0));
    LocalMux I__8219 (
            .O(N__33244),
            .I(M_this_external_address_qZ0Z_0));
    Odrv4 I__8218 (
            .O(N__33241),
            .I(M_this_external_address_qZ0Z_0));
    InMux I__8217 (
            .O(N__33234),
            .I(N__33231));
    LocalMux I__8216 (
            .O(N__33231),
            .I(N__33228));
    Span4Mux_h I__8215 (
            .O(N__33228),
            .I(N__33225));
    Odrv4 I__8214 (
            .O(N__33225),
            .I(un1_M_this_external_address_q_cry_0_THRU_CO));
    InMux I__8213 (
            .O(N__33222),
            .I(N__33217));
    IoInMux I__8212 (
            .O(N__33221),
            .I(N__33214));
    CascadeMux I__8211 (
            .O(N__33220),
            .I(N__33211));
    LocalMux I__8210 (
            .O(N__33217),
            .I(N__33208));
    LocalMux I__8209 (
            .O(N__33214),
            .I(N__33205));
    InMux I__8208 (
            .O(N__33211),
            .I(N__33202));
    Span4Mux_h I__8207 (
            .O(N__33208),
            .I(N__33199));
    Odrv12 I__8206 (
            .O(N__33205),
            .I(M_this_external_address_qZ0Z_1));
    LocalMux I__8205 (
            .O(N__33202),
            .I(M_this_external_address_qZ0Z_1));
    Odrv4 I__8204 (
            .O(N__33199),
            .I(M_this_external_address_qZ0Z_1));
    InMux I__8203 (
            .O(N__33192),
            .I(N__33189));
    LocalMux I__8202 (
            .O(N__33189),
            .I(N__33186));
    Span4Mux_h I__8201 (
            .O(N__33186),
            .I(N__33183));
    Odrv4 I__8200 (
            .O(N__33183),
            .I(un1_M_this_external_address_q_cry_1_THRU_CO));
    IoInMux I__8199 (
            .O(N__33180),
            .I(N__33177));
    LocalMux I__8198 (
            .O(N__33177),
            .I(N__33174));
    IoSpan4Mux I__8197 (
            .O(N__33174),
            .I(N__33169));
    InMux I__8196 (
            .O(N__33173),
            .I(N__33166));
    CascadeMux I__8195 (
            .O(N__33172),
            .I(N__33163));
    Span4Mux_s2_v I__8194 (
            .O(N__33169),
            .I(N__33160));
    LocalMux I__8193 (
            .O(N__33166),
            .I(N__33157));
    InMux I__8192 (
            .O(N__33163),
            .I(N__33154));
    Span4Mux_v I__8191 (
            .O(N__33160),
            .I(N__33149));
    Span4Mux_h I__8190 (
            .O(N__33157),
            .I(N__33149));
    LocalMux I__8189 (
            .O(N__33154),
            .I(M_this_external_address_qZ0Z_2));
    Odrv4 I__8188 (
            .O(N__33149),
            .I(M_this_external_address_qZ0Z_2));
    InMux I__8187 (
            .O(N__33144),
            .I(N__33141));
    LocalMux I__8186 (
            .O(N__33141),
            .I(N__33138));
    Span4Mux_h I__8185 (
            .O(N__33138),
            .I(N__33135));
    Odrv4 I__8184 (
            .O(N__33135),
            .I(un1_M_this_external_address_q_cry_2_THRU_CO));
    IoInMux I__8183 (
            .O(N__33132),
            .I(N__33129));
    LocalMux I__8182 (
            .O(N__33129),
            .I(N__33126));
    IoSpan4Mux I__8181 (
            .O(N__33126),
            .I(N__33121));
    InMux I__8180 (
            .O(N__33125),
            .I(N__33118));
    CascadeMux I__8179 (
            .O(N__33124),
            .I(N__33115));
    Span4Mux_s1_h I__8178 (
            .O(N__33121),
            .I(N__33112));
    LocalMux I__8177 (
            .O(N__33118),
            .I(N__33109));
    InMux I__8176 (
            .O(N__33115),
            .I(N__33106));
    Span4Mux_h I__8175 (
            .O(N__33112),
            .I(N__33101));
    Span4Mux_h I__8174 (
            .O(N__33109),
            .I(N__33101));
    LocalMux I__8173 (
            .O(N__33106),
            .I(M_this_external_address_qZ0Z_3));
    Odrv4 I__8172 (
            .O(N__33101),
            .I(M_this_external_address_qZ0Z_3));
    InMux I__8171 (
            .O(N__33096),
            .I(N__33093));
    LocalMux I__8170 (
            .O(N__33093),
            .I(N__33090));
    Span4Mux_v I__8169 (
            .O(N__33090),
            .I(N__33087));
    Odrv4 I__8168 (
            .O(N__33087),
            .I(un1_M_this_external_address_q_cry_3_THRU_CO));
    InMux I__8167 (
            .O(N__33084),
            .I(N__33079));
    IoInMux I__8166 (
            .O(N__33083),
            .I(N__33076));
    CascadeMux I__8165 (
            .O(N__33082),
            .I(N__33073));
    LocalMux I__8164 (
            .O(N__33079),
            .I(N__33070));
    LocalMux I__8163 (
            .O(N__33076),
            .I(N__33067));
    InMux I__8162 (
            .O(N__33073),
            .I(N__33064));
    Span4Mux_v I__8161 (
            .O(N__33070),
            .I(N__33061));
    Odrv12 I__8160 (
            .O(N__33067),
            .I(M_this_external_address_qZ0Z_4));
    LocalMux I__8159 (
            .O(N__33064),
            .I(M_this_external_address_qZ0Z_4));
    Odrv4 I__8158 (
            .O(N__33061),
            .I(M_this_external_address_qZ0Z_4));
    InMux I__8157 (
            .O(N__33054),
            .I(N__33051));
    LocalMux I__8156 (
            .O(N__33051),
            .I(N__33048));
    Span4Mux_v I__8155 (
            .O(N__33048),
            .I(N__33045));
    Odrv4 I__8154 (
            .O(N__33045),
            .I(un1_M_this_external_address_q_cry_4_THRU_CO));
    IoInMux I__8153 (
            .O(N__33042),
            .I(N__33039));
    LocalMux I__8152 (
            .O(N__33039),
            .I(N__33035));
    InMux I__8151 (
            .O(N__33038),
            .I(N__33031));
    Span4Mux_s1_h I__8150 (
            .O(N__33035),
            .I(N__33028));
    CascadeMux I__8149 (
            .O(N__33034),
            .I(N__33025));
    LocalMux I__8148 (
            .O(N__33031),
            .I(N__33022));
    Span4Mux_h I__8147 (
            .O(N__33028),
            .I(N__33019));
    InMux I__8146 (
            .O(N__33025),
            .I(N__33016));
    Span4Mux_h I__8145 (
            .O(N__33022),
            .I(N__33013));
    Odrv4 I__8144 (
            .O(N__33019),
            .I(M_this_external_address_qZ0Z_5));
    LocalMux I__8143 (
            .O(N__33016),
            .I(M_this_external_address_qZ0Z_5));
    Odrv4 I__8142 (
            .O(N__33013),
            .I(M_this_external_address_qZ0Z_5));
    CascadeMux I__8141 (
            .O(N__33006),
            .I(N__33003));
    InMux I__8140 (
            .O(N__33003),
            .I(N__33000));
    LocalMux I__8139 (
            .O(N__33000),
            .I(N__32997));
    Odrv12 I__8138 (
            .O(N__32997),
            .I(M_this_data_tmp_qZ0Z_23));
    InMux I__8137 (
            .O(N__32994),
            .I(N__32991));
    LocalMux I__8136 (
            .O(N__32991),
            .I(M_this_oam_ram_write_data_23));
    InMux I__8135 (
            .O(N__32988),
            .I(N__32982));
    InMux I__8134 (
            .O(N__32987),
            .I(N__32978));
    CascadeMux I__8133 (
            .O(N__32986),
            .I(N__32975));
    CascadeMux I__8132 (
            .O(N__32985),
            .I(N__32972));
    LocalMux I__8131 (
            .O(N__32982),
            .I(N__32968));
    InMux I__8130 (
            .O(N__32981),
            .I(N__32965));
    LocalMux I__8129 (
            .O(N__32978),
            .I(N__32962));
    InMux I__8128 (
            .O(N__32975),
            .I(N__32959));
    InMux I__8127 (
            .O(N__32972),
            .I(N__32956));
    CascadeMux I__8126 (
            .O(N__32971),
            .I(N__32951));
    Span4Mux_h I__8125 (
            .O(N__32968),
            .I(N__32946));
    LocalMux I__8124 (
            .O(N__32965),
            .I(N__32946));
    Span4Mux_v I__8123 (
            .O(N__32962),
            .I(N__32941));
    LocalMux I__8122 (
            .O(N__32959),
            .I(N__32941));
    LocalMux I__8121 (
            .O(N__32956),
            .I(N__32938));
    InMux I__8120 (
            .O(N__32955),
            .I(N__32935));
    InMux I__8119 (
            .O(N__32954),
            .I(N__32930));
    InMux I__8118 (
            .O(N__32951),
            .I(N__32930));
    Span4Mux_v I__8117 (
            .O(N__32946),
            .I(N__32927));
    Span4Mux_v I__8116 (
            .O(N__32941),
            .I(N__32923));
    Span4Mux_v I__8115 (
            .O(N__32938),
            .I(N__32918));
    LocalMux I__8114 (
            .O(N__32935),
            .I(N__32918));
    LocalMux I__8113 (
            .O(N__32930),
            .I(N__32913));
    Span4Mux_h I__8112 (
            .O(N__32927),
            .I(N__32909));
    InMux I__8111 (
            .O(N__32926),
            .I(N__32906));
    Span4Mux_h I__8110 (
            .O(N__32923),
            .I(N__32901));
    Span4Mux_v I__8109 (
            .O(N__32918),
            .I(N__32901));
    InMux I__8108 (
            .O(N__32917),
            .I(N__32898));
    InMux I__8107 (
            .O(N__32916),
            .I(N__32895));
    Span4Mux_v I__8106 (
            .O(N__32913),
            .I(N__32892));
    InMux I__8105 (
            .O(N__32912),
            .I(N__32889));
    Sp12to4 I__8104 (
            .O(N__32909),
            .I(N__32878));
    LocalMux I__8103 (
            .O(N__32906),
            .I(N__32878));
    Sp12to4 I__8102 (
            .O(N__32901),
            .I(N__32878));
    LocalMux I__8101 (
            .O(N__32898),
            .I(N__32878));
    LocalMux I__8100 (
            .O(N__32895),
            .I(N__32878));
    Span4Mux_h I__8099 (
            .O(N__32892),
            .I(N__32873));
    LocalMux I__8098 (
            .O(N__32889),
            .I(N__32873));
    Span12Mux_h I__8097 (
            .O(N__32878),
            .I(N__32868));
    Sp12to4 I__8096 (
            .O(N__32873),
            .I(N__32868));
    Odrv12 I__8095 (
            .O(N__32868),
            .I(port_data_c_1));
    InMux I__8094 (
            .O(N__32865),
            .I(N__32862));
    LocalMux I__8093 (
            .O(N__32862),
            .I(N_41_0));
    CascadeMux I__8092 (
            .O(N__32859),
            .I(N__32856));
    InMux I__8091 (
            .O(N__32856),
            .I(N__32853));
    LocalMux I__8090 (
            .O(N__32853),
            .I(N__32850));
    Odrv12 I__8089 (
            .O(N__32850),
            .I(M_this_data_tmp_qZ0Z_2));
    InMux I__8088 (
            .O(N__32847),
            .I(N__32844));
    LocalMux I__8087 (
            .O(N__32844),
            .I(N__32841));
    Span4Mux_h I__8086 (
            .O(N__32841),
            .I(N__32838));
    Odrv4 I__8085 (
            .O(N__32838),
            .I(un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0));
    InMux I__8084 (
            .O(N__32835),
            .I(N__32827));
    CascadeMux I__8083 (
            .O(N__32834),
            .I(N__32824));
    InMux I__8082 (
            .O(N__32833),
            .I(N__32820));
    CascadeMux I__8081 (
            .O(N__32832),
            .I(N__32817));
    InMux I__8080 (
            .O(N__32831),
            .I(N__32814));
    CascadeMux I__8079 (
            .O(N__32830),
            .I(N__32811));
    LocalMux I__8078 (
            .O(N__32827),
            .I(N__32808));
    InMux I__8077 (
            .O(N__32824),
            .I(N__32805));
    InMux I__8076 (
            .O(N__32823),
            .I(N__32802));
    LocalMux I__8075 (
            .O(N__32820),
            .I(N__32796));
    InMux I__8074 (
            .O(N__32817),
            .I(N__32793));
    LocalMux I__8073 (
            .O(N__32814),
            .I(N__32790));
    InMux I__8072 (
            .O(N__32811),
            .I(N__32787));
    Span4Mux_v I__8071 (
            .O(N__32808),
            .I(N__32782));
    LocalMux I__8070 (
            .O(N__32805),
            .I(N__32782));
    LocalMux I__8069 (
            .O(N__32802),
            .I(N__32779));
    InMux I__8068 (
            .O(N__32801),
            .I(N__32776));
    InMux I__8067 (
            .O(N__32800),
            .I(N__32773));
    InMux I__8066 (
            .O(N__32799),
            .I(N__32770));
    Span4Mux_v I__8065 (
            .O(N__32796),
            .I(N__32767));
    LocalMux I__8064 (
            .O(N__32793),
            .I(N__32764));
    Span4Mux_h I__8063 (
            .O(N__32790),
            .I(N__32759));
    LocalMux I__8062 (
            .O(N__32787),
            .I(N__32759));
    Span4Mux_h I__8061 (
            .O(N__32782),
            .I(N__32756));
    Span4Mux_v I__8060 (
            .O(N__32779),
            .I(N__32751));
    LocalMux I__8059 (
            .O(N__32776),
            .I(N__32751));
    LocalMux I__8058 (
            .O(N__32773),
            .I(N__32748));
    LocalMux I__8057 (
            .O(N__32770),
            .I(N__32745));
    Sp12to4 I__8056 (
            .O(N__32767),
            .I(N__32742));
    Span4Mux_v I__8055 (
            .O(N__32764),
            .I(N__32739));
    Span4Mux_v I__8054 (
            .O(N__32759),
            .I(N__32736));
    Span4Mux_v I__8053 (
            .O(N__32756),
            .I(N__32731));
    Span4Mux_h I__8052 (
            .O(N__32751),
            .I(N__32731));
    Span12Mux_h I__8051 (
            .O(N__32748),
            .I(N__32728));
    Span12Mux_v I__8050 (
            .O(N__32745),
            .I(N__32725));
    Span12Mux_h I__8049 (
            .O(N__32742),
            .I(N__32720));
    Sp12to4 I__8048 (
            .O(N__32739),
            .I(N__32720));
    Sp12to4 I__8047 (
            .O(N__32736),
            .I(N__32717));
    Span4Mux_v I__8046 (
            .O(N__32731),
            .I(N__32714));
    Span12Mux_v I__8045 (
            .O(N__32728),
            .I(N__32709));
    Span12Mux_h I__8044 (
            .O(N__32725),
            .I(N__32709));
    Span12Mux_h I__8043 (
            .O(N__32720),
            .I(N__32706));
    Span12Mux_h I__8042 (
            .O(N__32717),
            .I(N__32703));
    Span4Mux_h I__8041 (
            .O(N__32714),
            .I(N__32700));
    Odrv12 I__8040 (
            .O(N__32709),
            .I(port_data_c_3));
    Odrv12 I__8039 (
            .O(N__32706),
            .I(port_data_c_3));
    Odrv12 I__8038 (
            .O(N__32703),
            .I(port_data_c_3));
    Odrv4 I__8037 (
            .O(N__32700),
            .I(port_data_c_3));
    IoInMux I__8036 (
            .O(N__32691),
            .I(N__32688));
    LocalMux I__8035 (
            .O(N__32688),
            .I(N__32685));
    Span4Mux_s2_v I__8034 (
            .O(N__32685),
            .I(N__32681));
    InMux I__8033 (
            .O(N__32684),
            .I(N__32678));
    Span4Mux_v I__8032 (
            .O(N__32681),
            .I(N__32675));
    LocalMux I__8031 (
            .O(N__32678),
            .I(N__32672));
    Span4Mux_v I__8030 (
            .O(N__32675),
            .I(N__32669));
    Span4Mux_h I__8029 (
            .O(N__32672),
            .I(N__32666));
    Odrv4 I__8028 (
            .O(N__32669),
            .I(M_this_external_address_qZ0Z_11));
    Odrv4 I__8027 (
            .O(N__32666),
            .I(M_this_external_address_qZ0Z_11));
    InMux I__8026 (
            .O(N__32661),
            .I(N__32658));
    LocalMux I__8025 (
            .O(N__32658),
            .I(N__32655));
    Odrv4 I__8024 (
            .O(N__32655),
            .I(un1_M_this_external_address_q_cry_6_THRU_CO));
    IoInMux I__8023 (
            .O(N__32652),
            .I(N__32649));
    LocalMux I__8022 (
            .O(N__32649),
            .I(N__32646));
    IoSpan4Mux I__8021 (
            .O(N__32646),
            .I(N__32643));
    Span4Mux_s2_h I__8020 (
            .O(N__32643),
            .I(N__32640));
    Span4Mux_h I__8019 (
            .O(N__32640),
            .I(N__32637));
    Sp12to4 I__8018 (
            .O(N__32637),
            .I(N__32632));
    CascadeMux I__8017 (
            .O(N__32636),
            .I(N__32629));
    InMux I__8016 (
            .O(N__32635),
            .I(N__32626));
    Span12Mux_v I__8015 (
            .O(N__32632),
            .I(N__32623));
    InMux I__8014 (
            .O(N__32629),
            .I(N__32620));
    LocalMux I__8013 (
            .O(N__32626),
            .I(N__32617));
    Odrv12 I__8012 (
            .O(N__32623),
            .I(M_this_external_address_qZ0Z_7));
    LocalMux I__8011 (
            .O(N__32620),
            .I(M_this_external_address_qZ0Z_7));
    Odrv4 I__8010 (
            .O(N__32617),
            .I(M_this_external_address_qZ0Z_7));
    InMux I__8009 (
            .O(N__32610),
            .I(N__32607));
    LocalMux I__8008 (
            .O(N__32607),
            .I(N__32604));
    Span4Mux_h I__8007 (
            .O(N__32604),
            .I(N__32601));
    Odrv4 I__8006 (
            .O(N__32601),
            .I(un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0));
    CascadeMux I__8005 (
            .O(N__32598),
            .I(N__32595));
    InMux I__8004 (
            .O(N__32595),
            .I(N__32589));
    CascadeMux I__8003 (
            .O(N__32594),
            .I(N__32585));
    InMux I__8002 (
            .O(N__32593),
            .I(N__32582));
    CascadeMux I__8001 (
            .O(N__32592),
            .I(N__32579));
    LocalMux I__8000 (
            .O(N__32589),
            .I(N__32575));
    InMux I__7999 (
            .O(N__32588),
            .I(N__32572));
    InMux I__7998 (
            .O(N__32585),
            .I(N__32569));
    LocalMux I__7997 (
            .O(N__32582),
            .I(N__32565));
    InMux I__7996 (
            .O(N__32579),
            .I(N__32562));
    InMux I__7995 (
            .O(N__32578),
            .I(N__32559));
    Span4Mux_v I__7994 (
            .O(N__32575),
            .I(N__32556));
    LocalMux I__7993 (
            .O(N__32572),
            .I(N__32551));
    LocalMux I__7992 (
            .O(N__32569),
            .I(N__32551));
    CascadeMux I__7991 (
            .O(N__32568),
            .I(N__32548));
    Span4Mux_v I__7990 (
            .O(N__32565),
            .I(N__32544));
    LocalMux I__7989 (
            .O(N__32562),
            .I(N__32538));
    LocalMux I__7988 (
            .O(N__32559),
            .I(N__32538));
    Span4Mux_v I__7987 (
            .O(N__32556),
            .I(N__32533));
    Span4Mux_v I__7986 (
            .O(N__32551),
            .I(N__32533));
    InMux I__7985 (
            .O(N__32548),
            .I(N__32530));
    CascadeMux I__7984 (
            .O(N__32547),
            .I(N__32526));
    Span4Mux_v I__7983 (
            .O(N__32544),
            .I(N__32523));
    InMux I__7982 (
            .O(N__32543),
            .I(N__32520));
    Span4Mux_v I__7981 (
            .O(N__32538),
            .I(N__32513));
    Span4Mux_h I__7980 (
            .O(N__32533),
            .I(N__32513));
    LocalMux I__7979 (
            .O(N__32530),
            .I(N__32513));
    InMux I__7978 (
            .O(N__32529),
            .I(N__32510));
    InMux I__7977 (
            .O(N__32526),
            .I(N__32507));
    Sp12to4 I__7976 (
            .O(N__32523),
            .I(N__32502));
    LocalMux I__7975 (
            .O(N__32520),
            .I(N__32502));
    Sp12to4 I__7974 (
            .O(N__32513),
            .I(N__32499));
    LocalMux I__7973 (
            .O(N__32510),
            .I(N__32494));
    LocalMux I__7972 (
            .O(N__32507),
            .I(N__32494));
    Span12Mux_h I__7971 (
            .O(N__32502),
            .I(N__32489));
    Span12Mux_v I__7970 (
            .O(N__32499),
            .I(N__32489));
    Span12Mux_v I__7969 (
            .O(N__32494),
            .I(N__32486));
    Odrv12 I__7968 (
            .O(N__32489),
            .I(port_data_c_4));
    Odrv12 I__7967 (
            .O(N__32486),
            .I(port_data_c_4));
    IoInMux I__7966 (
            .O(N__32481),
            .I(N__32477));
    InMux I__7965 (
            .O(N__32480),
            .I(N__32474));
    LocalMux I__7964 (
            .O(N__32477),
            .I(N__32471));
    LocalMux I__7963 (
            .O(N__32474),
            .I(N__32468));
    Span12Mux_s6_h I__7962 (
            .O(N__32471),
            .I(N__32465));
    Span4Mux_h I__7961 (
            .O(N__32468),
            .I(N__32462));
    Odrv12 I__7960 (
            .O(N__32465),
            .I(M_this_external_address_qZ0Z_12));
    Odrv4 I__7959 (
            .O(N__32462),
            .I(M_this_external_address_qZ0Z_12));
    InMux I__7958 (
            .O(N__32457),
            .I(N__32454));
    LocalMux I__7957 (
            .O(N__32454),
            .I(N__32451));
    Span4Mux_h I__7956 (
            .O(N__32451),
            .I(N__32448));
    Odrv4 I__7955 (
            .O(N__32448),
            .I(un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0));
    IoInMux I__7954 (
            .O(N__32445),
            .I(N__32441));
    InMux I__7953 (
            .O(N__32444),
            .I(N__32438));
    LocalMux I__7952 (
            .O(N__32441),
            .I(N__32435));
    LocalMux I__7951 (
            .O(N__32438),
            .I(N__32432));
    Span12Mux_s6_h I__7950 (
            .O(N__32435),
            .I(N__32429));
    Span4Mux_h I__7949 (
            .O(N__32432),
            .I(N__32426));
    Odrv12 I__7948 (
            .O(N__32429),
            .I(M_this_external_address_qZ0Z_13));
    Odrv4 I__7947 (
            .O(N__32426),
            .I(M_this_external_address_qZ0Z_13));
    InMux I__7946 (
            .O(N__32421),
            .I(N__32418));
    LocalMux I__7945 (
            .O(N__32418),
            .I(N__32415));
    Span4Mux_h I__7944 (
            .O(N__32415),
            .I(N__32412));
    Odrv4 I__7943 (
            .O(N__32412),
            .I(un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0));
    CascadeMux I__7942 (
            .O(N__32409),
            .I(N__32404));
    InMux I__7941 (
            .O(N__32408),
            .I(N__32400));
    CascadeMux I__7940 (
            .O(N__32407),
            .I(N__32397));
    InMux I__7939 (
            .O(N__32404),
            .I(N__32394));
    CascadeMux I__7938 (
            .O(N__32403),
            .I(N__32390));
    LocalMux I__7937 (
            .O(N__32400),
            .I(N__32385));
    InMux I__7936 (
            .O(N__32397),
            .I(N__32382));
    LocalMux I__7935 (
            .O(N__32394),
            .I(N__32379));
    InMux I__7934 (
            .O(N__32393),
            .I(N__32374));
    InMux I__7933 (
            .O(N__32390),
            .I(N__32374));
    CascadeMux I__7932 (
            .O(N__32389),
            .I(N__32371));
    InMux I__7931 (
            .O(N__32388),
            .I(N__32368));
    Span4Mux_v I__7930 (
            .O(N__32385),
            .I(N__32365));
    LocalMux I__7929 (
            .O(N__32382),
            .I(N__32362));
    Span4Mux_h I__7928 (
            .O(N__32379),
            .I(N__32359));
    LocalMux I__7927 (
            .O(N__32374),
            .I(N__32356));
    InMux I__7926 (
            .O(N__32371),
            .I(N__32353));
    LocalMux I__7925 (
            .O(N__32368),
            .I(N__32349));
    Sp12to4 I__7924 (
            .O(N__32365),
            .I(N__32345));
    Span4Mux_v I__7923 (
            .O(N__32362),
            .I(N__32342));
    Span4Mux_v I__7922 (
            .O(N__32359),
            .I(N__32335));
    Span4Mux_h I__7921 (
            .O(N__32356),
            .I(N__32335));
    LocalMux I__7920 (
            .O(N__32353),
            .I(N__32335));
    CascadeMux I__7919 (
            .O(N__32352),
            .I(N__32332));
    Span4Mux_h I__7918 (
            .O(N__32349),
            .I(N__32328));
    InMux I__7917 (
            .O(N__32348),
            .I(N__32325));
    Span12Mux_h I__7916 (
            .O(N__32345),
            .I(N__32322));
    Span4Mux_v I__7915 (
            .O(N__32342),
            .I(N__32319));
    Span4Mux_h I__7914 (
            .O(N__32335),
            .I(N__32316));
    InMux I__7913 (
            .O(N__32332),
            .I(N__32313));
    InMux I__7912 (
            .O(N__32331),
            .I(N__32310));
    Span4Mux_v I__7911 (
            .O(N__32328),
            .I(N__32305));
    LocalMux I__7910 (
            .O(N__32325),
            .I(N__32305));
    Span12Mux_h I__7909 (
            .O(N__32322),
            .I(N__32302));
    Span4Mux_v I__7908 (
            .O(N__32319),
            .I(N__32299));
    Sp12to4 I__7907 (
            .O(N__32316),
            .I(N__32290));
    LocalMux I__7906 (
            .O(N__32313),
            .I(N__32290));
    LocalMux I__7905 (
            .O(N__32310),
            .I(N__32290));
    Sp12to4 I__7904 (
            .O(N__32305),
            .I(N__32290));
    Span12Mux_v I__7903 (
            .O(N__32302),
            .I(N__32287));
    Sp12to4 I__7902 (
            .O(N__32299),
            .I(N__32282));
    Span12Mux_v I__7901 (
            .O(N__32290),
            .I(N__32282));
    Odrv12 I__7900 (
            .O(N__32287),
            .I(port_data_c_6));
    Odrv12 I__7899 (
            .O(N__32282),
            .I(port_data_c_6));
    IoInMux I__7898 (
            .O(N__32277),
            .I(N__32274));
    LocalMux I__7897 (
            .O(N__32274),
            .I(N__32271));
    IoSpan4Mux I__7896 (
            .O(N__32271),
            .I(N__32267));
    InMux I__7895 (
            .O(N__32270),
            .I(N__32264));
    Span4Mux_s2_h I__7894 (
            .O(N__32267),
            .I(N__32261));
    LocalMux I__7893 (
            .O(N__32264),
            .I(N__32258));
    Span4Mux_v I__7892 (
            .O(N__32261),
            .I(N__32255));
    Span4Mux_v I__7891 (
            .O(N__32258),
            .I(N__32252));
    Odrv4 I__7890 (
            .O(N__32255),
            .I(M_this_external_address_qZ0Z_14));
    Odrv4 I__7889 (
            .O(N__32252),
            .I(M_this_external_address_qZ0Z_14));
    InMux I__7888 (
            .O(N__32247),
            .I(N__32244));
    LocalMux I__7887 (
            .O(N__32244),
            .I(N_63_0));
    InMux I__7886 (
            .O(N__32241),
            .I(N__32238));
    LocalMux I__7885 (
            .O(N__32238),
            .I(N_75_0));
    InMux I__7884 (
            .O(N__32235),
            .I(N__32232));
    LocalMux I__7883 (
            .O(N__32232),
            .I(M_this_oam_ram_write_data_11));
    CascadeMux I__7882 (
            .O(N__32229),
            .I(N__32226));
    InMux I__7881 (
            .O(N__32226),
            .I(N__32223));
    LocalMux I__7880 (
            .O(N__32223),
            .I(M_this_data_tmp_qZ0Z_11));
    InMux I__7879 (
            .O(N__32220),
            .I(N__32217));
    LocalMux I__7878 (
            .O(N__32217),
            .I(N__32214));
    Odrv4 I__7877 (
            .O(N__32214),
            .I(M_this_data_tmp_qZ0Z_12));
    CascadeMux I__7876 (
            .O(N__32211),
            .I(N__32208));
    InMux I__7875 (
            .O(N__32208),
            .I(N__32205));
    LocalMux I__7874 (
            .O(N__32205),
            .I(M_this_data_tmp_qZ0Z_9));
    CascadeMux I__7873 (
            .O(N__32202),
            .I(N__32199));
    InMux I__7872 (
            .O(N__32199),
            .I(N__32196));
    LocalMux I__7871 (
            .O(N__32196),
            .I(N__32193));
    Odrv4 I__7870 (
            .O(N__32193),
            .I(M_this_data_tmp_qZ0Z_14));
    CEMux I__7869 (
            .O(N__32190),
            .I(N__32185));
    CEMux I__7868 (
            .O(N__32189),
            .I(N__32180));
    CEMux I__7867 (
            .O(N__32188),
            .I(N__32177));
    LocalMux I__7866 (
            .O(N__32185),
            .I(N__32174));
    CEMux I__7865 (
            .O(N__32184),
            .I(N__32171));
    CEMux I__7864 (
            .O(N__32183),
            .I(N__32168));
    LocalMux I__7863 (
            .O(N__32180),
            .I(N__32165));
    LocalMux I__7862 (
            .O(N__32177),
            .I(N__32162));
    Span4Mux_v I__7861 (
            .O(N__32174),
            .I(N__32159));
    LocalMux I__7860 (
            .O(N__32171),
            .I(N__32156));
    LocalMux I__7859 (
            .O(N__32168),
            .I(N__32153));
    Span4Mux_h I__7858 (
            .O(N__32165),
            .I(N__32150));
    Span4Mux_v I__7857 (
            .O(N__32162),
            .I(N__32143));
    Span4Mux_h I__7856 (
            .O(N__32159),
            .I(N__32143));
    Span4Mux_v I__7855 (
            .O(N__32156),
            .I(N__32143));
    Span4Mux_h I__7854 (
            .O(N__32153),
            .I(N__32140));
    Sp12to4 I__7853 (
            .O(N__32150),
            .I(N__32137));
    Span4Mux_h I__7852 (
            .O(N__32143),
            .I(N__32134));
    Odrv4 I__7851 (
            .O(N__32140),
            .I(N_1134_0));
    Odrv12 I__7850 (
            .O(N__32137),
            .I(N_1134_0));
    Odrv4 I__7849 (
            .O(N__32134),
            .I(N_1134_0));
    InMux I__7848 (
            .O(N__32127),
            .I(N__32124));
    LocalMux I__7847 (
            .O(N__32124),
            .I(N_39_0));
    InMux I__7846 (
            .O(N__32121),
            .I(N__32118));
    LocalMux I__7845 (
            .O(N__32118),
            .I(M_this_oam_ram_write_data_27));
    InMux I__7844 (
            .O(N__32115),
            .I(N__32112));
    LocalMux I__7843 (
            .O(N__32112),
            .I(M_this_oam_ram_write_data_8));
    CascadeMux I__7842 (
            .O(N__32109),
            .I(N__32106));
    InMux I__7841 (
            .O(N__32106),
            .I(N__32103));
    LocalMux I__7840 (
            .O(N__32103),
            .I(M_this_data_tmp_qZ0Z_8));
    InMux I__7839 (
            .O(N__32100),
            .I(N__32097));
    LocalMux I__7838 (
            .O(N__32097),
            .I(N_79_0));
    CascadeMux I__7837 (
            .O(N__32094),
            .I(N__32091));
    InMux I__7836 (
            .O(N__32091),
            .I(N__32088));
    LocalMux I__7835 (
            .O(N__32088),
            .I(M_this_data_tmp_qZ0Z_0));
    InMux I__7834 (
            .O(N__32085),
            .I(N__32082));
    LocalMux I__7833 (
            .O(N__32082),
            .I(N__32079));
    Span4Mux_v I__7832 (
            .O(N__32079),
            .I(N__32076));
    Odrv4 I__7831 (
            .O(N__32076),
            .I(N_43_0));
    InMux I__7830 (
            .O(N__32073),
            .I(N__32070));
    LocalMux I__7829 (
            .O(N__32070),
            .I(N__32067));
    Odrv4 I__7828 (
            .O(N__32067),
            .I(N_77_0));
    InMux I__7827 (
            .O(N__32064),
            .I(N__32061));
    LocalMux I__7826 (
            .O(N__32061),
            .I(M_this_data_tmp_qZ0Z_1));
    InMux I__7825 (
            .O(N__32058),
            .I(N__32055));
    LocalMux I__7824 (
            .O(N__32055),
            .I(N_58_0));
    InMux I__7823 (
            .O(N__32052),
            .I(N__32049));
    LocalMux I__7822 (
            .O(N__32049),
            .I(M_this_oam_ram_write_data_14));
    InMux I__7821 (
            .O(N__32046),
            .I(bfn_24_23_0_));
    IoInMux I__7820 (
            .O(N__32043),
            .I(N__32040));
    LocalMux I__7819 (
            .O(N__32040),
            .I(N__32037));
    Span4Mux_s1_v I__7818 (
            .O(N__32037),
            .I(N__32034));
    Span4Mux_v I__7817 (
            .O(N__32034),
            .I(N__32030));
    InMux I__7816 (
            .O(N__32033),
            .I(N__32027));
    Span4Mux_v I__7815 (
            .O(N__32030),
            .I(N__32022));
    LocalMux I__7814 (
            .O(N__32027),
            .I(N__32022));
    Odrv4 I__7813 (
            .O(N__32022),
            .I(M_this_external_address_qZ0Z_9));
    InMux I__7812 (
            .O(N__32019),
            .I(N__32016));
    LocalMux I__7811 (
            .O(N__32016),
            .I(N__32013));
    Odrv12 I__7810 (
            .O(N__32013),
            .I(un1_M_this_external_address_q_cry_8_c_RNI09PBZ0));
    InMux I__7809 (
            .O(N__32010),
            .I(un1_M_this_external_address_q_cry_8));
    InMux I__7808 (
            .O(N__32007),
            .I(un1_M_this_external_address_q_cry_9));
    InMux I__7807 (
            .O(N__32004),
            .I(un1_M_this_external_address_q_cry_10));
    InMux I__7806 (
            .O(N__32001),
            .I(un1_M_this_external_address_q_cry_11));
    InMux I__7805 (
            .O(N__31998),
            .I(un1_M_this_external_address_q_cry_12));
    InMux I__7804 (
            .O(N__31995),
            .I(un1_M_this_external_address_q_cry_13));
    InMux I__7803 (
            .O(N__31992),
            .I(un1_M_this_external_address_q_cry_14));
    InMux I__7802 (
            .O(N__31989),
            .I(N__31985));
    InMux I__7801 (
            .O(N__31988),
            .I(N__31980));
    LocalMux I__7800 (
            .O(N__31985),
            .I(N__31977));
    InMux I__7799 (
            .O(N__31984),
            .I(N__31974));
    InMux I__7798 (
            .O(N__31983),
            .I(N__31971));
    LocalMux I__7797 (
            .O(N__31980),
            .I(N__31964));
    Span4Mux_v I__7796 (
            .O(N__31977),
            .I(N__31961));
    LocalMux I__7795 (
            .O(N__31974),
            .I(N__31958));
    LocalMux I__7794 (
            .O(N__31971),
            .I(N__31955));
    InMux I__7793 (
            .O(N__31970),
            .I(N__31952));
    InMux I__7792 (
            .O(N__31969),
            .I(N__31949));
    InMux I__7791 (
            .O(N__31968),
            .I(N__31944));
    InMux I__7790 (
            .O(N__31967),
            .I(N__31941));
    Span4Mux_v I__7789 (
            .O(N__31964),
            .I(N__31937));
    Span4Mux_v I__7788 (
            .O(N__31961),
            .I(N__31932));
    Span4Mux_v I__7787 (
            .O(N__31958),
            .I(N__31932));
    Span4Mux_v I__7786 (
            .O(N__31955),
            .I(N__31929));
    LocalMux I__7785 (
            .O(N__31952),
            .I(N__31924));
    LocalMux I__7784 (
            .O(N__31949),
            .I(N__31924));
    InMux I__7783 (
            .O(N__31948),
            .I(N__31921));
    InMux I__7782 (
            .O(N__31947),
            .I(N__31918));
    LocalMux I__7781 (
            .O(N__31944),
            .I(N__31915));
    LocalMux I__7780 (
            .O(N__31941),
            .I(N__31912));
    InMux I__7779 (
            .O(N__31940),
            .I(N__31909));
    Odrv4 I__7778 (
            .O(N__31937),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv4 I__7777 (
            .O(N__31932),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv4 I__7776 (
            .O(N__31929),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv12 I__7775 (
            .O(N__31924),
            .I(M_this_sprites_address_qZ0Z_12));
    LocalMux I__7774 (
            .O(N__31921),
            .I(M_this_sprites_address_qZ0Z_12));
    LocalMux I__7773 (
            .O(N__31918),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv4 I__7772 (
            .O(N__31915),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv4 I__7771 (
            .O(N__31912),
            .I(M_this_sprites_address_qZ0Z_12));
    LocalMux I__7770 (
            .O(N__31909),
            .I(M_this_sprites_address_qZ0Z_12));
    InMux I__7769 (
            .O(N__31890),
            .I(N__31887));
    LocalMux I__7768 (
            .O(N__31887),
            .I(N__31882));
    InMux I__7767 (
            .O(N__31886),
            .I(N__31879));
    InMux I__7766 (
            .O(N__31885),
            .I(N__31876));
    Span4Mux_v I__7765 (
            .O(N__31882),
            .I(N__31870));
    LocalMux I__7764 (
            .O(N__31879),
            .I(N__31870));
    LocalMux I__7763 (
            .O(N__31876),
            .I(N__31867));
    InMux I__7762 (
            .O(N__31875),
            .I(N__31864));
    Span4Mux_h I__7761 (
            .O(N__31870),
            .I(N__31858));
    Span4Mux_h I__7760 (
            .O(N__31867),
            .I(N__31853));
    LocalMux I__7759 (
            .O(N__31864),
            .I(N__31853));
    InMux I__7758 (
            .O(N__31863),
            .I(N__31850));
    InMux I__7757 (
            .O(N__31862),
            .I(N__31847));
    CascadeMux I__7756 (
            .O(N__31861),
            .I(N__31840));
    Span4Mux_v I__7755 (
            .O(N__31858),
            .I(N__31835));
    Span4Mux_h I__7754 (
            .O(N__31853),
            .I(N__31835));
    LocalMux I__7753 (
            .O(N__31850),
            .I(N__31830));
    LocalMux I__7752 (
            .O(N__31847),
            .I(N__31830));
    InMux I__7751 (
            .O(N__31846),
            .I(N__31827));
    InMux I__7750 (
            .O(N__31845),
            .I(N__31824));
    InMux I__7749 (
            .O(N__31844),
            .I(N__31821));
    InMux I__7748 (
            .O(N__31843),
            .I(N__31818));
    InMux I__7747 (
            .O(N__31840),
            .I(N__31815));
    Odrv4 I__7746 (
            .O(N__31835),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv12 I__7745 (
            .O(N__31830),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__7744 (
            .O(N__31827),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__7743 (
            .O(N__31824),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__7742 (
            .O(N__31821),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__7741 (
            .O(N__31818),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__7740 (
            .O(N__31815),
            .I(M_this_sprites_address_qZ0Z_11));
    CascadeMux I__7739 (
            .O(N__31800),
            .I(N__31796));
    CascadeMux I__7738 (
            .O(N__31799),
            .I(N__31792));
    InMux I__7737 (
            .O(N__31796),
            .I(N__31787));
    CascadeMux I__7736 (
            .O(N__31795),
            .I(N__31784));
    InMux I__7735 (
            .O(N__31792),
            .I(N__31780));
    CascadeMux I__7734 (
            .O(N__31791),
            .I(N__31776));
    CascadeMux I__7733 (
            .O(N__31790),
            .I(N__31773));
    LocalMux I__7732 (
            .O(N__31787),
            .I(N__31770));
    InMux I__7731 (
            .O(N__31784),
            .I(N__31767));
    InMux I__7730 (
            .O(N__31783),
            .I(N__31764));
    LocalMux I__7729 (
            .O(N__31780),
            .I(N__31761));
    CascadeMux I__7728 (
            .O(N__31779),
            .I(N__31758));
    InMux I__7727 (
            .O(N__31776),
            .I(N__31755));
    InMux I__7726 (
            .O(N__31773),
            .I(N__31750));
    Span4Mux_v I__7725 (
            .O(N__31770),
            .I(N__31746));
    LocalMux I__7724 (
            .O(N__31767),
            .I(N__31743));
    LocalMux I__7723 (
            .O(N__31764),
            .I(N__31740));
    Span4Mux_v I__7722 (
            .O(N__31761),
            .I(N__31737));
    InMux I__7721 (
            .O(N__31758),
            .I(N__31734));
    LocalMux I__7720 (
            .O(N__31755),
            .I(N__31731));
    CascadeMux I__7719 (
            .O(N__31754),
            .I(N__31728));
    CascadeMux I__7718 (
            .O(N__31753),
            .I(N__31725));
    LocalMux I__7717 (
            .O(N__31750),
            .I(N__31721));
    InMux I__7716 (
            .O(N__31749),
            .I(N__31718));
    Span4Mux_v I__7715 (
            .O(N__31746),
            .I(N__31711));
    Span4Mux_v I__7714 (
            .O(N__31743),
            .I(N__31711));
    Span4Mux_h I__7713 (
            .O(N__31740),
            .I(N__31711));
    Span4Mux_v I__7712 (
            .O(N__31737),
            .I(N__31708));
    LocalMux I__7711 (
            .O(N__31734),
            .I(N__31705));
    Span4Mux_v I__7710 (
            .O(N__31731),
            .I(N__31702));
    InMux I__7709 (
            .O(N__31728),
            .I(N__31699));
    InMux I__7708 (
            .O(N__31725),
            .I(N__31696));
    InMux I__7707 (
            .O(N__31724),
            .I(N__31693));
    Span4Mux_v I__7706 (
            .O(N__31721),
            .I(N__31686));
    LocalMux I__7705 (
            .O(N__31718),
            .I(N__31686));
    Span4Mux_h I__7704 (
            .O(N__31711),
            .I(N__31686));
    Odrv4 I__7703 (
            .O(N__31708),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv12 I__7702 (
            .O(N__31705),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__7701 (
            .O(N__31702),
            .I(M_this_sprites_address_qZ0Z_13));
    LocalMux I__7700 (
            .O(N__31699),
            .I(M_this_sprites_address_qZ0Z_13));
    LocalMux I__7699 (
            .O(N__31696),
            .I(M_this_sprites_address_qZ0Z_13));
    LocalMux I__7698 (
            .O(N__31693),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__7697 (
            .O(N__31686),
            .I(M_this_sprites_address_qZ0Z_13));
    InMux I__7696 (
            .O(N__31671),
            .I(N__31668));
    LocalMux I__7695 (
            .O(N__31668),
            .I(N__31664));
    InMux I__7694 (
            .O(N__31667),
            .I(N__31661));
    Span4Mux_v I__7693 (
            .O(N__31664),
            .I(N__31656));
    LocalMux I__7692 (
            .O(N__31661),
            .I(N__31653));
    InMux I__7691 (
            .O(N__31660),
            .I(N__31650));
    InMux I__7690 (
            .O(N__31659),
            .I(N__31646));
    Span4Mux_v I__7689 (
            .O(N__31656),
            .I(N__31640));
    Span4Mux_v I__7688 (
            .O(N__31653),
            .I(N__31640));
    LocalMux I__7687 (
            .O(N__31650),
            .I(N__31637));
    InMux I__7686 (
            .O(N__31649),
            .I(N__31634));
    LocalMux I__7685 (
            .O(N__31646),
            .I(N__31631));
    InMux I__7684 (
            .O(N__31645),
            .I(N__31628));
    Span4Mux_h I__7683 (
            .O(N__31640),
            .I(N__31621));
    Span4Mux_v I__7682 (
            .O(N__31637),
            .I(N__31621));
    LocalMux I__7681 (
            .O(N__31634),
            .I(N__31618));
    Span4Mux_v I__7680 (
            .O(N__31631),
            .I(N__31615));
    LocalMux I__7679 (
            .O(N__31628),
            .I(N__31612));
    InMux I__7678 (
            .O(N__31627),
            .I(N__31609));
    InMux I__7677 (
            .O(N__31626),
            .I(N__31606));
    Odrv4 I__7676 (
            .O(N__31621),
            .I(M_this_sprites_ram_write_en_0_0));
    Odrv12 I__7675 (
            .O(N__31618),
            .I(M_this_sprites_ram_write_en_0_0));
    Odrv4 I__7674 (
            .O(N__31615),
            .I(M_this_sprites_ram_write_en_0_0));
    Odrv4 I__7673 (
            .O(N__31612),
            .I(M_this_sprites_ram_write_en_0_0));
    LocalMux I__7672 (
            .O(N__31609),
            .I(M_this_sprites_ram_write_en_0_0));
    LocalMux I__7671 (
            .O(N__31606),
            .I(M_this_sprites_ram_write_en_0_0));
    CEMux I__7670 (
            .O(N__31593),
            .I(N__31589));
    CEMux I__7669 (
            .O(N__31592),
            .I(N__31586));
    LocalMux I__7668 (
            .O(N__31589),
            .I(N__31581));
    LocalMux I__7667 (
            .O(N__31586),
            .I(N__31581));
    Odrv4 I__7666 (
            .O(N__31581),
            .I(\this_sprites_ram.mem_WE_2 ));
    InMux I__7665 (
            .O(N__31578),
            .I(N__31575));
    LocalMux I__7664 (
            .O(N__31575),
            .I(N__31572));
    Span4Mux_v I__7663 (
            .O(N__31572),
            .I(N__31569));
    Odrv4 I__7662 (
            .O(N__31569),
            .I(M_this_oam_ram_write_data_30));
    InMux I__7661 (
            .O(N__31566),
            .I(un1_M_this_external_address_q_cry_0));
    InMux I__7660 (
            .O(N__31563),
            .I(un1_M_this_external_address_q_cry_1));
    InMux I__7659 (
            .O(N__31560),
            .I(un1_M_this_external_address_q_cry_2));
    InMux I__7658 (
            .O(N__31557),
            .I(un1_M_this_external_address_q_cry_3));
    InMux I__7657 (
            .O(N__31554),
            .I(un1_M_this_external_address_q_cry_4));
    InMux I__7656 (
            .O(N__31551),
            .I(un1_M_this_external_address_q_cry_5));
    InMux I__7655 (
            .O(N__31548),
            .I(un1_M_this_external_address_q_cry_6));
    InMux I__7654 (
            .O(N__31545),
            .I(N__31542));
    LocalMux I__7653 (
            .O(N__31542),
            .I(N__31537));
    InMux I__7652 (
            .O(N__31541),
            .I(N__31529));
    InMux I__7651 (
            .O(N__31540),
            .I(N__31529));
    Span4Mux_h I__7650 (
            .O(N__31537),
            .I(N__31526));
    InMux I__7649 (
            .O(N__31536),
            .I(N__31519));
    InMux I__7648 (
            .O(N__31535),
            .I(N__31519));
    InMux I__7647 (
            .O(N__31534),
            .I(N__31519));
    LocalMux I__7646 (
            .O(N__31529),
            .I(N__31516));
    Odrv4 I__7645 (
            .O(N__31526),
            .I(M_this_oam_ram_read_data_19));
    LocalMux I__7644 (
            .O(N__31519),
            .I(M_this_oam_ram_read_data_19));
    Odrv4 I__7643 (
            .O(N__31516),
            .I(M_this_oam_ram_read_data_19));
    CascadeMux I__7642 (
            .O(N__31509),
            .I(N__31506));
    InMux I__7641 (
            .O(N__31506),
            .I(N__31503));
    LocalMux I__7640 (
            .O(N__31503),
            .I(N__31500));
    Span4Mux_v I__7639 (
            .O(N__31500),
            .I(N__31497));
    Odrv4 I__7638 (
            .O(N__31497),
            .I(M_this_oam_ram_read_data_i_19));
    InMux I__7637 (
            .O(N__31494),
            .I(N__31491));
    LocalMux I__7636 (
            .O(N__31491),
            .I(M_this_data_tmp_qZ0Z_16));
    CascadeMux I__7635 (
            .O(N__31488),
            .I(N__31485));
    InMux I__7634 (
            .O(N__31485),
            .I(N__31482));
    LocalMux I__7633 (
            .O(N__31482),
            .I(M_this_data_tmp_qZ0Z_19));
    CascadeMux I__7632 (
            .O(N__31479),
            .I(N__31476));
    InMux I__7631 (
            .O(N__31476),
            .I(N__31473));
    LocalMux I__7630 (
            .O(N__31473),
            .I(M_this_data_tmp_qZ0Z_18));
    InMux I__7629 (
            .O(N__31470),
            .I(N__31467));
    LocalMux I__7628 (
            .O(N__31467),
            .I(M_this_data_tmp_qZ0Z_22));
    CascadeMux I__7627 (
            .O(N__31464),
            .I(N__31461));
    InMux I__7626 (
            .O(N__31461),
            .I(N__31458));
    LocalMux I__7625 (
            .O(N__31458),
            .I(M_this_data_tmp_qZ0Z_17));
    InMux I__7624 (
            .O(N__31455),
            .I(N__31452));
    LocalMux I__7623 (
            .O(N__31452),
            .I(N_54_0));
    CEMux I__7622 (
            .O(N__31449),
            .I(N__31446));
    LocalMux I__7621 (
            .O(N__31446),
            .I(N__31442));
    CEMux I__7620 (
            .O(N__31445),
            .I(N__31439));
    Span4Mux_v I__7619 (
            .O(N__31442),
            .I(N__31433));
    LocalMux I__7618 (
            .O(N__31439),
            .I(N__31433));
    CEMux I__7617 (
            .O(N__31438),
            .I(N__31430));
    Span4Mux_h I__7616 (
            .O(N__31433),
            .I(N__31427));
    LocalMux I__7615 (
            .O(N__31430),
            .I(N__31424));
    Span4Mux_h I__7614 (
            .O(N__31427),
            .I(N__31421));
    Odrv12 I__7613 (
            .O(N__31424),
            .I(N_1126_0));
    Odrv4 I__7612 (
            .O(N__31421),
            .I(N_1126_0));
    CascadeMux I__7611 (
            .O(N__31416),
            .I(N__31412));
    InMux I__7610 (
            .O(N__31415),
            .I(N__31409));
    InMux I__7609 (
            .O(N__31412),
            .I(N__31406));
    LocalMux I__7608 (
            .O(N__31409),
            .I(N__31401));
    LocalMux I__7607 (
            .O(N__31406),
            .I(N__31401));
    Span4Mux_v I__7606 (
            .O(N__31401),
            .I(N__31398));
    Odrv4 I__7605 (
            .O(N__31398),
            .I(M_this_oam_ram_read_data_23));
    CascadeMux I__7604 (
            .O(N__31395),
            .I(\this_ppu.un1_oam_data_c2_cascade_ ));
    InMux I__7603 (
            .O(N__31392),
            .I(N__31389));
    LocalMux I__7602 (
            .O(N__31389),
            .I(N__31386));
    Span4Mux_h I__7601 (
            .O(N__31386),
            .I(N__31383));
    Odrv4 I__7600 (
            .O(N__31383),
            .I(\this_ppu.un1_M_vaddress_q_3_7 ));
    InMux I__7599 (
            .O(N__31380),
            .I(N__31377));
    LocalMux I__7598 (
            .O(N__31377),
            .I(M_this_oam_ram_write_data_22));
    InMux I__7597 (
            .O(N__31374),
            .I(N__31369));
    InMux I__7596 (
            .O(N__31373),
            .I(N__31366));
    CascadeMux I__7595 (
            .O(N__31372),
            .I(N__31363));
    LocalMux I__7594 (
            .O(N__31369),
            .I(N__31358));
    LocalMux I__7593 (
            .O(N__31366),
            .I(N__31358));
    InMux I__7592 (
            .O(N__31363),
            .I(N__31355));
    Span4Mux_v I__7591 (
            .O(N__31358),
            .I(N__31352));
    LocalMux I__7590 (
            .O(N__31355),
            .I(M_this_oam_ram_read_data_22));
    Odrv4 I__7589 (
            .O(N__31352),
            .I(M_this_oam_ram_read_data_22));
    CascadeMux I__7588 (
            .O(N__31347),
            .I(N__31344));
    InMux I__7587 (
            .O(N__31344),
            .I(N__31341));
    LocalMux I__7586 (
            .O(N__31341),
            .I(N__31338));
    Span4Mux_h I__7585 (
            .O(N__31338),
            .I(N__31335));
    Odrv4 I__7584 (
            .O(N__31335),
            .I(\this_ppu.un1_M_vaddress_q_3_6 ));
    InMux I__7583 (
            .O(N__31332),
            .I(N__31329));
    LocalMux I__7582 (
            .O(N__31329),
            .I(M_this_oam_ram_write_data_31));
    InMux I__7581 (
            .O(N__31326),
            .I(N__31323));
    LocalMux I__7580 (
            .O(N__31323),
            .I(N_52_0));
    InMux I__7579 (
            .O(N__31320),
            .I(N__31317));
    LocalMux I__7578 (
            .O(N__31317),
            .I(M_this_oam_ram_write_data_16));
    CEMux I__7577 (
            .O(N__31314),
            .I(N__31311));
    LocalMux I__7576 (
            .O(N__31311),
            .I(N__31307));
    CEMux I__7575 (
            .O(N__31310),
            .I(N__31304));
    Span4Mux_h I__7574 (
            .O(N__31307),
            .I(N__31299));
    LocalMux I__7573 (
            .O(N__31304),
            .I(N__31299));
    Span4Mux_v I__7572 (
            .O(N__31299),
            .I(N__31296));
    Span4Mux_v I__7571 (
            .O(N__31296),
            .I(N__31293));
    Odrv4 I__7570 (
            .O(N__31293),
            .I(N_158_0));
    InMux I__7569 (
            .O(N__31290),
            .I(N__31286));
    InMux I__7568 (
            .O(N__31289),
            .I(N__31283));
    LocalMux I__7567 (
            .O(N__31286),
            .I(N__31279));
    LocalMux I__7566 (
            .O(N__31283),
            .I(N__31275));
    InMux I__7565 (
            .O(N__31282),
            .I(N__31272));
    Span4Mux_h I__7564 (
            .O(N__31279),
            .I(N__31269));
    InMux I__7563 (
            .O(N__31278),
            .I(N__31266));
    Odrv4 I__7562 (
            .O(N__31275),
            .I(M_this_oam_ram_read_data_21));
    LocalMux I__7561 (
            .O(N__31272),
            .I(M_this_oam_ram_read_data_21));
    Odrv4 I__7560 (
            .O(N__31269),
            .I(M_this_oam_ram_read_data_21));
    LocalMux I__7559 (
            .O(N__31266),
            .I(M_this_oam_ram_read_data_21));
    InMux I__7558 (
            .O(N__31257),
            .I(N__31253));
    CascadeMux I__7557 (
            .O(N__31256),
            .I(N__31250));
    LocalMux I__7556 (
            .O(N__31253),
            .I(N__31244));
    InMux I__7555 (
            .O(N__31250),
            .I(N__31239));
    InMux I__7554 (
            .O(N__31249),
            .I(N__31239));
    InMux I__7553 (
            .O(N__31248),
            .I(N__31234));
    InMux I__7552 (
            .O(N__31247),
            .I(N__31234));
    Span4Mux_h I__7551 (
            .O(N__31244),
            .I(N__31231));
    LocalMux I__7550 (
            .O(N__31239),
            .I(N__31228));
    LocalMux I__7549 (
            .O(N__31234),
            .I(M_this_oam_ram_read_data_20));
    Odrv4 I__7548 (
            .O(N__31231),
            .I(M_this_oam_ram_read_data_20));
    Odrv4 I__7547 (
            .O(N__31228),
            .I(M_this_oam_ram_read_data_20));
    CascadeMux I__7546 (
            .O(N__31221),
            .I(N__31218));
    InMux I__7545 (
            .O(N__31218),
            .I(N__31215));
    LocalMux I__7544 (
            .O(N__31215),
            .I(N__31212));
    Span4Mux_h I__7543 (
            .O(N__31212),
            .I(N__31209));
    Odrv4 I__7542 (
            .O(N__31209),
            .I(\this_ppu.un1_M_vaddress_q_3_5 ));
    CascadeMux I__7541 (
            .O(N__31206),
            .I(N__31202));
    CascadeMux I__7540 (
            .O(N__31205),
            .I(N__31198));
    InMux I__7539 (
            .O(N__31202),
            .I(N__31195));
    InMux I__7538 (
            .O(N__31201),
            .I(N__31192));
    InMux I__7537 (
            .O(N__31198),
            .I(N__31189));
    LocalMux I__7536 (
            .O(N__31195),
            .I(N__31186));
    LocalMux I__7535 (
            .O(N__31192),
            .I(N__31183));
    LocalMux I__7534 (
            .O(N__31189),
            .I(N__31180));
    Span4Mux_h I__7533 (
            .O(N__31186),
            .I(N__31177));
    Span4Mux_v I__7532 (
            .O(N__31183),
            .I(N__31172));
    Span4Mux_h I__7531 (
            .O(N__31180),
            .I(N__31172));
    Odrv4 I__7530 (
            .O(N__31177),
            .I(M_this_oam_ram_read_data_17));
    Odrv4 I__7529 (
            .O(N__31172),
            .I(M_this_oam_ram_read_data_17));
    InMux I__7528 (
            .O(N__31167),
            .I(N__31164));
    LocalMux I__7527 (
            .O(N__31164),
            .I(M_this_oam_ram_read_data_i_17));
    InMux I__7526 (
            .O(N__31161),
            .I(N__31158));
    LocalMux I__7525 (
            .O(N__31158),
            .I(N__31155));
    Span4Mux_h I__7524 (
            .O(N__31155),
            .I(N__31152));
    Span4Mux_h I__7523 (
            .O(N__31152),
            .I(N__31149));
    Span4Mux_h I__7522 (
            .O(N__31149),
            .I(N__31145));
    InMux I__7521 (
            .O(N__31148),
            .I(N__31142));
    Odrv4 I__7520 (
            .O(N__31145),
            .I(M_this_oam_ram_read_data_2));
    LocalMux I__7519 (
            .O(N__31142),
            .I(M_this_oam_ram_read_data_2));
    InMux I__7518 (
            .O(N__31137),
            .I(N__31134));
    LocalMux I__7517 (
            .O(N__31134),
            .I(N__31131));
    Span4Mux_v I__7516 (
            .O(N__31131),
            .I(N__31128));
    Sp12to4 I__7515 (
            .O(N__31128),
            .I(N__31124));
    InMux I__7514 (
            .O(N__31127),
            .I(N__31121));
    Odrv12 I__7513 (
            .O(N__31124),
            .I(M_this_oam_ram_read_data_1));
    LocalMux I__7512 (
            .O(N__31121),
            .I(M_this_oam_ram_read_data_1));
    InMux I__7511 (
            .O(N__31116),
            .I(N__31113));
    LocalMux I__7510 (
            .O(N__31113),
            .I(N__31110));
    Span4Mux_v I__7509 (
            .O(N__31110),
            .I(N__31106));
    CascadeMux I__7508 (
            .O(N__31109),
            .I(N__31103));
    Span4Mux_h I__7507 (
            .O(N__31106),
            .I(N__31100));
    InMux I__7506 (
            .O(N__31103),
            .I(N__31097));
    Span4Mux_h I__7505 (
            .O(N__31100),
            .I(N__31094));
    LocalMux I__7504 (
            .O(N__31097),
            .I(M_this_oam_ram_read_data_0));
    Odrv4 I__7503 (
            .O(N__31094),
            .I(M_this_oam_ram_read_data_0));
    InMux I__7502 (
            .O(N__31089),
            .I(N__31086));
    LocalMux I__7501 (
            .O(N__31086),
            .I(N__31083));
    Span12Mux_v I__7500 (
            .O(N__31083),
            .I(N__31080));
    Span12Mux_h I__7499 (
            .O(N__31080),
            .I(N__31076));
    InMux I__7498 (
            .O(N__31079),
            .I(N__31073));
    Odrv12 I__7497 (
            .O(N__31076),
            .I(M_this_oam_ram_read_data_3));
    LocalMux I__7496 (
            .O(N__31073),
            .I(M_this_oam_ram_read_data_3));
    InMux I__7495 (
            .O(N__31068),
            .I(N__31065));
    LocalMux I__7494 (
            .O(N__31065),
            .I(N__31062));
    Span4Mux_v I__7493 (
            .O(N__31062),
            .I(N__31059));
    Odrv4 I__7492 (
            .O(N__31059),
            .I(\this_ppu.un9lto7Z0Z_5 ));
    CascadeMux I__7491 (
            .O(N__31056),
            .I(N__31053));
    InMux I__7490 (
            .O(N__31053),
            .I(N__31050));
    LocalMux I__7489 (
            .O(N__31050),
            .I(N__31047));
    Span4Mux_h I__7488 (
            .O(N__31047),
            .I(N__31044));
    Odrv4 I__7487 (
            .O(N__31044),
            .I(\this_ppu.un1_M_haddress_q_2_6 ));
    CascadeMux I__7486 (
            .O(N__31041),
            .I(N__31038));
    InMux I__7485 (
            .O(N__31038),
            .I(N__31035));
    LocalMux I__7484 (
            .O(N__31035),
            .I(N__31032));
    Span4Mux_h I__7483 (
            .O(N__31032),
            .I(N__31028));
    InMux I__7482 (
            .O(N__31031),
            .I(N__31025));
    Odrv4 I__7481 (
            .O(N__31028),
            .I(M_this_oam_ram_read_data_4));
    LocalMux I__7480 (
            .O(N__31025),
            .I(M_this_oam_ram_read_data_4));
    InMux I__7479 (
            .O(N__31020),
            .I(N__31017));
    LocalMux I__7478 (
            .O(N__31017),
            .I(N__31014));
    Span4Mux_h I__7477 (
            .O(N__31014),
            .I(N__31010));
    InMux I__7476 (
            .O(N__31013),
            .I(N__31007));
    Odrv4 I__7475 (
            .O(N__31010),
            .I(M_this_oam_ram_read_data_6));
    LocalMux I__7474 (
            .O(N__31007),
            .I(M_this_oam_ram_read_data_6));
    InMux I__7473 (
            .O(N__31002),
            .I(N__30999));
    LocalMux I__7472 (
            .O(N__30999),
            .I(N__30996));
    Span4Mux_v I__7471 (
            .O(N__30996),
            .I(N__30992));
    CascadeMux I__7470 (
            .O(N__30995),
            .I(N__30989));
    Span4Mux_h I__7469 (
            .O(N__30992),
            .I(N__30986));
    InMux I__7468 (
            .O(N__30989),
            .I(N__30983));
    Odrv4 I__7467 (
            .O(N__30986),
            .I(M_this_oam_ram_read_data_7));
    LocalMux I__7466 (
            .O(N__30983),
            .I(M_this_oam_ram_read_data_7));
    InMux I__7465 (
            .O(N__30978),
            .I(N__30975));
    LocalMux I__7464 (
            .O(N__30975),
            .I(N__30972));
    Span4Mux_h I__7463 (
            .O(N__30972),
            .I(N__30969));
    Span4Mux_h I__7462 (
            .O(N__30969),
            .I(N__30965));
    InMux I__7461 (
            .O(N__30968),
            .I(N__30962));
    Odrv4 I__7460 (
            .O(N__30965),
            .I(M_this_oam_ram_read_data_5));
    LocalMux I__7459 (
            .O(N__30962),
            .I(M_this_oam_ram_read_data_5));
    InMux I__7458 (
            .O(N__30957),
            .I(N__30954));
    LocalMux I__7457 (
            .O(N__30954),
            .I(N__30951));
    Span4Mux_h I__7456 (
            .O(N__30951),
            .I(N__30948));
    Odrv4 I__7455 (
            .O(N__30948),
            .I(\this_ppu.un9lto7Z0Z_4 ));
    CascadeMux I__7454 (
            .O(N__30945),
            .I(N__30942));
    InMux I__7453 (
            .O(N__30942),
            .I(N__30939));
    LocalMux I__7452 (
            .O(N__30939),
            .I(N__30936));
    Span4Mux_v I__7451 (
            .O(N__30936),
            .I(N__30933));
    Odrv4 I__7450 (
            .O(N__30933),
            .I(\this_ppu.un1_M_vaddress_q_3_4 ));
    InMux I__7449 (
            .O(N__30930),
            .I(N__30924));
    InMux I__7448 (
            .O(N__30929),
            .I(N__30921));
    InMux I__7447 (
            .O(N__30928),
            .I(N__30916));
    InMux I__7446 (
            .O(N__30927),
            .I(N__30916));
    LocalMux I__7445 (
            .O(N__30924),
            .I(N__30912));
    LocalMux I__7444 (
            .O(N__30921),
            .I(N__30909));
    LocalMux I__7443 (
            .O(N__30916),
            .I(N__30906));
    InMux I__7442 (
            .O(N__30915),
            .I(N__30902));
    Span4Mux_v I__7441 (
            .O(N__30912),
            .I(N__30899));
    Span4Mux_h I__7440 (
            .O(N__30909),
            .I(N__30896));
    Span4Mux_h I__7439 (
            .O(N__30906),
            .I(N__30893));
    InMux I__7438 (
            .O(N__30905),
            .I(N__30890));
    LocalMux I__7437 (
            .O(N__30902),
            .I(M_this_oam_ram_read_data_11));
    Odrv4 I__7436 (
            .O(N__30899),
            .I(M_this_oam_ram_read_data_11));
    Odrv4 I__7435 (
            .O(N__30896),
            .I(M_this_oam_ram_read_data_11));
    Odrv4 I__7434 (
            .O(N__30893),
            .I(M_this_oam_ram_read_data_11));
    LocalMux I__7433 (
            .O(N__30890),
            .I(M_this_oam_ram_read_data_11));
    InMux I__7432 (
            .O(N__30879),
            .I(N__30875));
    InMux I__7431 (
            .O(N__30878),
            .I(N__30872));
    LocalMux I__7430 (
            .O(N__30875),
            .I(N__30865));
    LocalMux I__7429 (
            .O(N__30872),
            .I(N__30865));
    InMux I__7428 (
            .O(N__30871),
            .I(N__30862));
    InMux I__7427 (
            .O(N__30870),
            .I(N__30858));
    Span4Mux_v I__7426 (
            .O(N__30865),
            .I(N__30855));
    LocalMux I__7425 (
            .O(N__30862),
            .I(N__30852));
    InMux I__7424 (
            .O(N__30861),
            .I(N__30849));
    LocalMux I__7423 (
            .O(N__30858),
            .I(M_this_oam_ram_read_data_12));
    Odrv4 I__7422 (
            .O(N__30855),
            .I(M_this_oam_ram_read_data_12));
    Odrv12 I__7421 (
            .O(N__30852),
            .I(M_this_oam_ram_read_data_12));
    LocalMux I__7420 (
            .O(N__30849),
            .I(M_this_oam_ram_read_data_12));
    CascadeMux I__7419 (
            .O(N__30840),
            .I(N__30837));
    InMux I__7418 (
            .O(N__30837),
            .I(N__30834));
    LocalMux I__7417 (
            .O(N__30834),
            .I(N__30831));
    Span4Mux_h I__7416 (
            .O(N__30831),
            .I(N__30827));
    InMux I__7415 (
            .O(N__30830),
            .I(N__30824));
    Odrv4 I__7414 (
            .O(N__30827),
            .I(M_this_oam_ram_read_data_15));
    LocalMux I__7413 (
            .O(N__30824),
            .I(M_this_oam_ram_read_data_15));
    CascadeMux I__7412 (
            .O(N__30819),
            .I(N__30816));
    InMux I__7411 (
            .O(N__30816),
            .I(N__30812));
    CascadeMux I__7410 (
            .O(N__30815),
            .I(N__30808));
    LocalMux I__7409 (
            .O(N__30812),
            .I(N__30805));
    InMux I__7408 (
            .O(N__30811),
            .I(N__30802));
    InMux I__7407 (
            .O(N__30808),
            .I(N__30799));
    Span4Mux_h I__7406 (
            .O(N__30805),
            .I(N__30796));
    LocalMux I__7405 (
            .O(N__30802),
            .I(M_this_oam_ram_read_data_14));
    LocalMux I__7404 (
            .O(N__30799),
            .I(M_this_oam_ram_read_data_14));
    Odrv4 I__7403 (
            .O(N__30796),
            .I(M_this_oam_ram_read_data_14));
    CascadeMux I__7402 (
            .O(N__30789),
            .I(\this_ppu.un1_oam_data_1_c2_cascade_ ));
    CascadeMux I__7401 (
            .O(N__30786),
            .I(N__30783));
    InMux I__7400 (
            .O(N__30783),
            .I(N__30779));
    InMux I__7399 (
            .O(N__30782),
            .I(N__30776));
    LocalMux I__7398 (
            .O(N__30779),
            .I(N__30771));
    LocalMux I__7397 (
            .O(N__30776),
            .I(N__30768));
    InMux I__7396 (
            .O(N__30775),
            .I(N__30765));
    InMux I__7395 (
            .O(N__30774),
            .I(N__30762));
    Span4Mux_v I__7394 (
            .O(N__30771),
            .I(N__30759));
    Span4Mux_h I__7393 (
            .O(N__30768),
            .I(N__30756));
    LocalMux I__7392 (
            .O(N__30765),
            .I(M_this_oam_ram_read_data_13));
    LocalMux I__7391 (
            .O(N__30762),
            .I(M_this_oam_ram_read_data_13));
    Odrv4 I__7390 (
            .O(N__30759),
            .I(M_this_oam_ram_read_data_13));
    Odrv4 I__7389 (
            .O(N__30756),
            .I(M_this_oam_ram_read_data_13));
    InMux I__7388 (
            .O(N__30747),
            .I(N__30744));
    LocalMux I__7387 (
            .O(N__30744),
            .I(N__30741));
    Odrv4 I__7386 (
            .O(N__30741),
            .I(\this_ppu.un1_M_haddress_q_2_7 ));
    CascadeMux I__7385 (
            .O(N__30738),
            .I(N__30735));
    InMux I__7384 (
            .O(N__30735),
            .I(N__30732));
    LocalMux I__7383 (
            .O(N__30732),
            .I(N__30729));
    Span4Mux_v I__7382 (
            .O(N__30729),
            .I(N__30726));
    Odrv4 I__7381 (
            .O(N__30726),
            .I(M_this_data_tmp_qZ0Z_6));
    InMux I__7380 (
            .O(N__30723),
            .I(N__30720));
    LocalMux I__7379 (
            .O(N__30720),
            .I(N_67_0));
    CascadeMux I__7378 (
            .O(N__30717),
            .I(N__30714));
    CascadeBuf I__7377 (
            .O(N__30714),
            .I(N__30711));
    CascadeMux I__7376 (
            .O(N__30711),
            .I(N__30707));
    CascadeMux I__7375 (
            .O(N__30710),
            .I(N__30704));
    InMux I__7374 (
            .O(N__30707),
            .I(N__30701));
    InMux I__7373 (
            .O(N__30704),
            .I(N__30698));
    LocalMux I__7372 (
            .O(N__30701),
            .I(N__30695));
    LocalMux I__7371 (
            .O(N__30698),
            .I(M_this_oam_address_qZ0Z_5));
    Odrv12 I__7370 (
            .O(N__30695),
            .I(M_this_oam_address_qZ0Z_5));
    InMux I__7369 (
            .O(N__30690),
            .I(N__30686));
    InMux I__7368 (
            .O(N__30689),
            .I(N__30679));
    LocalMux I__7367 (
            .O(N__30686),
            .I(N__30676));
    InMux I__7366 (
            .O(N__30685),
            .I(N__30671));
    InMux I__7365 (
            .O(N__30684),
            .I(N__30671));
    InMux I__7364 (
            .O(N__30683),
            .I(N__30668));
    InMux I__7363 (
            .O(N__30682),
            .I(N__30665));
    LocalMux I__7362 (
            .O(N__30679),
            .I(N__30662));
    Span4Mux_v I__7361 (
            .O(N__30676),
            .I(N__30655));
    LocalMux I__7360 (
            .O(N__30671),
            .I(N__30655));
    LocalMux I__7359 (
            .O(N__30668),
            .I(N__30655));
    LocalMux I__7358 (
            .O(N__30665),
            .I(N__30652));
    Span12Mux_v I__7357 (
            .O(N__30662),
            .I(N__30649));
    Span4Mux_h I__7356 (
            .O(N__30655),
            .I(N__30646));
    Odrv12 I__7355 (
            .O(N__30652),
            .I(N_1152_0));
    Odrv12 I__7354 (
            .O(N__30649),
            .I(N_1152_0));
    Odrv4 I__7353 (
            .O(N__30646),
            .I(N_1152_0));
    CascadeMux I__7352 (
            .O(N__30639),
            .I(N__30636));
    CascadeBuf I__7351 (
            .O(N__30636),
            .I(N__30631));
    CascadeMux I__7350 (
            .O(N__30635),
            .I(N__30628));
    InMux I__7349 (
            .O(N__30634),
            .I(N__30625));
    CascadeMux I__7348 (
            .O(N__30631),
            .I(N__30622));
    InMux I__7347 (
            .O(N__30628),
            .I(N__30618));
    LocalMux I__7346 (
            .O(N__30625),
            .I(N__30615));
    InMux I__7345 (
            .O(N__30622),
            .I(N__30612));
    InMux I__7344 (
            .O(N__30621),
            .I(N__30609));
    LocalMux I__7343 (
            .O(N__30618),
            .I(N__30602));
    Span12Mux_v I__7342 (
            .O(N__30615),
            .I(N__30602));
    LocalMux I__7341 (
            .O(N__30612),
            .I(N__30602));
    LocalMux I__7340 (
            .O(N__30609),
            .I(M_this_oam_address_qZ0Z_3));
    Odrv12 I__7339 (
            .O(N__30602),
            .I(M_this_oam_address_qZ0Z_3));
    CascadeMux I__7338 (
            .O(N__30597),
            .I(N__30594));
    CascadeBuf I__7337 (
            .O(N__30594),
            .I(N__30591));
    CascadeMux I__7336 (
            .O(N__30591),
            .I(N__30587));
    InMux I__7335 (
            .O(N__30590),
            .I(N__30582));
    InMux I__7334 (
            .O(N__30587),
            .I(N__30578));
    InMux I__7333 (
            .O(N__30586),
            .I(N__30575));
    InMux I__7332 (
            .O(N__30585),
            .I(N__30572));
    LocalMux I__7331 (
            .O(N__30582),
            .I(N__30569));
    InMux I__7330 (
            .O(N__30581),
            .I(N__30566));
    LocalMux I__7329 (
            .O(N__30578),
            .I(N__30563));
    LocalMux I__7328 (
            .O(N__30575),
            .I(M_this_oam_address_qZ0Z_2));
    LocalMux I__7327 (
            .O(N__30572),
            .I(M_this_oam_address_qZ0Z_2));
    Odrv12 I__7326 (
            .O(N__30569),
            .I(M_this_oam_address_qZ0Z_2));
    LocalMux I__7325 (
            .O(N__30566),
            .I(M_this_oam_address_qZ0Z_2));
    Odrv12 I__7324 (
            .O(N__30563),
            .I(M_this_oam_address_qZ0Z_2));
    InMux I__7323 (
            .O(N__30552),
            .I(N__30547));
    InMux I__7322 (
            .O(N__30551),
            .I(N__30542));
    InMux I__7321 (
            .O(N__30550),
            .I(N__30542));
    LocalMux I__7320 (
            .O(N__30547),
            .I(un1_M_this_oam_address_q_c2));
    LocalMux I__7319 (
            .O(N__30542),
            .I(un1_M_this_oam_address_q_c2));
    InMux I__7318 (
            .O(N__30537),
            .I(N__30534));
    LocalMux I__7317 (
            .O(N__30534),
            .I(un1_M_this_oam_address_q_c4));
    InMux I__7316 (
            .O(N__30531),
            .I(N__30528));
    LocalMux I__7315 (
            .O(N__30528),
            .I(N__30525));
    Odrv12 I__7314 (
            .O(N__30525),
            .I(N_50_0));
    InMux I__7313 (
            .O(N__30522),
            .I(N__30519));
    LocalMux I__7312 (
            .O(N__30519),
            .I(N__30516));
    Span4Mux_v I__7311 (
            .O(N__30516),
            .I(N__30513));
    Odrv4 I__7310 (
            .O(N__30513),
            .I(N_46_0));
    CascadeMux I__7309 (
            .O(N__30510),
            .I(N__30507));
    InMux I__7308 (
            .O(N__30507),
            .I(N__30504));
    LocalMux I__7307 (
            .O(N__30504),
            .I(M_this_data_tmp_qZ0Z_21));
    CascadeMux I__7306 (
            .O(N__30501),
            .I(N__30498));
    InMux I__7305 (
            .O(N__30498),
            .I(N__30495));
    LocalMux I__7304 (
            .O(N__30495),
            .I(N__30492));
    Odrv4 I__7303 (
            .O(N__30492),
            .I(M_this_data_tmp_qZ0Z_10));
    InMux I__7302 (
            .O(N__30489),
            .I(N__30486));
    LocalMux I__7301 (
            .O(N__30486),
            .I(N__30483));
    Span4Mux_v I__7300 (
            .O(N__30483),
            .I(N__30480));
    Odrv4 I__7299 (
            .O(N__30480),
            .I(\this_sprites_ram.mem_out_bus5_3 ));
    InMux I__7298 (
            .O(N__30477),
            .I(N__30474));
    LocalMux I__7297 (
            .O(N__30474),
            .I(N__30471));
    Span4Mux_v I__7296 (
            .O(N__30471),
            .I(N__30468));
    Odrv4 I__7295 (
            .O(N__30468),
            .I(\this_sprites_ram.mem_out_bus1_3 ));
    InMux I__7294 (
            .O(N__30465),
            .I(N__30461));
    InMux I__7293 (
            .O(N__30464),
            .I(N__30450));
    LocalMux I__7292 (
            .O(N__30461),
            .I(N__30446));
    InMux I__7291 (
            .O(N__30460),
            .I(N__30443));
    InMux I__7290 (
            .O(N__30459),
            .I(N__30440));
    InMux I__7289 (
            .O(N__30458),
            .I(N__30431));
    InMux I__7288 (
            .O(N__30457),
            .I(N__30431));
    InMux I__7287 (
            .O(N__30456),
            .I(N__30431));
    InMux I__7286 (
            .O(N__30455),
            .I(N__30431));
    InMux I__7285 (
            .O(N__30454),
            .I(N__30426));
    InMux I__7284 (
            .O(N__30453),
            .I(N__30426));
    LocalMux I__7283 (
            .O(N__30450),
            .I(N__30420));
    InMux I__7282 (
            .O(N__30449),
            .I(N__30415));
    Span4Mux_h I__7281 (
            .O(N__30446),
            .I(N__30404));
    LocalMux I__7280 (
            .O(N__30443),
            .I(N__30404));
    LocalMux I__7279 (
            .O(N__30440),
            .I(N__30404));
    LocalMux I__7278 (
            .O(N__30431),
            .I(N__30404));
    LocalMux I__7277 (
            .O(N__30426),
            .I(N__30404));
    InMux I__7276 (
            .O(N__30425),
            .I(N__30397));
    InMux I__7275 (
            .O(N__30424),
            .I(N__30397));
    InMux I__7274 (
            .O(N__30423),
            .I(N__30397));
    Span4Mux_h I__7273 (
            .O(N__30420),
            .I(N__30394));
    InMux I__7272 (
            .O(N__30419),
            .I(N__30389));
    InMux I__7271 (
            .O(N__30418),
            .I(N__30389));
    LocalMux I__7270 (
            .O(N__30415),
            .I(N__30386));
    Span4Mux_h I__7269 (
            .O(N__30404),
            .I(N__30383));
    LocalMux I__7268 (
            .O(N__30397),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__7267 (
            .O(N__30394),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    LocalMux I__7266 (
            .O(N__30389),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__7265 (
            .O(N__30386),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__7264 (
            .O(N__30383),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    InMux I__7263 (
            .O(N__30372),
            .I(N__30369));
    LocalMux I__7262 (
            .O(N__30369),
            .I(N__30366));
    Span4Mux_h I__7261 (
            .O(N__30366),
            .I(N__30363));
    Span4Mux_h I__7260 (
            .O(N__30363),
            .I(N__30360));
    Odrv4 I__7259 (
            .O(N__30360),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ));
    CEMux I__7258 (
            .O(N__30357),
            .I(N__30353));
    CEMux I__7257 (
            .O(N__30356),
            .I(N__30350));
    LocalMux I__7256 (
            .O(N__30353),
            .I(N__30347));
    LocalMux I__7255 (
            .O(N__30350),
            .I(N__30344));
    Span4Mux_v I__7254 (
            .O(N__30347),
            .I(N__30339));
    Span4Mux_h I__7253 (
            .O(N__30344),
            .I(N__30339));
    Odrv4 I__7252 (
            .O(N__30339),
            .I(\this_sprites_ram.mem_WE_10 ));
    CascadeMux I__7251 (
            .O(N__30336),
            .I(N__30333));
    InMux I__7250 (
            .O(N__30333),
            .I(N__30329));
    InMux I__7249 (
            .O(N__30332),
            .I(N__30326));
    LocalMux I__7248 (
            .O(N__30329),
            .I(N__30323));
    LocalMux I__7247 (
            .O(N__30326),
            .I(\this_ppu.M_this_ppu_map_addr_i_5 ));
    Odrv4 I__7246 (
            .O(N__30323),
            .I(\this_ppu.M_this_ppu_map_addr_i_5 ));
    CascadeMux I__7245 (
            .O(N__30318),
            .I(N__30315));
    InMux I__7244 (
            .O(N__30315),
            .I(N__30311));
    InMux I__7243 (
            .O(N__30314),
            .I(N__30308));
    LocalMux I__7242 (
            .O(N__30311),
            .I(N__30305));
    LocalMux I__7241 (
            .O(N__30308),
            .I(\this_ppu.M_this_ppu_map_addr_i_6 ));
    Odrv4 I__7240 (
            .O(N__30305),
            .I(\this_ppu.M_this_ppu_map_addr_i_6 ));
    CascadeMux I__7239 (
            .O(N__30300),
            .I(N__30297));
    InMux I__7238 (
            .O(N__30297),
            .I(N__30293));
    InMux I__7237 (
            .O(N__30296),
            .I(N__30290));
    LocalMux I__7236 (
            .O(N__30293),
            .I(N__30287));
    LocalMux I__7235 (
            .O(N__30290),
            .I(\this_ppu.M_this_ppu_map_addr_i_7 ));
    Odrv4 I__7234 (
            .O(N__30287),
            .I(\this_ppu.M_this_ppu_map_addr_i_7 ));
    CascadeMux I__7233 (
            .O(N__30282),
            .I(N__30279));
    InMux I__7232 (
            .O(N__30279),
            .I(N__30275));
    InMux I__7231 (
            .O(N__30278),
            .I(N__30272));
    LocalMux I__7230 (
            .O(N__30275),
            .I(N__30269));
    LocalMux I__7229 (
            .O(N__30272),
            .I(\this_ppu.M_this_ppu_map_addr_i_8 ));
    Odrv4 I__7228 (
            .O(N__30269),
            .I(\this_ppu.M_this_ppu_map_addr_i_8 ));
    CascadeMux I__7227 (
            .O(N__30264),
            .I(N__30260));
    InMux I__7226 (
            .O(N__30263),
            .I(N__30257));
    InMux I__7225 (
            .O(N__30260),
            .I(N__30254));
    LocalMux I__7224 (
            .O(N__30257),
            .I(N__30251));
    LocalMux I__7223 (
            .O(N__30254),
            .I(\this_ppu.M_this_ppu_map_addr_i_9 ));
    Odrv4 I__7222 (
            .O(N__30251),
            .I(\this_ppu.M_this_ppu_map_addr_i_9 ));
    InMux I__7221 (
            .O(N__30246),
            .I(bfn_23_20_0_));
    CascadeMux I__7220 (
            .O(N__30243),
            .I(N__30240));
    InMux I__7219 (
            .O(N__30240),
            .I(N__30237));
    LocalMux I__7218 (
            .O(N__30237),
            .I(\this_ppu.un1_M_vaddress_q_cry_7_THRU_CO ));
    InMux I__7217 (
            .O(N__30234),
            .I(N__30231));
    LocalMux I__7216 (
            .O(N__30231),
            .I(N__30228));
    Span12Mux_s9_h I__7215 (
            .O(N__30228),
            .I(N__30225));
    Odrv12 I__7214 (
            .O(N__30225),
            .I(N_61_0));
    InMux I__7213 (
            .O(N__30222),
            .I(N__30219));
    LocalMux I__7212 (
            .O(N__30219),
            .I(N__30216));
    Span4Mux_v I__7211 (
            .O(N__30216),
            .I(N__30213));
    Odrv4 I__7210 (
            .O(N__30213),
            .I(M_this_data_tmp_qZ0Z_3));
    InMux I__7209 (
            .O(N__30210),
            .I(N__30207));
    LocalMux I__7208 (
            .O(N__30207),
            .I(N__30204));
    Span4Mux_v I__7207 (
            .O(N__30204),
            .I(N__30201));
    Odrv4 I__7206 (
            .O(N__30201),
            .I(N_73_0));
    CascadeMux I__7205 (
            .O(N__30198),
            .I(N__30195));
    CascadeBuf I__7204 (
            .O(N__30195),
            .I(N__30192));
    CascadeMux I__7203 (
            .O(N__30192),
            .I(N__30188));
    InMux I__7202 (
            .O(N__30191),
            .I(N__30185));
    InMux I__7201 (
            .O(N__30188),
            .I(N__30182));
    LocalMux I__7200 (
            .O(N__30185),
            .I(N__30176));
    LocalMux I__7199 (
            .O(N__30182),
            .I(N__30176));
    InMux I__7198 (
            .O(N__30181),
            .I(N__30173));
    Span4Mux_h I__7197 (
            .O(N__30176),
            .I(N__30170));
    LocalMux I__7196 (
            .O(N__30173),
            .I(M_this_oam_address_qZ0Z_4));
    Odrv4 I__7195 (
            .O(N__30170),
            .I(M_this_oam_address_qZ0Z_4));
    CascadeMux I__7194 (
            .O(N__30165),
            .I(N__30157));
    CascadeMux I__7193 (
            .O(N__30164),
            .I(N__30154));
    CascadeMux I__7192 (
            .O(N__30163),
            .I(N__30149));
    CascadeMux I__7191 (
            .O(N__30162),
            .I(N__30146));
    InMux I__7190 (
            .O(N__30161),
            .I(N__30142));
    InMux I__7189 (
            .O(N__30160),
            .I(N__30137));
    InMux I__7188 (
            .O(N__30157),
            .I(N__30137));
    InMux I__7187 (
            .O(N__30154),
            .I(N__30133));
    CascadeMux I__7186 (
            .O(N__30153),
            .I(N__30130));
    InMux I__7185 (
            .O(N__30152),
            .I(N__30127));
    InMux I__7184 (
            .O(N__30149),
            .I(N__30124));
    InMux I__7183 (
            .O(N__30146),
            .I(N__30121));
    CascadeMux I__7182 (
            .O(N__30145),
            .I(N__30118));
    LocalMux I__7181 (
            .O(N__30142),
            .I(N__30113));
    LocalMux I__7180 (
            .O(N__30137),
            .I(N__30113));
    CascadeMux I__7179 (
            .O(N__30136),
            .I(N__30109));
    LocalMux I__7178 (
            .O(N__30133),
            .I(N__30105));
    InMux I__7177 (
            .O(N__30130),
            .I(N__30102));
    LocalMux I__7176 (
            .O(N__30127),
            .I(N__30097));
    LocalMux I__7175 (
            .O(N__30124),
            .I(N__30097));
    LocalMux I__7174 (
            .O(N__30121),
            .I(N__30094));
    InMux I__7173 (
            .O(N__30118),
            .I(N__30091));
    Span4Mux_v I__7172 (
            .O(N__30113),
            .I(N__30088));
    InMux I__7171 (
            .O(N__30112),
            .I(N__30083));
    InMux I__7170 (
            .O(N__30109),
            .I(N__30083));
    InMux I__7169 (
            .O(N__30108),
            .I(N__30078));
    Span4Mux_h I__7168 (
            .O(N__30105),
            .I(N__30075));
    LocalMux I__7167 (
            .O(N__30102),
            .I(N__30072));
    Span4Mux_v I__7166 (
            .O(N__30097),
            .I(N__30069));
    Span4Mux_h I__7165 (
            .O(N__30094),
            .I(N__30064));
    LocalMux I__7164 (
            .O(N__30091),
            .I(N__30064));
    Span4Mux_h I__7163 (
            .O(N__30088),
            .I(N__30059));
    LocalMux I__7162 (
            .O(N__30083),
            .I(N__30059));
    CascadeMux I__7161 (
            .O(N__30082),
            .I(N__30056));
    InMux I__7160 (
            .O(N__30081),
            .I(N__30052));
    LocalMux I__7159 (
            .O(N__30078),
            .I(N__30045));
    Span4Mux_h I__7158 (
            .O(N__30075),
            .I(N__30045));
    Span4Mux_h I__7157 (
            .O(N__30072),
            .I(N__30045));
    Span4Mux_h I__7156 (
            .O(N__30069),
            .I(N__30038));
    Span4Mux_h I__7155 (
            .O(N__30064),
            .I(N__30038));
    Span4Mux_h I__7154 (
            .O(N__30059),
            .I(N__30038));
    InMux I__7153 (
            .O(N__30056),
            .I(N__30033));
    InMux I__7152 (
            .O(N__30055),
            .I(N__30033));
    LocalMux I__7151 (
            .O(N__30052),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    Odrv4 I__7150 (
            .O(N__30045),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    Odrv4 I__7149 (
            .O(N__30038),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    LocalMux I__7148 (
            .O(N__30033),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    CascadeMux I__7147 (
            .O(N__30024),
            .I(\this_ppu.un2_vscroll_axb_0_cascade_ ));
    InMux I__7146 (
            .O(N__30021),
            .I(N__30013));
    InMux I__7145 (
            .O(N__30020),
            .I(N__30010));
    InMux I__7144 (
            .O(N__30019),
            .I(N__30007));
    CascadeMux I__7143 (
            .O(N__30018),
            .I(N__30003));
    InMux I__7142 (
            .O(N__30017),
            .I(N__29992));
    InMux I__7141 (
            .O(N__30016),
            .I(N__29992));
    LocalMux I__7140 (
            .O(N__30013),
            .I(N__29987));
    LocalMux I__7139 (
            .O(N__30010),
            .I(N__29982));
    LocalMux I__7138 (
            .O(N__30007),
            .I(N__29982));
    InMux I__7137 (
            .O(N__30006),
            .I(N__29979));
    InMux I__7136 (
            .O(N__30003),
            .I(N__29975));
    InMux I__7135 (
            .O(N__30002),
            .I(N__29972));
    InMux I__7134 (
            .O(N__30001),
            .I(N__29969));
    InMux I__7133 (
            .O(N__30000),
            .I(N__29966));
    InMux I__7132 (
            .O(N__29999),
            .I(N__29963));
    InMux I__7131 (
            .O(N__29998),
            .I(N__29958));
    InMux I__7130 (
            .O(N__29997),
            .I(N__29958));
    LocalMux I__7129 (
            .O(N__29992),
            .I(N__29955));
    InMux I__7128 (
            .O(N__29991),
            .I(N__29952));
    InMux I__7127 (
            .O(N__29990),
            .I(N__29949));
    Span4Mux_v I__7126 (
            .O(N__29987),
            .I(N__29942));
    Span4Mux_h I__7125 (
            .O(N__29982),
            .I(N__29942));
    LocalMux I__7124 (
            .O(N__29979),
            .I(N__29942));
    InMux I__7123 (
            .O(N__29978),
            .I(N__29938));
    LocalMux I__7122 (
            .O(N__29975),
            .I(N__29931));
    LocalMux I__7121 (
            .O(N__29972),
            .I(N__29931));
    LocalMux I__7120 (
            .O(N__29969),
            .I(N__29931));
    LocalMux I__7119 (
            .O(N__29966),
            .I(N__29928));
    LocalMux I__7118 (
            .O(N__29963),
            .I(N__29919));
    LocalMux I__7117 (
            .O(N__29958),
            .I(N__29919));
    Span4Mux_v I__7116 (
            .O(N__29955),
            .I(N__29919));
    LocalMux I__7115 (
            .O(N__29952),
            .I(N__29919));
    LocalMux I__7114 (
            .O(N__29949),
            .I(N__29916));
    Span4Mux_h I__7113 (
            .O(N__29942),
            .I(N__29913));
    InMux I__7112 (
            .O(N__29941),
            .I(N__29910));
    LocalMux I__7111 (
            .O(N__29938),
            .I(N__29907));
    Span12Mux_h I__7110 (
            .O(N__29931),
            .I(N__29904));
    Span4Mux_v I__7109 (
            .O(N__29928),
            .I(N__29899));
    Span4Mux_h I__7108 (
            .O(N__29919),
            .I(N__29899));
    Span4Mux_h I__7107 (
            .O(N__29916),
            .I(N__29896));
    Odrv4 I__7106 (
            .O(N__29913),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    LocalMux I__7105 (
            .O(N__29910),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv4 I__7104 (
            .O(N__29907),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv12 I__7103 (
            .O(N__29904),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv4 I__7102 (
            .O(N__29899),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv4 I__7101 (
            .O(N__29896),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    CascadeMux I__7100 (
            .O(N__29883),
            .I(N__29879));
    CascadeMux I__7099 (
            .O(N__29882),
            .I(N__29876));
    InMux I__7098 (
            .O(N__29879),
            .I(N__29871));
    InMux I__7097 (
            .O(N__29876),
            .I(N__29866));
    CascadeMux I__7096 (
            .O(N__29875),
            .I(N__29863));
    CascadeMux I__7095 (
            .O(N__29874),
            .I(N__29859));
    LocalMux I__7094 (
            .O(N__29871),
            .I(N__29855));
    CascadeMux I__7093 (
            .O(N__29870),
            .I(N__29852));
    CascadeMux I__7092 (
            .O(N__29869),
            .I(N__29848));
    LocalMux I__7091 (
            .O(N__29866),
            .I(N__29844));
    InMux I__7090 (
            .O(N__29863),
            .I(N__29841));
    CascadeMux I__7089 (
            .O(N__29862),
            .I(N__29838));
    InMux I__7088 (
            .O(N__29859),
            .I(N__29835));
    CascadeMux I__7087 (
            .O(N__29858),
            .I(N__29832));
    Span4Mux_h I__7086 (
            .O(N__29855),
            .I(N__29829));
    InMux I__7085 (
            .O(N__29852),
            .I(N__29826));
    CascadeMux I__7084 (
            .O(N__29851),
            .I(N__29823));
    InMux I__7083 (
            .O(N__29848),
            .I(N__29819));
    CascadeMux I__7082 (
            .O(N__29847),
            .I(N__29816));
    Span4Mux_v I__7081 (
            .O(N__29844),
            .I(N__29809));
    LocalMux I__7080 (
            .O(N__29841),
            .I(N__29809));
    InMux I__7079 (
            .O(N__29838),
            .I(N__29805));
    LocalMux I__7078 (
            .O(N__29835),
            .I(N__29802));
    InMux I__7077 (
            .O(N__29832),
            .I(N__29799));
    Span4Mux_v I__7076 (
            .O(N__29829),
            .I(N__29793));
    LocalMux I__7075 (
            .O(N__29826),
            .I(N__29793));
    InMux I__7074 (
            .O(N__29823),
            .I(N__29790));
    CascadeMux I__7073 (
            .O(N__29822),
            .I(N__29787));
    LocalMux I__7072 (
            .O(N__29819),
            .I(N__29784));
    InMux I__7071 (
            .O(N__29816),
            .I(N__29781));
    CascadeMux I__7070 (
            .O(N__29815),
            .I(N__29778));
    CascadeMux I__7069 (
            .O(N__29814),
            .I(N__29774));
    Span4Mux_h I__7068 (
            .O(N__29809),
            .I(N__29771));
    CascadeMux I__7067 (
            .O(N__29808),
            .I(N__29768));
    LocalMux I__7066 (
            .O(N__29805),
            .I(N__29765));
    Span4Mux_h I__7065 (
            .O(N__29802),
            .I(N__29762));
    LocalMux I__7064 (
            .O(N__29799),
            .I(N__29759));
    CascadeMux I__7063 (
            .O(N__29798),
            .I(N__29756));
    Span4Mux_h I__7062 (
            .O(N__29793),
            .I(N__29753));
    LocalMux I__7061 (
            .O(N__29790),
            .I(N__29750));
    InMux I__7060 (
            .O(N__29787),
            .I(N__29747));
    Span4Mux_h I__7059 (
            .O(N__29784),
            .I(N__29744));
    LocalMux I__7058 (
            .O(N__29781),
            .I(N__29741));
    InMux I__7057 (
            .O(N__29778),
            .I(N__29738));
    CascadeMux I__7056 (
            .O(N__29777),
            .I(N__29735));
    InMux I__7055 (
            .O(N__29774),
            .I(N__29732));
    Sp12to4 I__7054 (
            .O(N__29771),
            .I(N__29729));
    InMux I__7053 (
            .O(N__29768),
            .I(N__29726));
    Span4Mux_h I__7052 (
            .O(N__29765),
            .I(N__29723));
    Span4Mux_v I__7051 (
            .O(N__29762),
            .I(N__29718));
    Span4Mux_h I__7050 (
            .O(N__29759),
            .I(N__29718));
    InMux I__7049 (
            .O(N__29756),
            .I(N__29715));
    Span4Mux_h I__7048 (
            .O(N__29753),
            .I(N__29712));
    Span4Mux_h I__7047 (
            .O(N__29750),
            .I(N__29709));
    LocalMux I__7046 (
            .O(N__29747),
            .I(N__29706));
    Span4Mux_v I__7045 (
            .O(N__29744),
            .I(N__29701));
    Span4Mux_h I__7044 (
            .O(N__29741),
            .I(N__29701));
    LocalMux I__7043 (
            .O(N__29738),
            .I(N__29698));
    InMux I__7042 (
            .O(N__29735),
            .I(N__29695));
    LocalMux I__7041 (
            .O(N__29732),
            .I(N__29692));
    Span12Mux_h I__7040 (
            .O(N__29729),
            .I(N__29687));
    LocalMux I__7039 (
            .O(N__29726),
            .I(N__29687));
    Span4Mux_v I__7038 (
            .O(N__29723),
            .I(N__29684));
    Span4Mux_v I__7037 (
            .O(N__29718),
            .I(N__29681));
    LocalMux I__7036 (
            .O(N__29715),
            .I(N__29678));
    Span4Mux_h I__7035 (
            .O(N__29712),
            .I(N__29675));
    Span4Mux_v I__7034 (
            .O(N__29709),
            .I(N__29670));
    Span4Mux_h I__7033 (
            .O(N__29706),
            .I(N__29670));
    Span4Mux_v I__7032 (
            .O(N__29701),
            .I(N__29665));
    Span4Mux_h I__7031 (
            .O(N__29698),
            .I(N__29665));
    LocalMux I__7030 (
            .O(N__29695),
            .I(N__29662));
    Span12Mux_s9_h I__7029 (
            .O(N__29692),
            .I(N__29657));
    Span12Mux_s9_h I__7028 (
            .O(N__29687),
            .I(N__29657));
    Span4Mux_v I__7027 (
            .O(N__29684),
            .I(N__29650));
    Span4Mux_v I__7026 (
            .O(N__29681),
            .I(N__29650));
    Span4Mux_h I__7025 (
            .O(N__29678),
            .I(N__29650));
    Span4Mux_h I__7024 (
            .O(N__29675),
            .I(N__29641));
    Span4Mux_v I__7023 (
            .O(N__29670),
            .I(N__29641));
    Span4Mux_v I__7022 (
            .O(N__29665),
            .I(N__29641));
    Span4Mux_h I__7021 (
            .O(N__29662),
            .I(N__29641));
    Odrv12 I__7020 (
            .O(N__29657),
            .I(M_this_ppu_sprites_addr_3));
    Odrv4 I__7019 (
            .O(N__29650),
            .I(M_this_ppu_sprites_addr_3));
    Odrv4 I__7018 (
            .O(N__29641),
            .I(M_this_ppu_sprites_addr_3));
    InMux I__7017 (
            .O(N__29634),
            .I(N__29619));
    InMux I__7016 (
            .O(N__29633),
            .I(N__29619));
    InMux I__7015 (
            .O(N__29632),
            .I(N__29619));
    InMux I__7014 (
            .O(N__29631),
            .I(N__29619));
    InMux I__7013 (
            .O(N__29630),
            .I(N__29616));
    InMux I__7012 (
            .O(N__29629),
            .I(N__29613));
    InMux I__7011 (
            .O(N__29628),
            .I(N__29610));
    LocalMux I__7010 (
            .O(N__29619),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    LocalMux I__7009 (
            .O(N__29616),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    LocalMux I__7008 (
            .O(N__29613),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    LocalMux I__7007 (
            .O(N__29610),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    InMux I__7006 (
            .O(N__29601),
            .I(N__29595));
    InMux I__7005 (
            .O(N__29600),
            .I(N__29595));
    LocalMux I__7004 (
            .O(N__29595),
            .I(N__29591));
    CascadeMux I__7003 (
            .O(N__29594),
            .I(N__29588));
    Span4Mux_h I__7002 (
            .O(N__29591),
            .I(N__29585));
    InMux I__7001 (
            .O(N__29588),
            .I(N__29582));
    Odrv4 I__7000 (
            .O(N__29585),
            .I(\this_ppu.un1_M_vaddress_q_2_c2 ));
    LocalMux I__6999 (
            .O(N__29582),
            .I(\this_ppu.un1_M_vaddress_q_2_c2 ));
    CascadeMux I__6998 (
            .O(N__29577),
            .I(N__29574));
    CascadeBuf I__6997 (
            .O(N__29574),
            .I(N__29571));
    CascadeMux I__6996 (
            .O(N__29571),
            .I(N__29568));
    InMux I__6995 (
            .O(N__29568),
            .I(N__29565));
    LocalMux I__6994 (
            .O(N__29565),
            .I(N__29561));
    CascadeMux I__6993 (
            .O(N__29564),
            .I(N__29558));
    Span12Mux_s10_h I__6992 (
            .O(N__29561),
            .I(N__29552));
    InMux I__6991 (
            .O(N__29558),
            .I(N__29547));
    InMux I__6990 (
            .O(N__29557),
            .I(N__29547));
    InMux I__6989 (
            .O(N__29556),
            .I(N__29544));
    InMux I__6988 (
            .O(N__29555),
            .I(N__29541));
    Span12Mux_h I__6987 (
            .O(N__29552),
            .I(N__29538));
    LocalMux I__6986 (
            .O(N__29547),
            .I(M_this_ppu_map_addr_5));
    LocalMux I__6985 (
            .O(N__29544),
            .I(M_this_ppu_map_addr_5));
    LocalMux I__6984 (
            .O(N__29541),
            .I(M_this_ppu_map_addr_5));
    Odrv12 I__6983 (
            .O(N__29538),
            .I(M_this_ppu_map_addr_5));
    CascadeMux I__6982 (
            .O(N__29529),
            .I(N__29526));
    CascadeBuf I__6981 (
            .O(N__29526),
            .I(N__29523));
    CascadeMux I__6980 (
            .O(N__29523),
            .I(N__29520));
    InMux I__6979 (
            .O(N__29520),
            .I(N__29517));
    LocalMux I__6978 (
            .O(N__29517),
            .I(N__29514));
    Span4Mux_h I__6977 (
            .O(N__29514),
            .I(N__29511));
    Sp12to4 I__6976 (
            .O(N__29511),
            .I(N__29508));
    Span12Mux_s10_v I__6975 (
            .O(N__29508),
            .I(N__29502));
    InMux I__6974 (
            .O(N__29507),
            .I(N__29499));
    InMux I__6973 (
            .O(N__29506),
            .I(N__29496));
    InMux I__6972 (
            .O(N__29505),
            .I(N__29493));
    Span12Mux_h I__6971 (
            .O(N__29502),
            .I(N__29490));
    LocalMux I__6970 (
            .O(N__29499),
            .I(M_this_ppu_map_addr_6));
    LocalMux I__6969 (
            .O(N__29496),
            .I(M_this_ppu_map_addr_6));
    LocalMux I__6968 (
            .O(N__29493),
            .I(M_this_ppu_map_addr_6));
    Odrv12 I__6967 (
            .O(N__29490),
            .I(M_this_ppu_map_addr_6));
    InMux I__6966 (
            .O(N__29481),
            .I(N__29478));
    LocalMux I__6965 (
            .O(N__29478),
            .I(N__29475));
    Span4Mux_v I__6964 (
            .O(N__29475),
            .I(N__29468));
    InMux I__6963 (
            .O(N__29474),
            .I(N__29465));
    InMux I__6962 (
            .O(N__29473),
            .I(N__29460));
    InMux I__6961 (
            .O(N__29472),
            .I(N__29460));
    CascadeMux I__6960 (
            .O(N__29471),
            .I(N__29457));
    Span4Mux_h I__6959 (
            .O(N__29468),
            .I(N__29451));
    LocalMux I__6958 (
            .O(N__29465),
            .I(N__29451));
    LocalMux I__6957 (
            .O(N__29460),
            .I(N__29448));
    InMux I__6956 (
            .O(N__29457),
            .I(N__29443));
    InMux I__6955 (
            .O(N__29456),
            .I(N__29443));
    Odrv4 I__6954 (
            .O(N__29451),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    Odrv4 I__6953 (
            .O(N__29448),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__6952 (
            .O(N__29443),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    CascadeMux I__6951 (
            .O(N__29436),
            .I(N__29431));
    CascadeMux I__6950 (
            .O(N__29435),
            .I(N__29428));
    CascadeMux I__6949 (
            .O(N__29434),
            .I(N__29424));
    InMux I__6948 (
            .O(N__29431),
            .I(N__29421));
    InMux I__6947 (
            .O(N__29428),
            .I(N__29418));
    InMux I__6946 (
            .O(N__29427),
            .I(N__29413));
    InMux I__6945 (
            .O(N__29424),
            .I(N__29413));
    LocalMux I__6944 (
            .O(N__29421),
            .I(N__29410));
    LocalMux I__6943 (
            .O(N__29418),
            .I(N__29407));
    LocalMux I__6942 (
            .O(N__29413),
            .I(N__29404));
    Sp12to4 I__6941 (
            .O(N__29410),
            .I(N__29399));
    Span4Mux_h I__6940 (
            .O(N__29407),
            .I(N__29396));
    Span4Mux_v I__6939 (
            .O(N__29404),
            .I(N__29393));
    InMux I__6938 (
            .O(N__29403),
            .I(N__29388));
    InMux I__6937 (
            .O(N__29402),
            .I(N__29388));
    Odrv12 I__6936 (
            .O(N__29399),
            .I(\this_ppu.M_last_q ));
    Odrv4 I__6935 (
            .O(N__29396),
            .I(\this_ppu.M_last_q ));
    Odrv4 I__6934 (
            .O(N__29393),
            .I(\this_ppu.M_last_q ));
    LocalMux I__6933 (
            .O(N__29388),
            .I(\this_ppu.M_last_q ));
    InMux I__6932 (
            .O(N__29379),
            .I(N__29376));
    LocalMux I__6931 (
            .O(N__29376),
            .I(N__29373));
    Span4Mux_v I__6930 (
            .O(N__29373),
            .I(N__29367));
    InMux I__6929 (
            .O(N__29372),
            .I(N__29364));
    InMux I__6928 (
            .O(N__29371),
            .I(N__29359));
    InMux I__6927 (
            .O(N__29370),
            .I(N__29359));
    Span4Mux_h I__6926 (
            .O(N__29367),
            .I(N__29352));
    LocalMux I__6925 (
            .O(N__29364),
            .I(N__29352));
    LocalMux I__6924 (
            .O(N__29359),
            .I(N__29349));
    InMux I__6923 (
            .O(N__29358),
            .I(N__29344));
    InMux I__6922 (
            .O(N__29357),
            .I(N__29344));
    Odrv4 I__6921 (
            .O(N__29352),
            .I(M_this_vga_signals_line_clk_0));
    Odrv4 I__6920 (
            .O(N__29349),
            .I(M_this_vga_signals_line_clk_0));
    LocalMux I__6919 (
            .O(N__29344),
            .I(M_this_vga_signals_line_clk_0));
    CascadeMux I__6918 (
            .O(N__29337),
            .I(N__29334));
    InMux I__6917 (
            .O(N__29334),
            .I(N__29331));
    LocalMux I__6916 (
            .O(N__29331),
            .I(N__29328));
    Span4Mux_v I__6915 (
            .O(N__29328),
            .I(N__29323));
    InMux I__6914 (
            .O(N__29327),
            .I(N__29320));
    InMux I__6913 (
            .O(N__29326),
            .I(N__29316));
    Sp12to4 I__6912 (
            .O(N__29323),
            .I(N__29313));
    LocalMux I__6911 (
            .O(N__29320),
            .I(N__29310));
    InMux I__6910 (
            .O(N__29319),
            .I(N__29307));
    LocalMux I__6909 (
            .O(N__29316),
            .I(N__29299));
    Span12Mux_h I__6908 (
            .O(N__29313),
            .I(N__29296));
    Span4Mux_h I__6907 (
            .O(N__29310),
            .I(N__29291));
    LocalMux I__6906 (
            .O(N__29307),
            .I(N__29291));
    InMux I__6905 (
            .O(N__29306),
            .I(N__29284));
    InMux I__6904 (
            .O(N__29305),
            .I(N__29284));
    InMux I__6903 (
            .O(N__29304),
            .I(N__29284));
    InMux I__6902 (
            .O(N__29303),
            .I(N__29281));
    InMux I__6901 (
            .O(N__29302),
            .I(N__29278));
    Odrv4 I__6900 (
            .O(N__29299),
            .I(M_this_ppu_vram_addr_7));
    Odrv12 I__6899 (
            .O(N__29296),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__6898 (
            .O(N__29291),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__6897 (
            .O(N__29284),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__6896 (
            .O(N__29281),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__6895 (
            .O(N__29278),
            .I(M_this_ppu_vram_addr_7));
    SRMux I__6894 (
            .O(N__29265),
            .I(N__29261));
    SRMux I__6893 (
            .O(N__29264),
            .I(N__29258));
    LocalMux I__6892 (
            .O(N__29261),
            .I(N__29255));
    LocalMux I__6891 (
            .O(N__29258),
            .I(N__29252));
    Span4Mux_h I__6890 (
            .O(N__29255),
            .I(N__29249));
    Span4Mux_h I__6889 (
            .O(N__29252),
            .I(N__29246));
    Odrv4 I__6888 (
            .O(N__29249),
            .I(\this_ppu.M_state_q_RNI42KTAZ0Z_0 ));
    Odrv4 I__6887 (
            .O(N__29246),
            .I(\this_ppu.M_state_q_RNI42KTAZ0Z_0 ));
    CascadeMux I__6886 (
            .O(N__29241),
            .I(N__29238));
    InMux I__6885 (
            .O(N__29238),
            .I(N__29235));
    LocalMux I__6884 (
            .O(N__29235),
            .I(N__29232));
    Span4Mux_h I__6883 (
            .O(N__29232),
            .I(N__29229));
    Odrv4 I__6882 (
            .O(N__29229),
            .I(M_this_data_tmp_qZ0Z_4));
    InMux I__6881 (
            .O(N__29226),
            .I(N__29223));
    LocalMux I__6880 (
            .O(N__29223),
            .I(N__29220));
    Span4Mux_h I__6879 (
            .O(N__29220),
            .I(N__29217));
    Odrv4 I__6878 (
            .O(N__29217),
            .I(N_71_0));
    InMux I__6877 (
            .O(N__29214),
            .I(N__29210));
    InMux I__6876 (
            .O(N__29213),
            .I(N__29207));
    LocalMux I__6875 (
            .O(N__29210),
            .I(N__29204));
    LocalMux I__6874 (
            .O(N__29207),
            .I(\this_ppu.M_this_ppu_vram_addr_i_7 ));
    Odrv4 I__6873 (
            .O(N__29204),
            .I(\this_ppu.M_this_ppu_vram_addr_i_7 ));
    InMux I__6872 (
            .O(N__29199),
            .I(N__29194));
    CascadeMux I__6871 (
            .O(N__29198),
            .I(N__29190));
    CascadeMux I__6870 (
            .O(N__29197),
            .I(N__29187));
    LocalMux I__6869 (
            .O(N__29194),
            .I(N__29184));
    InMux I__6868 (
            .O(N__29193),
            .I(N__29181));
    InMux I__6867 (
            .O(N__29190),
            .I(N__29178));
    InMux I__6866 (
            .O(N__29187),
            .I(N__29175));
    Span4Mux_h I__6865 (
            .O(N__29184),
            .I(N__29172));
    LocalMux I__6864 (
            .O(N__29181),
            .I(N__29167));
    LocalMux I__6863 (
            .O(N__29178),
            .I(N__29167));
    LocalMux I__6862 (
            .O(N__29175),
            .I(N__29164));
    Span4Mux_v I__6861 (
            .O(N__29172),
            .I(N__29161));
    Span4Mux_h I__6860 (
            .O(N__29167),
            .I(N__29158));
    Span4Mux_h I__6859 (
            .O(N__29164),
            .I(N__29155));
    Odrv4 I__6858 (
            .O(N__29161),
            .I(M_this_oam_ram_read_data_16));
    Odrv4 I__6857 (
            .O(N__29158),
            .I(M_this_oam_ram_read_data_16));
    Odrv4 I__6856 (
            .O(N__29155),
            .I(M_this_oam_ram_read_data_16));
    InMux I__6855 (
            .O(N__29148),
            .I(N__29144));
    InMux I__6854 (
            .O(N__29147),
            .I(N__29141));
    LocalMux I__6853 (
            .O(N__29144),
            .I(N__29138));
    LocalMux I__6852 (
            .O(N__29141),
            .I(\this_ppu.M_vaddress_q_i_1 ));
    Odrv4 I__6851 (
            .O(N__29138),
            .I(\this_ppu.M_vaddress_q_i_1 ));
    InMux I__6850 (
            .O(N__29133),
            .I(N__29129));
    InMux I__6849 (
            .O(N__29132),
            .I(N__29126));
    LocalMux I__6848 (
            .O(N__29129),
            .I(N__29123));
    LocalMux I__6847 (
            .O(N__29126),
            .I(\this_ppu.M_vaddress_q_i_2 ));
    Odrv4 I__6846 (
            .O(N__29123),
            .I(\this_ppu.M_vaddress_q_i_2 ));
    CascadeMux I__6845 (
            .O(N__29118),
            .I(N__29113));
    CascadeMux I__6844 (
            .O(N__29117),
            .I(N__29110));
    InMux I__6843 (
            .O(N__29116),
            .I(N__29107));
    InMux I__6842 (
            .O(N__29113),
            .I(N__29104));
    InMux I__6841 (
            .O(N__29110),
            .I(N__29101));
    LocalMux I__6840 (
            .O(N__29107),
            .I(N__29098));
    LocalMux I__6839 (
            .O(N__29104),
            .I(N__29095));
    LocalMux I__6838 (
            .O(N__29101),
            .I(N__29092));
    Span4Mux_h I__6837 (
            .O(N__29098),
            .I(N__29089));
    Span4Mux_v I__6836 (
            .O(N__29095),
            .I(N__29086));
    Span4Mux_h I__6835 (
            .O(N__29092),
            .I(N__29083));
    Odrv4 I__6834 (
            .O(N__29089),
            .I(M_this_oam_ram_read_data_18));
    Odrv4 I__6833 (
            .O(N__29086),
            .I(M_this_oam_ram_read_data_18));
    Odrv4 I__6832 (
            .O(N__29083),
            .I(M_this_oam_ram_read_data_18));
    CascadeMux I__6831 (
            .O(N__29076),
            .I(N__29073));
    InMux I__6830 (
            .O(N__29073),
            .I(N__29070));
    LocalMux I__6829 (
            .O(N__29070),
            .I(N__29067));
    Odrv4 I__6828 (
            .O(N__29067),
            .I(M_this_data_tmp_qZ0Z_15));
    InMux I__6827 (
            .O(N__29064),
            .I(N__29061));
    LocalMux I__6826 (
            .O(N__29061),
            .I(N__29058));
    Span4Mux_v I__6825 (
            .O(N__29058),
            .I(N__29055));
    Sp12to4 I__6824 (
            .O(N__29055),
            .I(N__29052));
    Odrv12 I__6823 (
            .O(N__29052),
            .I(M_this_oam_ram_write_data_15));
    CascadeMux I__6822 (
            .O(N__29049),
            .I(N__29046));
    InMux I__6821 (
            .O(N__29046),
            .I(N__29043));
    LocalMux I__6820 (
            .O(N__29043),
            .I(\this_ppu.M_this_oam_ram_read_data_i_16 ));
    InMux I__6819 (
            .O(N__29040),
            .I(N__29037));
    LocalMux I__6818 (
            .O(N__29037),
            .I(\this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0 ));
    InMux I__6817 (
            .O(N__29034),
            .I(\this_ppu.un2_vscroll_cry_0 ));
    InMux I__6816 (
            .O(N__29031),
            .I(\this_ppu.un2_vscroll_cry_1 ));
    CascadeMux I__6815 (
            .O(N__29028),
            .I(N__29025));
    InMux I__6814 (
            .O(N__29025),
            .I(N__29022));
    LocalMux I__6813 (
            .O(N__29022),
            .I(N__29019));
    Span4Mux_v I__6812 (
            .O(N__29019),
            .I(N__29016));
    Sp12to4 I__6811 (
            .O(N__29016),
            .I(N__29013));
    Span12Mux_h I__6810 (
            .O(N__29013),
            .I(N__29010));
    Span12Mux_v I__6809 (
            .O(N__29010),
            .I(N__29007));
    Odrv12 I__6808 (
            .O(N__29007),
            .I(M_this_map_ram_read_data_6));
    CascadeMux I__6807 (
            .O(N__29004),
            .I(N__29000));
    InMux I__6806 (
            .O(N__29003),
            .I(N__28996));
    InMux I__6805 (
            .O(N__29000),
            .I(N__28993));
    InMux I__6804 (
            .O(N__28999),
            .I(N__28990));
    LocalMux I__6803 (
            .O(N__28996),
            .I(N__28986));
    LocalMux I__6802 (
            .O(N__28993),
            .I(N__28983));
    LocalMux I__6801 (
            .O(N__28990),
            .I(N__28980));
    InMux I__6800 (
            .O(N__28989),
            .I(N__28977));
    Span4Mux_h I__6799 (
            .O(N__28986),
            .I(N__28974));
    Span4Mux_v I__6798 (
            .O(N__28983),
            .I(N__28967));
    Span4Mux_h I__6797 (
            .O(N__28980),
            .I(N__28967));
    LocalMux I__6796 (
            .O(N__28977),
            .I(N__28967));
    Span4Mux_h I__6795 (
            .O(N__28974),
            .I(N__28964));
    Span4Mux_h I__6794 (
            .O(N__28967),
            .I(N__28961));
    Odrv4 I__6793 (
            .O(N__28964),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    Odrv4 I__6792 (
            .O(N__28961),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    InMux I__6791 (
            .O(N__28956),
            .I(N__28953));
    LocalMux I__6790 (
            .O(N__28953),
            .I(\this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0 ));
    CascadeMux I__6789 (
            .O(N__28950),
            .I(N__28945));
    CascadeMux I__6788 (
            .O(N__28949),
            .I(N__28941));
    CascadeMux I__6787 (
            .O(N__28948),
            .I(N__28938));
    InMux I__6786 (
            .O(N__28945),
            .I(N__28934));
    CascadeMux I__6785 (
            .O(N__28944),
            .I(N__28931));
    InMux I__6784 (
            .O(N__28941),
            .I(N__28927));
    InMux I__6783 (
            .O(N__28938),
            .I(N__28924));
    CascadeMux I__6782 (
            .O(N__28937),
            .I(N__28921));
    LocalMux I__6781 (
            .O(N__28934),
            .I(N__28915));
    InMux I__6780 (
            .O(N__28931),
            .I(N__28912));
    CascadeMux I__6779 (
            .O(N__28930),
            .I(N__28909));
    LocalMux I__6778 (
            .O(N__28927),
            .I(N__28906));
    LocalMux I__6777 (
            .O(N__28924),
            .I(N__28903));
    InMux I__6776 (
            .O(N__28921),
            .I(N__28900));
    CascadeMux I__6775 (
            .O(N__28920),
            .I(N__28897));
    CascadeMux I__6774 (
            .O(N__28919),
            .I(N__28893));
    CascadeMux I__6773 (
            .O(N__28918),
            .I(N__28890));
    Span4Mux_h I__6772 (
            .O(N__28915),
            .I(N__28885));
    LocalMux I__6771 (
            .O(N__28912),
            .I(N__28882));
    InMux I__6770 (
            .O(N__28909),
            .I(N__28879));
    Span4Mux_h I__6769 (
            .O(N__28906),
            .I(N__28875));
    Span4Mux_v I__6768 (
            .O(N__28903),
            .I(N__28870));
    LocalMux I__6767 (
            .O(N__28900),
            .I(N__28870));
    InMux I__6766 (
            .O(N__28897),
            .I(N__28867));
    CascadeMux I__6765 (
            .O(N__28896),
            .I(N__28864));
    InMux I__6764 (
            .O(N__28893),
            .I(N__28861));
    InMux I__6763 (
            .O(N__28890),
            .I(N__28858));
    CascadeMux I__6762 (
            .O(N__28889),
            .I(N__28855));
    CascadeMux I__6761 (
            .O(N__28888),
            .I(N__28852));
    Span4Mux_v I__6760 (
            .O(N__28885),
            .I(N__28845));
    Span4Mux_h I__6759 (
            .O(N__28882),
            .I(N__28845));
    LocalMux I__6758 (
            .O(N__28879),
            .I(N__28842));
    CascadeMux I__6757 (
            .O(N__28878),
            .I(N__28838));
    Span4Mux_h I__6756 (
            .O(N__28875),
            .I(N__28835));
    Span4Mux_v I__6755 (
            .O(N__28870),
            .I(N__28830));
    LocalMux I__6754 (
            .O(N__28867),
            .I(N__28830));
    InMux I__6753 (
            .O(N__28864),
            .I(N__28827));
    LocalMux I__6752 (
            .O(N__28861),
            .I(N__28822));
    LocalMux I__6751 (
            .O(N__28858),
            .I(N__28822));
    InMux I__6750 (
            .O(N__28855),
            .I(N__28819));
    InMux I__6749 (
            .O(N__28852),
            .I(N__28816));
    CascadeMux I__6748 (
            .O(N__28851),
            .I(N__28813));
    CascadeMux I__6747 (
            .O(N__28850),
            .I(N__28810));
    Span4Mux_v I__6746 (
            .O(N__28845),
            .I(N__28805));
    Span4Mux_h I__6745 (
            .O(N__28842),
            .I(N__28805));
    CascadeMux I__6744 (
            .O(N__28841),
            .I(N__28802));
    InMux I__6743 (
            .O(N__28838),
            .I(N__28799));
    Span4Mux_h I__6742 (
            .O(N__28835),
            .I(N__28796));
    Span4Mux_h I__6741 (
            .O(N__28830),
            .I(N__28791));
    LocalMux I__6740 (
            .O(N__28827),
            .I(N__28791));
    Span4Mux_v I__6739 (
            .O(N__28822),
            .I(N__28784));
    LocalMux I__6738 (
            .O(N__28819),
            .I(N__28784));
    LocalMux I__6737 (
            .O(N__28816),
            .I(N__28784));
    InMux I__6736 (
            .O(N__28813),
            .I(N__28781));
    InMux I__6735 (
            .O(N__28810),
            .I(N__28778));
    Span4Mux_h I__6734 (
            .O(N__28805),
            .I(N__28775));
    InMux I__6733 (
            .O(N__28802),
            .I(N__28772));
    LocalMux I__6732 (
            .O(N__28799),
            .I(N__28769));
    Span4Mux_h I__6731 (
            .O(N__28796),
            .I(N__28766));
    Span4Mux_v I__6730 (
            .O(N__28791),
            .I(N__28763));
    Span4Mux_v I__6729 (
            .O(N__28784),
            .I(N__28758));
    LocalMux I__6728 (
            .O(N__28781),
            .I(N__28758));
    LocalMux I__6727 (
            .O(N__28778),
            .I(N__28755));
    Span4Mux_h I__6726 (
            .O(N__28775),
            .I(N__28752));
    LocalMux I__6725 (
            .O(N__28772),
            .I(N__28749));
    Span12Mux_s9_h I__6724 (
            .O(N__28769),
            .I(N__28746));
    Span4Mux_v I__6723 (
            .O(N__28766),
            .I(N__28739));
    Span4Mux_v I__6722 (
            .O(N__28763),
            .I(N__28739));
    Span4Mux_v I__6721 (
            .O(N__28758),
            .I(N__28739));
    Span4Mux_h I__6720 (
            .O(N__28755),
            .I(N__28736));
    Span4Mux_h I__6719 (
            .O(N__28752),
            .I(N__28731));
    Span4Mux_h I__6718 (
            .O(N__28749),
            .I(N__28731));
    Odrv12 I__6717 (
            .O(N__28746),
            .I(M_this_ppu_sprites_addr_5));
    Odrv4 I__6716 (
            .O(N__28739),
            .I(M_this_ppu_sprites_addr_5));
    Odrv4 I__6715 (
            .O(N__28736),
            .I(M_this_ppu_sprites_addr_5));
    Odrv4 I__6714 (
            .O(N__28731),
            .I(M_this_ppu_sprites_addr_5));
    CascadeMux I__6713 (
            .O(N__28722),
            .I(N__28717));
    CascadeMux I__6712 (
            .O(N__28721),
            .I(N__28712));
    InMux I__6711 (
            .O(N__28720),
            .I(N__28708));
    InMux I__6710 (
            .O(N__28717),
            .I(N__28705));
    InMux I__6709 (
            .O(N__28716),
            .I(N__28702));
    InMux I__6708 (
            .O(N__28715),
            .I(N__28699));
    InMux I__6707 (
            .O(N__28712),
            .I(N__28694));
    InMux I__6706 (
            .O(N__28711),
            .I(N__28694));
    LocalMux I__6705 (
            .O(N__28708),
            .I(N__28689));
    LocalMux I__6704 (
            .O(N__28705),
            .I(N__28689));
    LocalMux I__6703 (
            .O(N__28702),
            .I(N__28686));
    LocalMux I__6702 (
            .O(N__28699),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    LocalMux I__6701 (
            .O(N__28694),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv4 I__6700 (
            .O(N__28689),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv4 I__6699 (
            .O(N__28686),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    CascadeMux I__6698 (
            .O(N__28677),
            .I(N__28673));
    InMux I__6697 (
            .O(N__28676),
            .I(N__28669));
    InMux I__6696 (
            .O(N__28673),
            .I(N__28665));
    InMux I__6695 (
            .O(N__28672),
            .I(N__28660));
    LocalMux I__6694 (
            .O(N__28669),
            .I(N__28657));
    CascadeMux I__6693 (
            .O(N__28668),
            .I(N__28654));
    LocalMux I__6692 (
            .O(N__28665),
            .I(N__28651));
    InMux I__6691 (
            .O(N__28664),
            .I(N__28646));
    InMux I__6690 (
            .O(N__28663),
            .I(N__28646));
    LocalMux I__6689 (
            .O(N__28660),
            .I(N__28643));
    Span4Mux_h I__6688 (
            .O(N__28657),
            .I(N__28639));
    InMux I__6687 (
            .O(N__28654),
            .I(N__28636));
    Span4Mux_h I__6686 (
            .O(N__28651),
            .I(N__28633));
    LocalMux I__6685 (
            .O(N__28646),
            .I(N__28628));
    Span4Mux_h I__6684 (
            .O(N__28643),
            .I(N__28628));
    InMux I__6683 (
            .O(N__28642),
            .I(N__28625));
    Span4Mux_h I__6682 (
            .O(N__28639),
            .I(N__28622));
    LocalMux I__6681 (
            .O(N__28636),
            .I(N__28617));
    Span4Mux_h I__6680 (
            .O(N__28633),
            .I(N__28617));
    Span4Mux_h I__6679 (
            .O(N__28628),
            .I(N__28614));
    LocalMux I__6678 (
            .O(N__28625),
            .I(\this_ppu.N_132_0 ));
    Odrv4 I__6677 (
            .O(N__28622),
            .I(\this_ppu.N_132_0 ));
    Odrv4 I__6676 (
            .O(N__28617),
            .I(\this_ppu.N_132_0 ));
    Odrv4 I__6675 (
            .O(N__28614),
            .I(\this_ppu.N_132_0 ));
    InMux I__6674 (
            .O(N__28605),
            .I(N__28602));
    LocalMux I__6673 (
            .O(N__28602),
            .I(N__28599));
    Span4Mux_h I__6672 (
            .O(N__28599),
            .I(N__28596));
    Odrv4 I__6671 (
            .O(N__28596),
            .I(N_56_0));
    CascadeMux I__6670 (
            .O(N__28593),
            .I(N__28590));
    InMux I__6669 (
            .O(N__28590),
            .I(N__28587));
    LocalMux I__6668 (
            .O(N__28587),
            .I(M_this_data_tmp_qZ0Z_13));
    CascadeMux I__6667 (
            .O(N__28584),
            .I(N__28580));
    CascadeMux I__6666 (
            .O(N__28583),
            .I(N__28576));
    InMux I__6665 (
            .O(N__28580),
            .I(N__28571));
    InMux I__6664 (
            .O(N__28579),
            .I(N__28571));
    InMux I__6663 (
            .O(N__28576),
            .I(N__28568));
    LocalMux I__6662 (
            .O(N__28571),
            .I(N__28562));
    LocalMux I__6661 (
            .O(N__28568),
            .I(N__28562));
    InMux I__6660 (
            .O(N__28567),
            .I(N__28558));
    Span4Mux_v I__6659 (
            .O(N__28562),
            .I(N__28554));
    InMux I__6658 (
            .O(N__28561),
            .I(N__28551));
    LocalMux I__6657 (
            .O(N__28558),
            .I(N__28548));
    InMux I__6656 (
            .O(N__28557),
            .I(N__28545));
    Span4Mux_h I__6655 (
            .O(N__28554),
            .I(N__28542));
    LocalMux I__6654 (
            .O(N__28551),
            .I(N__28539));
    Span4Mux_h I__6653 (
            .O(N__28548),
            .I(N__28534));
    LocalMux I__6652 (
            .O(N__28545),
            .I(N__28534));
    Odrv4 I__6651 (
            .O(N__28542),
            .I(M_this_state_d21_1));
    Odrv12 I__6650 (
            .O(N__28539),
            .I(M_this_state_d21_1));
    Odrv4 I__6649 (
            .O(N__28534),
            .I(M_this_state_d21_1));
    InMux I__6648 (
            .O(N__28527),
            .I(N__28524));
    LocalMux I__6647 (
            .O(N__28524),
            .I(N__28521));
    Span4Mux_v I__6646 (
            .O(N__28521),
            .I(N__28516));
    InMux I__6645 (
            .O(N__28520),
            .I(N__28511));
    InMux I__6644 (
            .O(N__28519),
            .I(N__28511));
    Sp12to4 I__6643 (
            .O(N__28516),
            .I(N__28506));
    LocalMux I__6642 (
            .O(N__28511),
            .I(N__28506));
    Odrv12 I__6641 (
            .O(N__28506),
            .I(port_address_in_4));
    InMux I__6640 (
            .O(N__28503),
            .I(N__28495));
    InMux I__6639 (
            .O(N__28502),
            .I(N__28495));
    InMux I__6638 (
            .O(N__28501),
            .I(N__28490));
    InMux I__6637 (
            .O(N__28500),
            .I(N__28490));
    LocalMux I__6636 (
            .O(N__28495),
            .I(N__28485));
    LocalMux I__6635 (
            .O(N__28490),
            .I(N__28485));
    Sp12to4 I__6634 (
            .O(N__28485),
            .I(N__28482));
    Odrv12 I__6633 (
            .O(N__28482),
            .I(port_address_in_2));
    CascadeMux I__6632 (
            .O(N__28479),
            .I(N__28475));
    InMux I__6631 (
            .O(N__28478),
            .I(N__28470));
    InMux I__6630 (
            .O(N__28475),
            .I(N__28470));
    LocalMux I__6629 (
            .O(N__28470),
            .I(N__28467));
    Odrv4 I__6628 (
            .O(N__28467),
            .I(M_this_state_d21_6_x));
    InMux I__6627 (
            .O(N__28464),
            .I(N__28461));
    LocalMux I__6626 (
            .O(N__28461),
            .I(N__28458));
    Odrv4 I__6625 (
            .O(N__28458),
            .I(M_this_substate_q_RNOZ0Z_2));
    CascadeMux I__6624 (
            .O(N__28455),
            .I(N__28451));
    InMux I__6623 (
            .O(N__28454),
            .I(N__28447));
    InMux I__6622 (
            .O(N__28451),
            .I(N__28442));
    InMux I__6621 (
            .O(N__28450),
            .I(N__28442));
    LocalMux I__6620 (
            .O(N__28447),
            .I(N__28436));
    LocalMux I__6619 (
            .O(N__28442),
            .I(N__28436));
    InMux I__6618 (
            .O(N__28441),
            .I(N__28433));
    Span4Mux_v I__6617 (
            .O(N__28436),
            .I(N__28428));
    LocalMux I__6616 (
            .O(N__28433),
            .I(N__28428));
    Span4Mux_h I__6615 (
            .O(N__28428),
            .I(N__28425));
    Span4Mux_v I__6614 (
            .O(N__28425),
            .I(N__28422));
    Span4Mux_h I__6613 (
            .O(N__28422),
            .I(N__28419));
    Odrv4 I__6612 (
            .O(N__28419),
            .I(port_address_in_3));
    CascadeMux I__6611 (
            .O(N__28416),
            .I(N__28411));
    CascadeMux I__6610 (
            .O(N__28415),
            .I(N__28408));
    InMux I__6609 (
            .O(N__28414),
            .I(N__28404));
    InMux I__6608 (
            .O(N__28411),
            .I(N__28399));
    InMux I__6607 (
            .O(N__28408),
            .I(N__28399));
    InMux I__6606 (
            .O(N__28407),
            .I(N__28396));
    LocalMux I__6605 (
            .O(N__28404),
            .I(N__28391));
    LocalMux I__6604 (
            .O(N__28399),
            .I(N__28386));
    LocalMux I__6603 (
            .O(N__28396),
            .I(N__28386));
    InMux I__6602 (
            .O(N__28395),
            .I(N__28383));
    InMux I__6601 (
            .O(N__28394),
            .I(N__28379));
    Span4Mux_h I__6600 (
            .O(N__28391),
            .I(N__28374));
    Span4Mux_h I__6599 (
            .O(N__28386),
            .I(N__28374));
    LocalMux I__6598 (
            .O(N__28383),
            .I(N__28371));
    InMux I__6597 (
            .O(N__28382),
            .I(N__28368));
    LocalMux I__6596 (
            .O(N__28379),
            .I(N__28365));
    Span4Mux_h I__6595 (
            .O(N__28374),
            .I(N__28357));
    Span4Mux_v I__6594 (
            .O(N__28371),
            .I(N__28357));
    LocalMux I__6593 (
            .O(N__28368),
            .I(N__28357));
    Span4Mux_v I__6592 (
            .O(N__28365),
            .I(N__28354));
    InMux I__6591 (
            .O(N__28364),
            .I(N__28351));
    Span4Mux_h I__6590 (
            .O(N__28357),
            .I(N__28348));
    Sp12to4 I__6589 (
            .O(N__28354),
            .I(N__28343));
    LocalMux I__6588 (
            .O(N__28351),
            .I(N__28343));
    Span4Mux_v I__6587 (
            .O(N__28348),
            .I(N__28340));
    Span12Mux_h I__6586 (
            .O(N__28343),
            .I(N__28337));
    Span4Mux_v I__6585 (
            .O(N__28340),
            .I(N__28334));
    Odrv12 I__6584 (
            .O(N__28337),
            .I(port_address_in_1));
    Odrv4 I__6583 (
            .O(N__28334),
            .I(port_address_in_1));
    CascadeMux I__6582 (
            .O(N__28329),
            .I(N__28326));
    InMux I__6581 (
            .O(N__28326),
            .I(N__28323));
    LocalMux I__6580 (
            .O(N__28323),
            .I(N__28320));
    Span4Mux_v I__6579 (
            .O(N__28320),
            .I(N__28317));
    Odrv4 I__6578 (
            .O(N__28317),
            .I(\this_vga_signals.M_this_state_d24Z0Z_1 ));
    CEMux I__6577 (
            .O(N__28314),
            .I(N__28310));
    CEMux I__6576 (
            .O(N__28313),
            .I(N__28307));
    LocalMux I__6575 (
            .O(N__28310),
            .I(N__28304));
    LocalMux I__6574 (
            .O(N__28307),
            .I(N__28301));
    Span4Mux_h I__6573 (
            .O(N__28304),
            .I(N__28298));
    Span4Mux_h I__6572 (
            .O(N__28301),
            .I(N__28295));
    Span4Mux_v I__6571 (
            .O(N__28298),
            .I(N__28292));
    Span4Mux_v I__6570 (
            .O(N__28295),
            .I(N__28289));
    Odrv4 I__6569 (
            .O(N__28292),
            .I(\this_sprites_ram.mem_WE_0 ));
    Odrv4 I__6568 (
            .O(N__28289),
            .I(\this_sprites_ram.mem_WE_0 ));
    CascadeMux I__6567 (
            .O(N__28284),
            .I(N__28280));
    InMux I__6566 (
            .O(N__28283),
            .I(N__28277));
    InMux I__6565 (
            .O(N__28280),
            .I(N__28274));
    LocalMux I__6564 (
            .O(N__28277),
            .I(\this_ppu.M_this_ppu_map_addr_i_1 ));
    LocalMux I__6563 (
            .O(N__28274),
            .I(\this_ppu.M_this_ppu_map_addr_i_1 ));
    InMux I__6562 (
            .O(N__28269),
            .I(N__28265));
    InMux I__6561 (
            .O(N__28268),
            .I(N__28262));
    LocalMux I__6560 (
            .O(N__28265),
            .I(\this_ppu.M_this_ppu_map_addr_i_2 ));
    LocalMux I__6559 (
            .O(N__28262),
            .I(\this_ppu.M_this_ppu_map_addr_i_2 ));
    InMux I__6558 (
            .O(N__28257),
            .I(N__28253));
    InMux I__6557 (
            .O(N__28256),
            .I(N__28250));
    LocalMux I__6556 (
            .O(N__28253),
            .I(\this_ppu.M_this_ppu_map_addr_i_3 ));
    LocalMux I__6555 (
            .O(N__28250),
            .I(\this_ppu.M_this_ppu_map_addr_i_3 ));
    CascadeMux I__6554 (
            .O(N__28245),
            .I(N__28242));
    InMux I__6553 (
            .O(N__28242),
            .I(N__28238));
    InMux I__6552 (
            .O(N__28241),
            .I(N__28235));
    LocalMux I__6551 (
            .O(N__28238),
            .I(\this_ppu.M_this_ppu_map_addr_i_4 ));
    LocalMux I__6550 (
            .O(N__28235),
            .I(\this_ppu.M_this_ppu_map_addr_i_4 ));
    InMux I__6549 (
            .O(N__28230),
            .I(bfn_22_20_0_));
    InMux I__6548 (
            .O(N__28227),
            .I(N__28224));
    LocalMux I__6547 (
            .O(N__28224),
            .I(\this_ppu.vscroll8_1 ));
    InMux I__6546 (
            .O(N__28221),
            .I(N__28218));
    LocalMux I__6545 (
            .O(N__28218),
            .I(N__28215));
    Span4Mux_h I__6544 (
            .O(N__28215),
            .I(N__28211));
    InMux I__6543 (
            .O(N__28214),
            .I(N__28208));
    Span4Mux_h I__6542 (
            .O(N__28211),
            .I(N__28205));
    LocalMux I__6541 (
            .O(N__28208),
            .I(N__28202));
    IoSpan4Mux I__6540 (
            .O(N__28205),
            .I(N__28199));
    Span12Mux_h I__6539 (
            .O(N__28202),
            .I(N__28196));
    Odrv4 I__6538 (
            .O(N__28199),
            .I(port_address_in_5));
    Odrv12 I__6537 (
            .O(N__28196),
            .I(port_address_in_5));
    InMux I__6536 (
            .O(N__28191),
            .I(N__28188));
    LocalMux I__6535 (
            .O(N__28188),
            .I(N__28184));
    InMux I__6534 (
            .O(N__28187),
            .I(N__28181));
    Span4Mux_h I__6533 (
            .O(N__28184),
            .I(N__28176));
    LocalMux I__6532 (
            .O(N__28181),
            .I(N__28176));
    Span4Mux_v I__6531 (
            .O(N__28176),
            .I(N__28173));
    Sp12to4 I__6530 (
            .O(N__28173),
            .I(N__28170));
    Odrv12 I__6529 (
            .O(N__28170),
            .I(port_address_in_6));
    CascadeMux I__6528 (
            .O(N__28167),
            .I(N__28164));
    InMux I__6527 (
            .O(N__28164),
            .I(N__28161));
    LocalMux I__6526 (
            .O(N__28161),
            .I(N__28157));
    InMux I__6525 (
            .O(N__28160),
            .I(N__28154));
    Span4Mux_v I__6524 (
            .O(N__28157),
            .I(N__28151));
    LocalMux I__6523 (
            .O(N__28154),
            .I(N__28148));
    Sp12to4 I__6522 (
            .O(N__28151),
            .I(N__28143));
    Span12Mux_v I__6521 (
            .O(N__28148),
            .I(N__28143));
    Span12Mux_v I__6520 (
            .O(N__28143),
            .I(N__28140));
    Odrv12 I__6519 (
            .O(N__28140),
            .I(port_address_in_7));
    InMux I__6518 (
            .O(N__28137),
            .I(N__28134));
    LocalMux I__6517 (
            .O(N__28134),
            .I(N__28130));
    InMux I__6516 (
            .O(N__28133),
            .I(N__28127));
    Span4Mux_h I__6515 (
            .O(N__28130),
            .I(N__28121));
    LocalMux I__6514 (
            .O(N__28127),
            .I(N__28121));
    InMux I__6513 (
            .O(N__28126),
            .I(N__28115));
    Span4Mux_h I__6512 (
            .O(N__28121),
            .I(N__28112));
    InMux I__6511 (
            .O(N__28120),
            .I(N__28109));
    InMux I__6510 (
            .O(N__28119),
            .I(N__28106));
    InMux I__6509 (
            .O(N__28118),
            .I(N__28103));
    LocalMux I__6508 (
            .O(N__28115),
            .I(M_this_state_qZ0Z_12));
    Odrv4 I__6507 (
            .O(N__28112),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__6506 (
            .O(N__28109),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__6505 (
            .O(N__28106),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__6504 (
            .O(N__28103),
            .I(M_this_state_qZ0Z_12));
    InMux I__6503 (
            .O(N__28092),
            .I(bfn_22_18_0_));
    InMux I__6502 (
            .O(N__28089),
            .I(N__28086));
    LocalMux I__6501 (
            .O(N__28086),
            .I(\this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO ));
    CascadeMux I__6500 (
            .O(N__28083),
            .I(N__28080));
    InMux I__6499 (
            .O(N__28080),
            .I(N__28077));
    LocalMux I__6498 (
            .O(N__28077),
            .I(N__28074));
    Odrv4 I__6497 (
            .O(N__28074),
            .I(\this_ppu.un1_M_haddress_q_2_5 ));
    CascadeMux I__6496 (
            .O(N__28071),
            .I(un1_M_this_oam_address_q_c3_cascade_));
    CascadeMux I__6495 (
            .O(N__28068),
            .I(N__28065));
    InMux I__6494 (
            .O(N__28065),
            .I(N__28062));
    LocalMux I__6493 (
            .O(N__28062),
            .I(N__28059));
    Odrv12 I__6492 (
            .O(N__28059),
            .I(M_this_data_tmp_qZ0Z_7));
    InMux I__6491 (
            .O(N__28056),
            .I(N__28053));
    LocalMux I__6490 (
            .O(N__28053),
            .I(N__28050));
    Span4Mux_h I__6489 (
            .O(N__28050),
            .I(N__28047));
    Odrv4 I__6488 (
            .O(N__28047),
            .I(N_65_0));
    InMux I__6487 (
            .O(N__28044),
            .I(N__28040));
    InMux I__6486 (
            .O(N__28043),
            .I(N__28037));
    LocalMux I__6485 (
            .O(N__28040),
            .I(\this_ppu.M_this_ppu_vram_addr_i_0 ));
    LocalMux I__6484 (
            .O(N__28037),
            .I(\this_ppu.M_this_ppu_vram_addr_i_0 ));
    CascadeMux I__6483 (
            .O(N__28032),
            .I(N__28027));
    InMux I__6482 (
            .O(N__28031),
            .I(N__28023));
    InMux I__6481 (
            .O(N__28030),
            .I(N__28020));
    InMux I__6480 (
            .O(N__28027),
            .I(N__28017));
    CascadeMux I__6479 (
            .O(N__28026),
            .I(N__28014));
    LocalMux I__6478 (
            .O(N__28023),
            .I(N__28007));
    LocalMux I__6477 (
            .O(N__28020),
            .I(N__28007));
    LocalMux I__6476 (
            .O(N__28017),
            .I(N__28007));
    InMux I__6475 (
            .O(N__28014),
            .I(N__28004));
    Span4Mux_v I__6474 (
            .O(N__28007),
            .I(N__27999));
    LocalMux I__6473 (
            .O(N__28004),
            .I(N__27999));
    Span4Mux_h I__6472 (
            .O(N__27999),
            .I(N__27996));
    Odrv4 I__6471 (
            .O(N__27996),
            .I(M_this_oam_ram_read_data_8));
    InMux I__6470 (
            .O(N__27993),
            .I(N__27989));
    InMux I__6469 (
            .O(N__27992),
            .I(N__27986));
    LocalMux I__6468 (
            .O(N__27989),
            .I(\this_ppu.M_this_ppu_vram_addr_i_1 ));
    LocalMux I__6467 (
            .O(N__27986),
            .I(\this_ppu.M_this_ppu_vram_addr_i_1 ));
    CascadeMux I__6466 (
            .O(N__27981),
            .I(N__27977));
    InMux I__6465 (
            .O(N__27980),
            .I(N__27973));
    InMux I__6464 (
            .O(N__27977),
            .I(N__27970));
    CascadeMux I__6463 (
            .O(N__27976),
            .I(N__27967));
    LocalMux I__6462 (
            .O(N__27973),
            .I(N__27962));
    LocalMux I__6461 (
            .O(N__27970),
            .I(N__27962));
    InMux I__6460 (
            .O(N__27967),
            .I(N__27959));
    Span4Mux_v I__6459 (
            .O(N__27962),
            .I(N__27954));
    LocalMux I__6458 (
            .O(N__27959),
            .I(N__27954));
    Span4Mux_h I__6457 (
            .O(N__27954),
            .I(N__27951));
    Odrv4 I__6456 (
            .O(N__27951),
            .I(M_this_oam_ram_read_data_9));
    InMux I__6455 (
            .O(N__27948),
            .I(N__27944));
    InMux I__6454 (
            .O(N__27947),
            .I(N__27941));
    LocalMux I__6453 (
            .O(N__27944),
            .I(\this_ppu.M_this_ppu_vram_addr_i_2 ));
    LocalMux I__6452 (
            .O(N__27941),
            .I(\this_ppu.M_this_ppu_vram_addr_i_2 ));
    CascadeMux I__6451 (
            .O(N__27936),
            .I(N__27933));
    InMux I__6450 (
            .O(N__27933),
            .I(N__27928));
    CascadeMux I__6449 (
            .O(N__27932),
            .I(N__27925));
    InMux I__6448 (
            .O(N__27931),
            .I(N__27922));
    LocalMux I__6447 (
            .O(N__27928),
            .I(N__27919));
    InMux I__6446 (
            .O(N__27925),
            .I(N__27916));
    LocalMux I__6445 (
            .O(N__27922),
            .I(N__27913));
    Span4Mux_v I__6444 (
            .O(N__27919),
            .I(N__27908));
    LocalMux I__6443 (
            .O(N__27916),
            .I(N__27908));
    Span4Mux_h I__6442 (
            .O(N__27913),
            .I(N__27905));
    Span4Mux_h I__6441 (
            .O(N__27908),
            .I(N__27902));
    Odrv4 I__6440 (
            .O(N__27905),
            .I(M_this_oam_ram_read_data_10));
    Odrv4 I__6439 (
            .O(N__27902),
            .I(M_this_oam_ram_read_data_10));
    CascadeMux I__6438 (
            .O(N__27897),
            .I(N__27893));
    InMux I__6437 (
            .O(N__27896),
            .I(N__27890));
    InMux I__6436 (
            .O(N__27893),
            .I(N__27887));
    LocalMux I__6435 (
            .O(N__27890),
            .I(\this_ppu.M_this_ppu_map_addr_i_0 ));
    LocalMux I__6434 (
            .O(N__27887),
            .I(\this_ppu.M_this_ppu_map_addr_i_0 ));
    InMux I__6433 (
            .O(N__27882),
            .I(N__27873));
    InMux I__6432 (
            .O(N__27881),
            .I(N__27873));
    InMux I__6431 (
            .O(N__27880),
            .I(N__27873));
    LocalMux I__6430 (
            .O(N__27873),
            .I(\this_ppu.un1_M_vaddress_q_2_c5 ));
    CascadeMux I__6429 (
            .O(N__27870),
            .I(N__27867));
    CascadeBuf I__6428 (
            .O(N__27867),
            .I(N__27864));
    CascadeMux I__6427 (
            .O(N__27864),
            .I(N__27861));
    InMux I__6426 (
            .O(N__27861),
            .I(N__27858));
    LocalMux I__6425 (
            .O(N__27858),
            .I(N__27854));
    InMux I__6424 (
            .O(N__27857),
            .I(N__27848));
    Span12Mux_h I__6423 (
            .O(N__27854),
            .I(N__27845));
    InMux I__6422 (
            .O(N__27853),
            .I(N__27838));
    InMux I__6421 (
            .O(N__27852),
            .I(N__27838));
    InMux I__6420 (
            .O(N__27851),
            .I(N__27838));
    LocalMux I__6419 (
            .O(N__27848),
            .I(N__27835));
    Span12Mux_v I__6418 (
            .O(N__27845),
            .I(N__27832));
    LocalMux I__6417 (
            .O(N__27838),
            .I(M_this_ppu_map_addr_7));
    Odrv4 I__6416 (
            .O(N__27835),
            .I(M_this_ppu_map_addr_7));
    Odrv12 I__6415 (
            .O(N__27832),
            .I(M_this_ppu_map_addr_7));
    CascadeMux I__6414 (
            .O(N__27825),
            .I(N__27822));
    CascadeBuf I__6413 (
            .O(N__27822),
            .I(N__27819));
    CascadeMux I__6412 (
            .O(N__27819),
            .I(N__27816));
    InMux I__6411 (
            .O(N__27816),
            .I(N__27813));
    LocalMux I__6410 (
            .O(N__27813),
            .I(N__27810));
    Sp12to4 I__6409 (
            .O(N__27810),
            .I(N__27805));
    CascadeMux I__6408 (
            .O(N__27809),
            .I(N__27802));
    InMux I__6407 (
            .O(N__27808),
            .I(N__27798));
    Span12Mux_h I__6406 (
            .O(N__27805),
            .I(N__27795));
    InMux I__6405 (
            .O(N__27802),
            .I(N__27790));
    InMux I__6404 (
            .O(N__27801),
            .I(N__27790));
    LocalMux I__6403 (
            .O(N__27798),
            .I(N__27787));
    Span12Mux_v I__6402 (
            .O(N__27795),
            .I(N__27784));
    LocalMux I__6401 (
            .O(N__27790),
            .I(M_this_ppu_map_addr_8));
    Odrv4 I__6400 (
            .O(N__27787),
            .I(M_this_ppu_map_addr_8));
    Odrv12 I__6399 (
            .O(N__27784),
            .I(M_this_ppu_map_addr_8));
    CascadeMux I__6398 (
            .O(N__27777),
            .I(N__27774));
    CascadeBuf I__6397 (
            .O(N__27774),
            .I(N__27771));
    CascadeMux I__6396 (
            .O(N__27771),
            .I(N__27768));
    InMux I__6395 (
            .O(N__27768),
            .I(N__27765));
    LocalMux I__6394 (
            .O(N__27765),
            .I(N__27761));
    InMux I__6393 (
            .O(N__27764),
            .I(N__27757));
    Span12Mux_h I__6392 (
            .O(N__27761),
            .I(N__27754));
    InMux I__6391 (
            .O(N__27760),
            .I(N__27751));
    LocalMux I__6390 (
            .O(N__27757),
            .I(N__27748));
    Span12Mux_v I__6389 (
            .O(N__27754),
            .I(N__27745));
    LocalMux I__6388 (
            .O(N__27751),
            .I(M_this_ppu_map_addr_9));
    Odrv4 I__6387 (
            .O(N__27748),
            .I(M_this_ppu_map_addr_9));
    Odrv12 I__6386 (
            .O(N__27745),
            .I(M_this_ppu_map_addr_9));
    InMux I__6385 (
            .O(N__27738),
            .I(N__27735));
    LocalMux I__6384 (
            .O(N__27735),
            .I(N__27732));
    Odrv4 I__6383 (
            .O(N__27732),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4 ));
    InMux I__6382 (
            .O(N__27729),
            .I(N__27716));
    InMux I__6381 (
            .O(N__27728),
            .I(N__27716));
    InMux I__6380 (
            .O(N__27727),
            .I(N__27707));
    InMux I__6379 (
            .O(N__27726),
            .I(N__27707));
    InMux I__6378 (
            .O(N__27725),
            .I(N__27707));
    InMux I__6377 (
            .O(N__27724),
            .I(N__27707));
    InMux I__6376 (
            .O(N__27723),
            .I(N__27704));
    InMux I__6375 (
            .O(N__27722),
            .I(N__27697));
    InMux I__6374 (
            .O(N__27721),
            .I(N__27697));
    LocalMux I__6373 (
            .O(N__27716),
            .I(N__27692));
    LocalMux I__6372 (
            .O(N__27707),
            .I(N__27692));
    LocalMux I__6371 (
            .O(N__27704),
            .I(N__27689));
    InMux I__6370 (
            .O(N__27703),
            .I(N__27686));
    InMux I__6369 (
            .O(N__27702),
            .I(N__27680));
    LocalMux I__6368 (
            .O(N__27697),
            .I(N__27677));
    Span4Mux_v I__6367 (
            .O(N__27692),
            .I(N__27670));
    Span4Mux_h I__6366 (
            .O(N__27689),
            .I(N__27670));
    LocalMux I__6365 (
            .O(N__27686),
            .I(N__27670));
    InMux I__6364 (
            .O(N__27685),
            .I(N__27663));
    InMux I__6363 (
            .O(N__27684),
            .I(N__27663));
    InMux I__6362 (
            .O(N__27683),
            .I(N__27663));
    LocalMux I__6361 (
            .O(N__27680),
            .I(\this_vga_signals.un1_M_this_state_q_14_0 ));
    Odrv4 I__6360 (
            .O(N__27677),
            .I(\this_vga_signals.un1_M_this_state_q_14_0 ));
    Odrv4 I__6359 (
            .O(N__27670),
            .I(\this_vga_signals.un1_M_this_state_q_14_0 ));
    LocalMux I__6358 (
            .O(N__27663),
            .I(\this_vga_signals.un1_M_this_state_q_14_0 ));
    CascadeMux I__6357 (
            .O(N__27654),
            .I(N__27651));
    InMux I__6356 (
            .O(N__27651),
            .I(N__27648));
    LocalMux I__6355 (
            .O(N__27648),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_4 ));
    InMux I__6354 (
            .O(N__27645),
            .I(N__27642));
    LocalMux I__6353 (
            .O(N__27642),
            .I(N__27639));
    Span4Mux_h I__6352 (
            .O(N__27639),
            .I(N__27636));
    Odrv4 I__6351 (
            .O(N__27636),
            .I(un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0));
    CascadeMux I__6350 (
            .O(N__27633),
            .I(N__27630));
    InMux I__6349 (
            .O(N__27630),
            .I(N__27626));
    CascadeMux I__6348 (
            .O(N__27629),
            .I(N__27623));
    LocalMux I__6347 (
            .O(N__27626),
            .I(N__27619));
    InMux I__6346 (
            .O(N__27623),
            .I(N__27616));
    CascadeMux I__6345 (
            .O(N__27622),
            .I(N__27613));
    Span4Mux_h I__6344 (
            .O(N__27619),
            .I(N__27606));
    LocalMux I__6343 (
            .O(N__27616),
            .I(N__27606));
    InMux I__6342 (
            .O(N__27613),
            .I(N__27603));
    CascadeMux I__6341 (
            .O(N__27612),
            .I(N__27600));
    CascadeMux I__6340 (
            .O(N__27611),
            .I(N__27596));
    Span4Mux_v I__6339 (
            .O(N__27606),
            .I(N__27591));
    LocalMux I__6338 (
            .O(N__27603),
            .I(N__27591));
    InMux I__6337 (
            .O(N__27600),
            .I(N__27588));
    CascadeMux I__6336 (
            .O(N__27599),
            .I(N__27585));
    InMux I__6335 (
            .O(N__27596),
            .I(N__27581));
    Span4Mux_h I__6334 (
            .O(N__27591),
            .I(N__27575));
    LocalMux I__6333 (
            .O(N__27588),
            .I(N__27575));
    InMux I__6332 (
            .O(N__27585),
            .I(N__27572));
    CascadeMux I__6331 (
            .O(N__27584),
            .I(N__27569));
    LocalMux I__6330 (
            .O(N__27581),
            .I(N__27565));
    CascadeMux I__6329 (
            .O(N__27580),
            .I(N__27562));
    Span4Mux_v I__6328 (
            .O(N__27575),
            .I(N__27556));
    LocalMux I__6327 (
            .O(N__27572),
            .I(N__27556));
    InMux I__6326 (
            .O(N__27569),
            .I(N__27553));
    CascadeMux I__6325 (
            .O(N__27568),
            .I(N__27550));
    Span4Mux_h I__6324 (
            .O(N__27565),
            .I(N__27545));
    InMux I__6323 (
            .O(N__27562),
            .I(N__27542));
    CascadeMux I__6322 (
            .O(N__27561),
            .I(N__27539));
    Span4Mux_h I__6321 (
            .O(N__27556),
            .I(N__27533));
    LocalMux I__6320 (
            .O(N__27553),
            .I(N__27533));
    InMux I__6319 (
            .O(N__27550),
            .I(N__27530));
    CascadeMux I__6318 (
            .O(N__27549),
            .I(N__27526));
    CascadeMux I__6317 (
            .O(N__27548),
            .I(N__27523));
    Span4Mux_v I__6316 (
            .O(N__27545),
            .I(N__27517));
    LocalMux I__6315 (
            .O(N__27542),
            .I(N__27517));
    InMux I__6314 (
            .O(N__27539),
            .I(N__27514));
    CascadeMux I__6313 (
            .O(N__27538),
            .I(N__27511));
    Span4Mux_v I__6312 (
            .O(N__27533),
            .I(N__27506));
    LocalMux I__6311 (
            .O(N__27530),
            .I(N__27506));
    CascadeMux I__6310 (
            .O(N__27529),
            .I(N__27503));
    InMux I__6309 (
            .O(N__27526),
            .I(N__27500));
    InMux I__6308 (
            .O(N__27523),
            .I(N__27497));
    CascadeMux I__6307 (
            .O(N__27522),
            .I(N__27494));
    Span4Mux_h I__6306 (
            .O(N__27517),
            .I(N__27488));
    LocalMux I__6305 (
            .O(N__27514),
            .I(N__27488));
    InMux I__6304 (
            .O(N__27511),
            .I(N__27485));
    Span4Mux_h I__6303 (
            .O(N__27506),
            .I(N__27482));
    InMux I__6302 (
            .O(N__27503),
            .I(N__27479));
    LocalMux I__6301 (
            .O(N__27500),
            .I(N__27476));
    LocalMux I__6300 (
            .O(N__27497),
            .I(N__27473));
    InMux I__6299 (
            .O(N__27494),
            .I(N__27470));
    CascadeMux I__6298 (
            .O(N__27493),
            .I(N__27467));
    Span4Mux_v I__6297 (
            .O(N__27488),
            .I(N__27461));
    LocalMux I__6296 (
            .O(N__27485),
            .I(N__27461));
    Span4Mux_v I__6295 (
            .O(N__27482),
            .I(N__27456));
    LocalMux I__6294 (
            .O(N__27479),
            .I(N__27456));
    Span4Mux_v I__6293 (
            .O(N__27476),
            .I(N__27449));
    Span4Mux_h I__6292 (
            .O(N__27473),
            .I(N__27449));
    LocalMux I__6291 (
            .O(N__27470),
            .I(N__27449));
    InMux I__6290 (
            .O(N__27467),
            .I(N__27446));
    InMux I__6289 (
            .O(N__27466),
            .I(N__27442));
    Sp12to4 I__6288 (
            .O(N__27461),
            .I(N__27438));
    Span4Mux_v I__6287 (
            .O(N__27456),
            .I(N__27431));
    Span4Mux_v I__6286 (
            .O(N__27449),
            .I(N__27431));
    LocalMux I__6285 (
            .O(N__27446),
            .I(N__27431));
    InMux I__6284 (
            .O(N__27445),
            .I(N__27428));
    LocalMux I__6283 (
            .O(N__27442),
            .I(N__27425));
    InMux I__6282 (
            .O(N__27441),
            .I(N__27422));
    Span12Mux_h I__6281 (
            .O(N__27438),
            .I(N__27415));
    Sp12to4 I__6280 (
            .O(N__27431),
            .I(N__27415));
    LocalMux I__6279 (
            .O(N__27428),
            .I(N__27415));
    Span4Mux_h I__6278 (
            .O(N__27425),
            .I(N__27412));
    LocalMux I__6277 (
            .O(N__27422),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv12 I__6276 (
            .O(N__27415),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv4 I__6275 (
            .O(N__27412),
            .I(M_this_sprites_address_qZ0Z_4));
    InMux I__6274 (
            .O(N__27405),
            .I(N__27401));
    InMux I__6273 (
            .O(N__27404),
            .I(N__27396));
    LocalMux I__6272 (
            .O(N__27401),
            .I(N__27393));
    InMux I__6271 (
            .O(N__27400),
            .I(N__27390));
    InMux I__6270 (
            .O(N__27399),
            .I(N__27387));
    LocalMux I__6269 (
            .O(N__27396),
            .I(N__27384));
    Span4Mux_v I__6268 (
            .O(N__27393),
            .I(N__27379));
    LocalMux I__6267 (
            .O(N__27390),
            .I(N__27379));
    LocalMux I__6266 (
            .O(N__27387),
            .I(N__27376));
    Odrv4 I__6265 (
            .O(N__27384),
            .I(\this_vga_signals.M_this_state_q_ns_8 ));
    Odrv4 I__6264 (
            .O(N__27379),
            .I(\this_vga_signals.M_this_state_q_ns_8 ));
    Odrv4 I__6263 (
            .O(N__27376),
            .I(\this_vga_signals.M_this_state_q_ns_8 ));
    InMux I__6262 (
            .O(N__27369),
            .I(N__27365));
    InMux I__6261 (
            .O(N__27368),
            .I(N__27362));
    LocalMux I__6260 (
            .O(N__27365),
            .I(N__27357));
    LocalMux I__6259 (
            .O(N__27362),
            .I(N__27354));
    InMux I__6258 (
            .O(N__27361),
            .I(N__27351));
    CascadeMux I__6257 (
            .O(N__27360),
            .I(N__27347));
    Span4Mux_h I__6256 (
            .O(N__27357),
            .I(N__27344));
    Span4Mux_v I__6255 (
            .O(N__27354),
            .I(N__27341));
    LocalMux I__6254 (
            .O(N__27351),
            .I(N__27338));
    InMux I__6253 (
            .O(N__27350),
            .I(N__27335));
    InMux I__6252 (
            .O(N__27347),
            .I(N__27332));
    Odrv4 I__6251 (
            .O(N__27344),
            .I(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ));
    Odrv4 I__6250 (
            .O(N__27341),
            .I(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ));
    Odrv12 I__6249 (
            .O(N__27338),
            .I(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ));
    LocalMux I__6248 (
            .O(N__27335),
            .I(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ));
    LocalMux I__6247 (
            .O(N__27332),
            .I(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ));
    InMux I__6246 (
            .O(N__27321),
            .I(N__27318));
    LocalMux I__6245 (
            .O(N__27318),
            .I(N__27313));
    InMux I__6244 (
            .O(N__27317),
            .I(N__27310));
    InMux I__6243 (
            .O(N__27316),
            .I(N__27306));
    Span4Mux_h I__6242 (
            .O(N__27313),
            .I(N__27302));
    LocalMux I__6241 (
            .O(N__27310),
            .I(N__27299));
    InMux I__6240 (
            .O(N__27309),
            .I(N__27296));
    LocalMux I__6239 (
            .O(N__27306),
            .I(N__27292));
    InMux I__6238 (
            .O(N__27305),
            .I(N__27289));
    Span4Mux_v I__6237 (
            .O(N__27302),
            .I(N__27284));
    Span4Mux_h I__6236 (
            .O(N__27299),
            .I(N__27284));
    LocalMux I__6235 (
            .O(N__27296),
            .I(N__27281));
    InMux I__6234 (
            .O(N__27295),
            .I(N__27278));
    Span4Mux_v I__6233 (
            .O(N__27292),
            .I(N__27273));
    LocalMux I__6232 (
            .O(N__27289),
            .I(N__27273));
    Span4Mux_v I__6231 (
            .O(N__27284),
            .I(N__27268));
    Span4Mux_h I__6230 (
            .O(N__27281),
            .I(N__27268));
    LocalMux I__6229 (
            .O(N__27278),
            .I(N__27265));
    Span4Mux_v I__6228 (
            .O(N__27273),
            .I(N__27260));
    Span4Mux_v I__6227 (
            .O(N__27268),
            .I(N__27255));
    Span4Mux_h I__6226 (
            .O(N__27265),
            .I(N__27255));
    InMux I__6225 (
            .O(N__27264),
            .I(N__27252));
    InMux I__6224 (
            .O(N__27263),
            .I(N__27249));
    Span4Mux_h I__6223 (
            .O(N__27260),
            .I(N__27246));
    Span4Mux_v I__6222 (
            .O(N__27255),
            .I(N__27243));
    LocalMux I__6221 (
            .O(N__27252),
            .I(N__27240));
    LocalMux I__6220 (
            .O(N__27249),
            .I(N__27237));
    Sp12to4 I__6219 (
            .O(N__27246),
            .I(N__27234));
    Span4Mux_v I__6218 (
            .O(N__27243),
            .I(N__27227));
    Span4Mux_h I__6217 (
            .O(N__27240),
            .I(N__27227));
    Span4Mux_h I__6216 (
            .O(N__27237),
            .I(N__27227));
    Odrv12 I__6215 (
            .O(N__27234),
            .I(M_this_sprites_ram_write_data_1));
    Odrv4 I__6214 (
            .O(N__27227),
            .I(M_this_sprites_ram_write_data_1));
    InMux I__6213 (
            .O(N__27222),
            .I(N__27219));
    LocalMux I__6212 (
            .O(N__27219),
            .I(N__27216));
    Span12Mux_v I__6211 (
            .O(N__27216),
            .I(N__27213));
    Span12Mux_h I__6210 (
            .O(N__27213),
            .I(N__27210));
    Span12Mux_v I__6209 (
            .O(N__27210),
            .I(N__27207));
    Odrv12 I__6208 (
            .O(N__27207),
            .I(M_this_map_ram_read_data_4));
    CascadeMux I__6207 (
            .O(N__27204),
            .I(N__27197));
    CascadeMux I__6206 (
            .O(N__27203),
            .I(N__27193));
    CascadeMux I__6205 (
            .O(N__27202),
            .I(N__27190));
    CascadeMux I__6204 (
            .O(N__27201),
            .I(N__27186));
    CascadeMux I__6203 (
            .O(N__27200),
            .I(N__27183));
    InMux I__6202 (
            .O(N__27197),
            .I(N__27179));
    CascadeMux I__6201 (
            .O(N__27196),
            .I(N__27176));
    InMux I__6200 (
            .O(N__27193),
            .I(N__27172));
    InMux I__6199 (
            .O(N__27190),
            .I(N__27169));
    CascadeMux I__6198 (
            .O(N__27189),
            .I(N__27166));
    InMux I__6197 (
            .O(N__27186),
            .I(N__27161));
    InMux I__6196 (
            .O(N__27183),
            .I(N__27158));
    CascadeMux I__6195 (
            .O(N__27182),
            .I(N__27155));
    LocalMux I__6194 (
            .O(N__27179),
            .I(N__27151));
    InMux I__6193 (
            .O(N__27176),
            .I(N__27148));
    CascadeMux I__6192 (
            .O(N__27175),
            .I(N__27145));
    LocalMux I__6191 (
            .O(N__27172),
            .I(N__27141));
    LocalMux I__6190 (
            .O(N__27169),
            .I(N__27138));
    InMux I__6189 (
            .O(N__27166),
            .I(N__27135));
    CascadeMux I__6188 (
            .O(N__27165),
            .I(N__27132));
    CascadeMux I__6187 (
            .O(N__27164),
            .I(N__27128));
    LocalMux I__6186 (
            .O(N__27161),
            .I(N__27123));
    LocalMux I__6185 (
            .O(N__27158),
            .I(N__27123));
    InMux I__6184 (
            .O(N__27155),
            .I(N__27120));
    CascadeMux I__6183 (
            .O(N__27154),
            .I(N__27116));
    Span4Mux_v I__6182 (
            .O(N__27151),
            .I(N__27111));
    LocalMux I__6181 (
            .O(N__27148),
            .I(N__27111));
    InMux I__6180 (
            .O(N__27145),
            .I(N__27108));
    CascadeMux I__6179 (
            .O(N__27144),
            .I(N__27105));
    Span4Mux_v I__6178 (
            .O(N__27141),
            .I(N__27098));
    Span4Mux_h I__6177 (
            .O(N__27138),
            .I(N__27098));
    LocalMux I__6176 (
            .O(N__27135),
            .I(N__27098));
    InMux I__6175 (
            .O(N__27132),
            .I(N__27095));
    CascadeMux I__6174 (
            .O(N__27131),
            .I(N__27092));
    InMux I__6173 (
            .O(N__27128),
            .I(N__27089));
    Span4Mux_v I__6172 (
            .O(N__27123),
            .I(N__27084));
    LocalMux I__6171 (
            .O(N__27120),
            .I(N__27084));
    CascadeMux I__6170 (
            .O(N__27119),
            .I(N__27081));
    InMux I__6169 (
            .O(N__27116),
            .I(N__27077));
    Span4Mux_h I__6168 (
            .O(N__27111),
            .I(N__27072));
    LocalMux I__6167 (
            .O(N__27108),
            .I(N__27072));
    InMux I__6166 (
            .O(N__27105),
            .I(N__27069));
    Span4Mux_v I__6165 (
            .O(N__27098),
            .I(N__27064));
    LocalMux I__6164 (
            .O(N__27095),
            .I(N__27064));
    InMux I__6163 (
            .O(N__27092),
            .I(N__27061));
    LocalMux I__6162 (
            .O(N__27089),
            .I(N__27058));
    Span4Mux_v I__6161 (
            .O(N__27084),
            .I(N__27055));
    InMux I__6160 (
            .O(N__27081),
            .I(N__27052));
    CascadeMux I__6159 (
            .O(N__27080),
            .I(N__27049));
    LocalMux I__6158 (
            .O(N__27077),
            .I(N__27046));
    Span4Mux_v I__6157 (
            .O(N__27072),
            .I(N__27041));
    LocalMux I__6156 (
            .O(N__27069),
            .I(N__27041));
    Span4Mux_h I__6155 (
            .O(N__27064),
            .I(N__27038));
    LocalMux I__6154 (
            .O(N__27061),
            .I(N__27035));
    Span12Mux_h I__6153 (
            .O(N__27058),
            .I(N__27032));
    Sp12to4 I__6152 (
            .O(N__27055),
            .I(N__27027));
    LocalMux I__6151 (
            .O(N__27052),
            .I(N__27027));
    InMux I__6150 (
            .O(N__27049),
            .I(N__27024));
    Span12Mux_s10_h I__6149 (
            .O(N__27046),
            .I(N__27021));
    Span4Mux_h I__6148 (
            .O(N__27041),
            .I(N__27018));
    Span4Mux_v I__6147 (
            .O(N__27038),
            .I(N__27013));
    Span4Mux_h I__6146 (
            .O(N__27035),
            .I(N__27013));
    Span12Mux_v I__6145 (
            .O(N__27032),
            .I(N__27006));
    Span12Mux_h I__6144 (
            .O(N__27027),
            .I(N__27006));
    LocalMux I__6143 (
            .O(N__27024),
            .I(N__27006));
    Odrv12 I__6142 (
            .O(N__27021),
            .I(M_this_ppu_sprites_addr_10));
    Odrv4 I__6141 (
            .O(N__27018),
            .I(M_this_ppu_sprites_addr_10));
    Odrv4 I__6140 (
            .O(N__27013),
            .I(M_this_ppu_sprites_addr_10));
    Odrv12 I__6139 (
            .O(N__27006),
            .I(M_this_ppu_sprites_addr_10));
    CascadeMux I__6138 (
            .O(N__26997),
            .I(N__26993));
    CascadeMux I__6137 (
            .O(N__26996),
            .I(N__26987));
    InMux I__6136 (
            .O(N__26993),
            .I(N__26982));
    CascadeMux I__6135 (
            .O(N__26992),
            .I(N__26979));
    CascadeMux I__6134 (
            .O(N__26991),
            .I(N__26974));
    CascadeMux I__6133 (
            .O(N__26990),
            .I(N__26971));
    InMux I__6132 (
            .O(N__26987),
            .I(N__26967));
    CascadeMux I__6131 (
            .O(N__26986),
            .I(N__26964));
    CascadeMux I__6130 (
            .O(N__26985),
            .I(N__26961));
    LocalMux I__6129 (
            .O(N__26982),
            .I(N__26957));
    InMux I__6128 (
            .O(N__26979),
            .I(N__26954));
    CascadeMux I__6127 (
            .O(N__26978),
            .I(N__26951));
    CascadeMux I__6126 (
            .O(N__26977),
            .I(N__26948));
    InMux I__6125 (
            .O(N__26974),
            .I(N__26943));
    InMux I__6124 (
            .O(N__26971),
            .I(N__26940));
    CascadeMux I__6123 (
            .O(N__26970),
            .I(N__26937));
    LocalMux I__6122 (
            .O(N__26967),
            .I(N__26934));
    InMux I__6121 (
            .O(N__26964),
            .I(N__26931));
    InMux I__6120 (
            .O(N__26961),
            .I(N__26928));
    CascadeMux I__6119 (
            .O(N__26960),
            .I(N__26925));
    Span4Mux_h I__6118 (
            .O(N__26957),
            .I(N__26920));
    LocalMux I__6117 (
            .O(N__26954),
            .I(N__26920));
    InMux I__6116 (
            .O(N__26951),
            .I(N__26917));
    InMux I__6115 (
            .O(N__26948),
            .I(N__26914));
    CascadeMux I__6114 (
            .O(N__26947),
            .I(N__26911));
    CascadeMux I__6113 (
            .O(N__26946),
            .I(N__26908));
    LocalMux I__6112 (
            .O(N__26943),
            .I(N__26904));
    LocalMux I__6111 (
            .O(N__26940),
            .I(N__26901));
    InMux I__6110 (
            .O(N__26937),
            .I(N__26898));
    Span4Mux_v I__6109 (
            .O(N__26934),
            .I(N__26892));
    LocalMux I__6108 (
            .O(N__26931),
            .I(N__26892));
    LocalMux I__6107 (
            .O(N__26928),
            .I(N__26889));
    InMux I__6106 (
            .O(N__26925),
            .I(N__26886));
    Span4Mux_v I__6105 (
            .O(N__26920),
            .I(N__26879));
    LocalMux I__6104 (
            .O(N__26917),
            .I(N__26879));
    LocalMux I__6103 (
            .O(N__26914),
            .I(N__26879));
    InMux I__6102 (
            .O(N__26911),
            .I(N__26876));
    InMux I__6101 (
            .O(N__26908),
            .I(N__26873));
    CascadeMux I__6100 (
            .O(N__26907),
            .I(N__26870));
    Span4Mux_v I__6099 (
            .O(N__26904),
            .I(N__26863));
    Span4Mux_v I__6098 (
            .O(N__26901),
            .I(N__26863));
    LocalMux I__6097 (
            .O(N__26898),
            .I(N__26863));
    CascadeMux I__6096 (
            .O(N__26897),
            .I(N__26860));
    Span4Mux_h I__6095 (
            .O(N__26892),
            .I(N__26856));
    Span4Mux_v I__6094 (
            .O(N__26889),
            .I(N__26851));
    LocalMux I__6093 (
            .O(N__26886),
            .I(N__26851));
    Span4Mux_v I__6092 (
            .O(N__26879),
            .I(N__26846));
    LocalMux I__6091 (
            .O(N__26876),
            .I(N__26846));
    LocalMux I__6090 (
            .O(N__26873),
            .I(N__26843));
    InMux I__6089 (
            .O(N__26870),
            .I(N__26840));
    Span4Mux_v I__6088 (
            .O(N__26863),
            .I(N__26837));
    InMux I__6087 (
            .O(N__26860),
            .I(N__26834));
    CascadeMux I__6086 (
            .O(N__26859),
            .I(N__26831));
    Span4Mux_v I__6085 (
            .O(N__26856),
            .I(N__26826));
    Span4Mux_h I__6084 (
            .O(N__26851),
            .I(N__26826));
    Span4Mux_h I__6083 (
            .O(N__26846),
            .I(N__26823));
    Span4Mux_v I__6082 (
            .O(N__26843),
            .I(N__26818));
    LocalMux I__6081 (
            .O(N__26840),
            .I(N__26818));
    Sp12to4 I__6080 (
            .O(N__26837),
            .I(N__26813));
    LocalMux I__6079 (
            .O(N__26834),
            .I(N__26813));
    InMux I__6078 (
            .O(N__26831),
            .I(N__26810));
    Span4Mux_v I__6077 (
            .O(N__26826),
            .I(N__26803));
    Span4Mux_v I__6076 (
            .O(N__26823),
            .I(N__26803));
    Span4Mux_h I__6075 (
            .O(N__26818),
            .I(N__26803));
    Span12Mux_h I__6074 (
            .O(N__26813),
            .I(N__26798));
    LocalMux I__6073 (
            .O(N__26810),
            .I(N__26798));
    Odrv4 I__6072 (
            .O(N__26803),
            .I(M_this_ppu_sprites_addr_4));
    Odrv12 I__6071 (
            .O(N__26798),
            .I(M_this_ppu_sprites_addr_4));
    CEMux I__6070 (
            .O(N__26793),
            .I(N__26790));
    LocalMux I__6069 (
            .O(N__26790),
            .I(N__26787));
    Span4Mux_v I__6068 (
            .O(N__26787),
            .I(N__26783));
    CEMux I__6067 (
            .O(N__26786),
            .I(N__26780));
    Span4Mux_h I__6066 (
            .O(N__26783),
            .I(N__26777));
    LocalMux I__6065 (
            .O(N__26780),
            .I(N__26774));
    Span4Mux_h I__6064 (
            .O(N__26777),
            .I(N__26771));
    Span4Mux_v I__6063 (
            .O(N__26774),
            .I(N__26768));
    Span4Mux_h I__6062 (
            .O(N__26771),
            .I(N__26763));
    Span4Mux_h I__6061 (
            .O(N__26768),
            .I(N__26763));
    Odrv4 I__6060 (
            .O(N__26763),
            .I(\this_sprites_ram.mem_WE_4 ));
    CascadeMux I__6059 (
            .O(N__26760),
            .I(N__26757));
    InMux I__6058 (
            .O(N__26757),
            .I(N__26754));
    LocalMux I__6057 (
            .O(N__26754),
            .I(N__26751));
    Odrv12 I__6056 (
            .O(N__26751),
            .I(M_this_state_d22));
    InMux I__6055 (
            .O(N__26748),
            .I(N__26745));
    LocalMux I__6054 (
            .O(N__26745),
            .I(N__26742));
    Odrv4 I__6053 (
            .O(N__26742),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11 ));
    InMux I__6052 (
            .O(N__26739),
            .I(N__26736));
    LocalMux I__6051 (
            .O(N__26736),
            .I(N__26732));
    InMux I__6050 (
            .O(N__26735),
            .I(N__26728));
    Span4Mux_v I__6049 (
            .O(N__26732),
            .I(N__26722));
    InMux I__6048 (
            .O(N__26731),
            .I(N__26719));
    LocalMux I__6047 (
            .O(N__26728),
            .I(N__26716));
    InMux I__6046 (
            .O(N__26727),
            .I(N__26709));
    InMux I__6045 (
            .O(N__26726),
            .I(N__26709));
    InMux I__6044 (
            .O(N__26725),
            .I(N__26709));
    Sp12to4 I__6043 (
            .O(N__26722),
            .I(N__26703));
    LocalMux I__6042 (
            .O(N__26719),
            .I(N__26703));
    Span4Mux_h I__6041 (
            .O(N__26716),
            .I(N__26698));
    LocalMux I__6040 (
            .O(N__26709),
            .I(N__26698));
    InMux I__6039 (
            .O(N__26708),
            .I(N__26695));
    Span12Mux_h I__6038 (
            .O(N__26703),
            .I(N__26690));
    Sp12to4 I__6037 (
            .O(N__26698),
            .I(N__26690));
    LocalMux I__6036 (
            .O(N__26695),
            .I(N__26687));
    Odrv12 I__6035 (
            .O(N__26690),
            .I(port_address_in_0));
    Odrv12 I__6034 (
            .O(N__26687),
            .I(port_address_in_0));
    CascadeMux I__6033 (
            .O(N__26682),
            .I(N__26678));
    InMux I__6032 (
            .O(N__26681),
            .I(N__26673));
    InMux I__6031 (
            .O(N__26678),
            .I(N__26673));
    LocalMux I__6030 (
            .O(N__26673),
            .I(\this_vga_signals.M_this_state_d21Z0Z_6 ));
    CascadeMux I__6029 (
            .O(N__26670),
            .I(N__26667));
    InMux I__6028 (
            .O(N__26667),
            .I(N__26663));
    CascadeMux I__6027 (
            .O(N__26666),
            .I(N__26660));
    LocalMux I__6026 (
            .O(N__26663),
            .I(N__26657));
    InMux I__6025 (
            .O(N__26660),
            .I(N__26654));
    Span4Mux_v I__6024 (
            .O(N__26657),
            .I(N__26651));
    LocalMux I__6023 (
            .O(N__26654),
            .I(N__26648));
    Span4Mux_h I__6022 (
            .O(N__26651),
            .I(N__26643));
    Span4Mux_v I__6021 (
            .O(N__26648),
            .I(N__26643));
    Odrv4 I__6020 (
            .O(N__26643),
            .I(\this_vga_signals.M_this_state_dZ0Z24 ));
    InMux I__6019 (
            .O(N__26640),
            .I(N__26637));
    LocalMux I__6018 (
            .O(N__26637),
            .I(N__26634));
    Odrv4 I__6017 (
            .O(N__26634),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8 ));
    CascadeMux I__6016 (
            .O(N__26631),
            .I(N__26628));
    InMux I__6015 (
            .O(N__26628),
            .I(N__26625));
    LocalMux I__6014 (
            .O(N__26625),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_8 ));
    InMux I__6013 (
            .O(N__26622),
            .I(N__26619));
    LocalMux I__6012 (
            .O(N__26619),
            .I(N__26616));
    Odrv4 I__6011 (
            .O(N__26616),
            .I(un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0));
    CascadeMux I__6010 (
            .O(N__26613),
            .I(N__26610));
    InMux I__6009 (
            .O(N__26610),
            .I(N__26605));
    CascadeMux I__6008 (
            .O(N__26609),
            .I(N__26602));
    CascadeMux I__6007 (
            .O(N__26608),
            .I(N__26599));
    LocalMux I__6006 (
            .O(N__26605),
            .I(N__26594));
    InMux I__6005 (
            .O(N__26602),
            .I(N__26591));
    InMux I__6004 (
            .O(N__26599),
            .I(N__26588));
    CascadeMux I__6003 (
            .O(N__26598),
            .I(N__26585));
    CascadeMux I__6002 (
            .O(N__26597),
            .I(N__26581));
    Span4Mux_h I__6001 (
            .O(N__26594),
            .I(N__26573));
    LocalMux I__6000 (
            .O(N__26591),
            .I(N__26573));
    LocalMux I__5999 (
            .O(N__26588),
            .I(N__26570));
    InMux I__5998 (
            .O(N__26585),
            .I(N__26567));
    CascadeMux I__5997 (
            .O(N__26584),
            .I(N__26564));
    InMux I__5996 (
            .O(N__26581),
            .I(N__26558));
    CascadeMux I__5995 (
            .O(N__26580),
            .I(N__26555));
    CascadeMux I__5994 (
            .O(N__26579),
            .I(N__26552));
    CascadeMux I__5993 (
            .O(N__26578),
            .I(N__26549));
    Span4Mux_v I__5992 (
            .O(N__26573),
            .I(N__26542));
    Span4Mux_h I__5991 (
            .O(N__26570),
            .I(N__26542));
    LocalMux I__5990 (
            .O(N__26567),
            .I(N__26542));
    InMux I__5989 (
            .O(N__26564),
            .I(N__26539));
    CascadeMux I__5988 (
            .O(N__26563),
            .I(N__26536));
    CascadeMux I__5987 (
            .O(N__26562),
            .I(N__26532));
    CascadeMux I__5986 (
            .O(N__26561),
            .I(N__26529));
    LocalMux I__5985 (
            .O(N__26558),
            .I(N__26524));
    InMux I__5984 (
            .O(N__26555),
            .I(N__26521));
    InMux I__5983 (
            .O(N__26552),
            .I(N__26518));
    InMux I__5982 (
            .O(N__26549),
            .I(N__26515));
    Span4Mux_v I__5981 (
            .O(N__26542),
            .I(N__26510));
    LocalMux I__5980 (
            .O(N__26539),
            .I(N__26510));
    InMux I__5979 (
            .O(N__26536),
            .I(N__26507));
    CascadeMux I__5978 (
            .O(N__26535),
            .I(N__26504));
    InMux I__5977 (
            .O(N__26532),
            .I(N__26501));
    InMux I__5976 (
            .O(N__26529),
            .I(N__26498));
    CascadeMux I__5975 (
            .O(N__26528),
            .I(N__26495));
    CascadeMux I__5974 (
            .O(N__26527),
            .I(N__26492));
    Span4Mux_v I__5973 (
            .O(N__26524),
            .I(N__26486));
    LocalMux I__5972 (
            .O(N__26521),
            .I(N__26486));
    LocalMux I__5971 (
            .O(N__26518),
            .I(N__26481));
    LocalMux I__5970 (
            .O(N__26515),
            .I(N__26481));
    Span4Mux_h I__5969 (
            .O(N__26510),
            .I(N__26476));
    LocalMux I__5968 (
            .O(N__26507),
            .I(N__26476));
    InMux I__5967 (
            .O(N__26504),
            .I(N__26473));
    LocalMux I__5966 (
            .O(N__26501),
            .I(N__26470));
    LocalMux I__5965 (
            .O(N__26498),
            .I(N__26467));
    InMux I__5964 (
            .O(N__26495),
            .I(N__26464));
    InMux I__5963 (
            .O(N__26492),
            .I(N__26461));
    CascadeMux I__5962 (
            .O(N__26491),
            .I(N__26458));
    Span4Mux_v I__5961 (
            .O(N__26486),
            .I(N__26453));
    Span4Mux_v I__5960 (
            .O(N__26481),
            .I(N__26453));
    Span4Mux_v I__5959 (
            .O(N__26476),
            .I(N__26448));
    LocalMux I__5958 (
            .O(N__26473),
            .I(N__26448));
    Span4Mux_v I__5957 (
            .O(N__26470),
            .I(N__26441));
    Span4Mux_h I__5956 (
            .O(N__26467),
            .I(N__26441));
    LocalMux I__5955 (
            .O(N__26464),
            .I(N__26441));
    LocalMux I__5954 (
            .O(N__26461),
            .I(N__26438));
    InMux I__5953 (
            .O(N__26458),
            .I(N__26435));
    Sp12to4 I__5952 (
            .O(N__26453),
            .I(N__26430));
    Span4Mux_h I__5951 (
            .O(N__26448),
            .I(N__26427));
    Span4Mux_v I__5950 (
            .O(N__26441),
            .I(N__26420));
    Span4Mux_v I__5949 (
            .O(N__26438),
            .I(N__26420));
    LocalMux I__5948 (
            .O(N__26435),
            .I(N__26420));
    InMux I__5947 (
            .O(N__26434),
            .I(N__26416));
    InMux I__5946 (
            .O(N__26433),
            .I(N__26413));
    Span12Mux_h I__5945 (
            .O(N__26430),
            .I(N__26410));
    Span4Mux_v I__5944 (
            .O(N__26427),
            .I(N__26405));
    Span4Mux_h I__5943 (
            .O(N__26420),
            .I(N__26405));
    InMux I__5942 (
            .O(N__26419),
            .I(N__26402));
    LocalMux I__5941 (
            .O(N__26416),
            .I(N__26399));
    LocalMux I__5940 (
            .O(N__26413),
            .I(N__26396));
    Odrv12 I__5939 (
            .O(N__26410),
            .I(M_this_sprites_address_qZ0Z_8));
    Odrv4 I__5938 (
            .O(N__26405),
            .I(M_this_sprites_address_qZ0Z_8));
    LocalMux I__5937 (
            .O(N__26402),
            .I(M_this_sprites_address_qZ0Z_8));
    Odrv4 I__5936 (
            .O(N__26399),
            .I(M_this_sprites_address_qZ0Z_8));
    Odrv4 I__5935 (
            .O(N__26396),
            .I(M_this_sprites_address_qZ0Z_8));
    CascadeMux I__5934 (
            .O(N__26385),
            .I(N__26380));
    InMux I__5933 (
            .O(N__26384),
            .I(N__26370));
    InMux I__5932 (
            .O(N__26383),
            .I(N__26365));
    InMux I__5931 (
            .O(N__26380),
            .I(N__26365));
    InMux I__5930 (
            .O(N__26379),
            .I(N__26362));
    InMux I__5929 (
            .O(N__26378),
            .I(N__26359));
    InMux I__5928 (
            .O(N__26377),
            .I(N__26353));
    InMux I__5927 (
            .O(N__26376),
            .I(N__26349));
    InMux I__5926 (
            .O(N__26375),
            .I(N__26346));
    InMux I__5925 (
            .O(N__26374),
            .I(N__26343));
    InMux I__5924 (
            .O(N__26373),
            .I(N__26340));
    LocalMux I__5923 (
            .O(N__26370),
            .I(N__26335));
    LocalMux I__5922 (
            .O(N__26365),
            .I(N__26335));
    LocalMux I__5921 (
            .O(N__26362),
            .I(N__26330));
    LocalMux I__5920 (
            .O(N__26359),
            .I(N__26330));
    InMux I__5919 (
            .O(N__26358),
            .I(N__26325));
    InMux I__5918 (
            .O(N__26357),
            .I(N__26325));
    InMux I__5917 (
            .O(N__26356),
            .I(N__26322));
    LocalMux I__5916 (
            .O(N__26353),
            .I(N__26319));
    InMux I__5915 (
            .O(N__26352),
            .I(N__26315));
    LocalMux I__5914 (
            .O(N__26349),
            .I(N__26310));
    LocalMux I__5913 (
            .O(N__26346),
            .I(N__26310));
    LocalMux I__5912 (
            .O(N__26343),
            .I(N__26307));
    LocalMux I__5911 (
            .O(N__26340),
            .I(N__26298));
    Span4Mux_v I__5910 (
            .O(N__26335),
            .I(N__26298));
    Span4Mux_h I__5909 (
            .O(N__26330),
            .I(N__26298));
    LocalMux I__5908 (
            .O(N__26325),
            .I(N__26298));
    LocalMux I__5907 (
            .O(N__26322),
            .I(N__26293));
    Span4Mux_h I__5906 (
            .O(N__26319),
            .I(N__26293));
    InMux I__5905 (
            .O(N__26318),
            .I(N__26287));
    LocalMux I__5904 (
            .O(N__26315),
            .I(N__26284));
    Span4Mux_h I__5903 (
            .O(N__26310),
            .I(N__26281));
    Span4Mux_h I__5902 (
            .O(N__26307),
            .I(N__26276));
    Span4Mux_h I__5901 (
            .O(N__26298),
            .I(N__26276));
    Span4Mux_h I__5900 (
            .O(N__26293),
            .I(N__26273));
    InMux I__5899 (
            .O(N__26292),
            .I(N__26268));
    InMux I__5898 (
            .O(N__26291),
            .I(N__26268));
    InMux I__5897 (
            .O(N__26290),
            .I(N__26265));
    LocalMux I__5896 (
            .O(N__26287),
            .I(M_this_state_qZ0Z_1));
    Odrv12 I__5895 (
            .O(N__26284),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__5894 (
            .O(N__26281),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__5893 (
            .O(N__26276),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__5892 (
            .O(N__26273),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__5891 (
            .O(N__26268),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__5890 (
            .O(N__26265),
            .I(M_this_state_qZ0Z_1));
    InMux I__5889 (
            .O(N__26250),
            .I(N__26247));
    LocalMux I__5888 (
            .O(N__26247),
            .I(N__26244));
    Span4Mux_v I__5887 (
            .O(N__26244),
            .I(N__26241));
    Odrv4 I__5886 (
            .O(N__26241),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1 ));
    CascadeMux I__5885 (
            .O(N__26238),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_1_cascade_ ));
    InMux I__5884 (
            .O(N__26235),
            .I(N__26232));
    LocalMux I__5883 (
            .O(N__26232),
            .I(N__26229));
    Span4Mux_h I__5882 (
            .O(N__26229),
            .I(N__26226));
    Odrv4 I__5881 (
            .O(N__26226),
            .I(un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0));
    CascadeMux I__5880 (
            .O(N__26223),
            .I(N__26219));
    CascadeMux I__5879 (
            .O(N__26222),
            .I(N__26216));
    InMux I__5878 (
            .O(N__26219),
            .I(N__26211));
    InMux I__5877 (
            .O(N__26216),
            .I(N__26208));
    CascadeMux I__5876 (
            .O(N__26215),
            .I(N__26205));
    CascadeMux I__5875 (
            .O(N__26214),
            .I(N__26202));
    LocalMux I__5874 (
            .O(N__26211),
            .I(N__26191));
    LocalMux I__5873 (
            .O(N__26208),
            .I(N__26191));
    InMux I__5872 (
            .O(N__26205),
            .I(N__26188));
    InMux I__5871 (
            .O(N__26202),
            .I(N__26185));
    CascadeMux I__5870 (
            .O(N__26201),
            .I(N__26182));
    CascadeMux I__5869 (
            .O(N__26200),
            .I(N__26179));
    CascadeMux I__5868 (
            .O(N__26199),
            .I(N__26173));
    CascadeMux I__5867 (
            .O(N__26198),
            .I(N__26170));
    CascadeMux I__5866 (
            .O(N__26197),
            .I(N__26167));
    CascadeMux I__5865 (
            .O(N__26196),
            .I(N__26164));
    Span4Mux_v I__5864 (
            .O(N__26191),
            .I(N__26157));
    LocalMux I__5863 (
            .O(N__26188),
            .I(N__26157));
    LocalMux I__5862 (
            .O(N__26185),
            .I(N__26157));
    InMux I__5861 (
            .O(N__26182),
            .I(N__26154));
    InMux I__5860 (
            .O(N__26179),
            .I(N__26151));
    CascadeMux I__5859 (
            .O(N__26178),
            .I(N__26148));
    CascadeMux I__5858 (
            .O(N__26177),
            .I(N__26144));
    CascadeMux I__5857 (
            .O(N__26176),
            .I(N__26141));
    InMux I__5856 (
            .O(N__26173),
            .I(N__26135));
    InMux I__5855 (
            .O(N__26170),
            .I(N__26132));
    InMux I__5854 (
            .O(N__26167),
            .I(N__26129));
    InMux I__5853 (
            .O(N__26164),
            .I(N__26126));
    Span4Mux_v I__5852 (
            .O(N__26157),
            .I(N__26119));
    LocalMux I__5851 (
            .O(N__26154),
            .I(N__26119));
    LocalMux I__5850 (
            .O(N__26151),
            .I(N__26119));
    InMux I__5849 (
            .O(N__26148),
            .I(N__26116));
    CascadeMux I__5848 (
            .O(N__26147),
            .I(N__26113));
    InMux I__5847 (
            .O(N__26144),
            .I(N__26110));
    InMux I__5846 (
            .O(N__26141),
            .I(N__26107));
    CascadeMux I__5845 (
            .O(N__26140),
            .I(N__26104));
    CascadeMux I__5844 (
            .O(N__26139),
            .I(N__26101));
    InMux I__5843 (
            .O(N__26138),
            .I(N__26098));
    LocalMux I__5842 (
            .O(N__26135),
            .I(N__26090));
    LocalMux I__5841 (
            .O(N__26132),
            .I(N__26090));
    LocalMux I__5840 (
            .O(N__26129),
            .I(N__26090));
    LocalMux I__5839 (
            .O(N__26126),
            .I(N__26087));
    Span4Mux_v I__5838 (
            .O(N__26119),
            .I(N__26082));
    LocalMux I__5837 (
            .O(N__26116),
            .I(N__26082));
    InMux I__5836 (
            .O(N__26113),
            .I(N__26079));
    LocalMux I__5835 (
            .O(N__26110),
            .I(N__26074));
    LocalMux I__5834 (
            .O(N__26107),
            .I(N__26074));
    InMux I__5833 (
            .O(N__26104),
            .I(N__26071));
    InMux I__5832 (
            .O(N__26101),
            .I(N__26068));
    LocalMux I__5831 (
            .O(N__26098),
            .I(N__26065));
    InMux I__5830 (
            .O(N__26097),
            .I(N__26062));
    Span12Mux_v I__5829 (
            .O(N__26090),
            .I(N__26057));
    Span12Mux_s9_v I__5828 (
            .O(N__26087),
            .I(N__26057));
    Span4Mux_v I__5827 (
            .O(N__26082),
            .I(N__26052));
    LocalMux I__5826 (
            .O(N__26079),
            .I(N__26052));
    Span4Mux_v I__5825 (
            .O(N__26074),
            .I(N__26045));
    LocalMux I__5824 (
            .O(N__26071),
            .I(N__26045));
    LocalMux I__5823 (
            .O(N__26068),
            .I(N__26045));
    Span4Mux_v I__5822 (
            .O(N__26065),
            .I(N__26039));
    LocalMux I__5821 (
            .O(N__26062),
            .I(N__26039));
    Span12Mux_h I__5820 (
            .O(N__26057),
            .I(N__26036));
    Span4Mux_v I__5819 (
            .O(N__26052),
            .I(N__26031));
    Span4Mux_v I__5818 (
            .O(N__26045),
            .I(N__26031));
    InMux I__5817 (
            .O(N__26044),
            .I(N__26028));
    Span4Mux_h I__5816 (
            .O(N__26039),
            .I(N__26025));
    Odrv12 I__5815 (
            .O(N__26036),
            .I(M_this_sprites_address_qZ0Z_1));
    Odrv4 I__5814 (
            .O(N__26031),
            .I(M_this_sprites_address_qZ0Z_1));
    LocalMux I__5813 (
            .O(N__26028),
            .I(M_this_sprites_address_qZ0Z_1));
    Odrv4 I__5812 (
            .O(N__26025),
            .I(M_this_sprites_address_qZ0Z_1));
    InMux I__5811 (
            .O(N__26016),
            .I(bfn_21_19_0_));
    InMux I__5810 (
            .O(N__26013),
            .I(N__26007));
    InMux I__5809 (
            .O(N__26012),
            .I(N__26000));
    InMux I__5808 (
            .O(N__26011),
            .I(N__26000));
    InMux I__5807 (
            .O(N__26010),
            .I(N__26000));
    LocalMux I__5806 (
            .O(N__26007),
            .I(\this_ppu.vscroll8 ));
    LocalMux I__5805 (
            .O(N__26000),
            .I(\this_ppu.vscroll8 ));
    CascadeMux I__5804 (
            .O(N__25995),
            .I(N__25991));
    InMux I__5803 (
            .O(N__25994),
            .I(N__25988));
    InMux I__5802 (
            .O(N__25991),
            .I(N__25985));
    LocalMux I__5801 (
            .O(N__25988),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    LocalMux I__5800 (
            .O(N__25985),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    InMux I__5799 (
            .O(N__25980),
            .I(N__25977));
    LocalMux I__5798 (
            .O(N__25977),
            .I(N__25974));
    Span4Mux_v I__5797 (
            .O(N__25974),
            .I(N__25971));
    Span4Mux_h I__5796 (
            .O(N__25971),
            .I(N__25968));
    Odrv4 I__5795 (
            .O(N__25968),
            .I(N_48_0));
    InMux I__5794 (
            .O(N__25965),
            .I(N__25962));
    LocalMux I__5793 (
            .O(N__25962),
            .I(N__25959));
    Span4Mux_h I__5792 (
            .O(N__25959),
            .I(N__25956));
    Odrv4 I__5791 (
            .O(N__25956),
            .I(M_this_oam_ram_write_data_28));
    CascadeMux I__5790 (
            .O(N__25953),
            .I(N__25948));
    InMux I__5789 (
            .O(N__25952),
            .I(N__25944));
    InMux I__5788 (
            .O(N__25951),
            .I(N__25937));
    InMux I__5787 (
            .O(N__25948),
            .I(N__25937));
    InMux I__5786 (
            .O(N__25947),
            .I(N__25937));
    LocalMux I__5785 (
            .O(N__25944),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    LocalMux I__5784 (
            .O(N__25937),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    CascadeMux I__5783 (
            .O(N__25932),
            .I(N__25927));
    InMux I__5782 (
            .O(N__25931),
            .I(N__25922));
    InMux I__5781 (
            .O(N__25930),
            .I(N__25918));
    InMux I__5780 (
            .O(N__25927),
            .I(N__25915));
    CascadeMux I__5779 (
            .O(N__25926),
            .I(N__25912));
    InMux I__5778 (
            .O(N__25925),
            .I(N__25907));
    LocalMux I__5777 (
            .O(N__25922),
            .I(N__25904));
    InMux I__5776 (
            .O(N__25921),
            .I(N__25901));
    LocalMux I__5775 (
            .O(N__25918),
            .I(N__25896));
    LocalMux I__5774 (
            .O(N__25915),
            .I(N__25896));
    InMux I__5773 (
            .O(N__25912),
            .I(N__25891));
    InMux I__5772 (
            .O(N__25911),
            .I(N__25891));
    InMux I__5771 (
            .O(N__25910),
            .I(N__25888));
    LocalMux I__5770 (
            .O(N__25907),
            .I(N__25885));
    Span4Mux_v I__5769 (
            .O(N__25904),
            .I(N__25880));
    LocalMux I__5768 (
            .O(N__25901),
            .I(N__25880));
    Span4Mux_v I__5767 (
            .O(N__25896),
            .I(N__25877));
    LocalMux I__5766 (
            .O(N__25891),
            .I(N__25874));
    LocalMux I__5765 (
            .O(N__25888),
            .I(N__25871));
    Span4Mux_h I__5764 (
            .O(N__25885),
            .I(N__25866));
    Span4Mux_h I__5763 (
            .O(N__25880),
            .I(N__25866));
    Odrv4 I__5762 (
            .O(N__25877),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    Odrv4 I__5761 (
            .O(N__25874),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    Odrv12 I__5760 (
            .O(N__25871),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    Odrv4 I__5759 (
            .O(N__25866),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    InMux I__5758 (
            .O(N__25857),
            .I(N__25853));
    InMux I__5757 (
            .O(N__25856),
            .I(N__25850));
    LocalMux I__5756 (
            .O(N__25853),
            .I(N__25847));
    LocalMux I__5755 (
            .O(N__25850),
            .I(N__25843));
    Span12Mux_h I__5754 (
            .O(N__25847),
            .I(N__25840));
    InMux I__5753 (
            .O(N__25846),
            .I(N__25837));
    Odrv12 I__5752 (
            .O(N__25843),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_7 ));
    Odrv12 I__5751 (
            .O(N__25840),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_7 ));
    LocalMux I__5750 (
            .O(N__25837),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_7 ));
    InMux I__5749 (
            .O(N__25830),
            .I(N__25827));
    LocalMux I__5748 (
            .O(N__25827),
            .I(\this_ppu.N_148 ));
    CascadeMux I__5747 (
            .O(N__25824),
            .I(N__25821));
    InMux I__5746 (
            .O(N__25821),
            .I(N__25818));
    LocalMux I__5745 (
            .O(N__25818),
            .I(N__25815));
    Odrv4 I__5744 (
            .O(N__25815),
            .I(M_this_data_tmp_qZ0Z_20));
    CascadeMux I__5743 (
            .O(N__25812),
            .I(N__25809));
    InMux I__5742 (
            .O(N__25809),
            .I(N__25804));
    CascadeMux I__5741 (
            .O(N__25808),
            .I(N__25801));
    CascadeMux I__5740 (
            .O(N__25807),
            .I(N__25795));
    LocalMux I__5739 (
            .O(N__25804),
            .I(N__25791));
    InMux I__5738 (
            .O(N__25801),
            .I(N__25788));
    CascadeMux I__5737 (
            .O(N__25800),
            .I(N__25785));
    CascadeMux I__5736 (
            .O(N__25799),
            .I(N__25781));
    CascadeMux I__5735 (
            .O(N__25798),
            .I(N__25777));
    InMux I__5734 (
            .O(N__25795),
            .I(N__25772));
    CascadeMux I__5733 (
            .O(N__25794),
            .I(N__25769));
    Span4Mux_s2_v I__5732 (
            .O(N__25791),
            .I(N__25764));
    LocalMux I__5731 (
            .O(N__25788),
            .I(N__25764));
    InMux I__5730 (
            .O(N__25785),
            .I(N__25761));
    CascadeMux I__5729 (
            .O(N__25784),
            .I(N__25758));
    InMux I__5728 (
            .O(N__25781),
            .I(N__25754));
    CascadeMux I__5727 (
            .O(N__25780),
            .I(N__25751));
    InMux I__5726 (
            .O(N__25777),
            .I(N__25748));
    CascadeMux I__5725 (
            .O(N__25776),
            .I(N__25745));
    CascadeMux I__5724 (
            .O(N__25775),
            .I(N__25742));
    LocalMux I__5723 (
            .O(N__25772),
            .I(N__25737));
    InMux I__5722 (
            .O(N__25769),
            .I(N__25734));
    Span4Mux_v I__5721 (
            .O(N__25764),
            .I(N__25729));
    LocalMux I__5720 (
            .O(N__25761),
            .I(N__25729));
    InMux I__5719 (
            .O(N__25758),
            .I(N__25726));
    CascadeMux I__5718 (
            .O(N__25757),
            .I(N__25723));
    LocalMux I__5717 (
            .O(N__25754),
            .I(N__25719));
    InMux I__5716 (
            .O(N__25751),
            .I(N__25716));
    LocalMux I__5715 (
            .O(N__25748),
            .I(N__25712));
    InMux I__5714 (
            .O(N__25745),
            .I(N__25709));
    InMux I__5713 (
            .O(N__25742),
            .I(N__25706));
    CascadeMux I__5712 (
            .O(N__25741),
            .I(N__25703));
    CascadeMux I__5711 (
            .O(N__25740),
            .I(N__25700));
    Span4Mux_h I__5710 (
            .O(N__25737),
            .I(N__25697));
    LocalMux I__5709 (
            .O(N__25734),
            .I(N__25694));
    Span4Mux_h I__5708 (
            .O(N__25729),
            .I(N__25689));
    LocalMux I__5707 (
            .O(N__25726),
            .I(N__25689));
    InMux I__5706 (
            .O(N__25723),
            .I(N__25686));
    CascadeMux I__5705 (
            .O(N__25722),
            .I(N__25683));
    Span4Mux_v I__5704 (
            .O(N__25719),
            .I(N__25678));
    LocalMux I__5703 (
            .O(N__25716),
            .I(N__25678));
    CascadeMux I__5702 (
            .O(N__25715),
            .I(N__25675));
    Span4Mux_v I__5701 (
            .O(N__25712),
            .I(N__25670));
    LocalMux I__5700 (
            .O(N__25709),
            .I(N__25670));
    LocalMux I__5699 (
            .O(N__25706),
            .I(N__25667));
    InMux I__5698 (
            .O(N__25703),
            .I(N__25664));
    InMux I__5697 (
            .O(N__25700),
            .I(N__25661));
    Span4Mux_h I__5696 (
            .O(N__25697),
            .I(N__25658));
    Span4Mux_h I__5695 (
            .O(N__25694),
            .I(N__25655));
    Span4Mux_v I__5694 (
            .O(N__25689),
            .I(N__25650));
    LocalMux I__5693 (
            .O(N__25686),
            .I(N__25650));
    InMux I__5692 (
            .O(N__25683),
            .I(N__25647));
    Span4Mux_h I__5691 (
            .O(N__25678),
            .I(N__25644));
    InMux I__5690 (
            .O(N__25675),
            .I(N__25641));
    Span4Mux_v I__5689 (
            .O(N__25670),
            .I(N__25632));
    Span4Mux_v I__5688 (
            .O(N__25667),
            .I(N__25632));
    LocalMux I__5687 (
            .O(N__25664),
            .I(N__25632));
    LocalMux I__5686 (
            .O(N__25661),
            .I(N__25632));
    Span4Mux_v I__5685 (
            .O(N__25658),
            .I(N__25627));
    Span4Mux_h I__5684 (
            .O(N__25655),
            .I(N__25627));
    Span4Mux_v I__5683 (
            .O(N__25650),
            .I(N__25622));
    LocalMux I__5682 (
            .O(N__25647),
            .I(N__25622));
    Span4Mux_v I__5681 (
            .O(N__25644),
            .I(N__25619));
    LocalMux I__5680 (
            .O(N__25641),
            .I(N__25616));
    Span4Mux_v I__5679 (
            .O(N__25632),
            .I(N__25613));
    Span4Mux_h I__5678 (
            .O(N__25627),
            .I(N__25608));
    Span4Mux_h I__5677 (
            .O(N__25622),
            .I(N__25608));
    Sp12to4 I__5676 (
            .O(N__25619),
            .I(N__25605));
    Span12Mux_s11_h I__5675 (
            .O(N__25616),
            .I(N__25602));
    Span4Mux_h I__5674 (
            .O(N__25613),
            .I(N__25597));
    Span4Mux_h I__5673 (
            .O(N__25608),
            .I(N__25597));
    Odrv12 I__5672 (
            .O(N__25605),
            .I(M_this_ppu_sprites_addr_1));
    Odrv12 I__5671 (
            .O(N__25602),
            .I(M_this_ppu_sprites_addr_1));
    Odrv4 I__5670 (
            .O(N__25597),
            .I(M_this_ppu_sprites_addr_1));
    CascadeMux I__5669 (
            .O(N__25590),
            .I(N__25587));
    InMux I__5668 (
            .O(N__25587),
            .I(N__25584));
    LocalMux I__5667 (
            .O(N__25584),
            .I(N__25581));
    Span12Mux_v I__5666 (
            .O(N__25581),
            .I(N__25577));
    CascadeMux I__5665 (
            .O(N__25580),
            .I(N__25574));
    Span12Mux_h I__5664 (
            .O(N__25577),
            .I(N__25564));
    InMux I__5663 (
            .O(N__25574),
            .I(N__25553));
    InMux I__5662 (
            .O(N__25573),
            .I(N__25553));
    InMux I__5661 (
            .O(N__25572),
            .I(N__25553));
    InMux I__5660 (
            .O(N__25571),
            .I(N__25553));
    InMux I__5659 (
            .O(N__25570),
            .I(N__25553));
    InMux I__5658 (
            .O(N__25569),
            .I(N__25550));
    InMux I__5657 (
            .O(N__25568),
            .I(N__25547));
    InMux I__5656 (
            .O(N__25567),
            .I(N__25544));
    Odrv12 I__5655 (
            .O(N__25564),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__5654 (
            .O(N__25553),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__5653 (
            .O(N__25550),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__5652 (
            .O(N__25547),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__5651 (
            .O(N__25544),
            .I(M_this_ppu_vram_addr_0));
    CascadeMux I__5650 (
            .O(N__25533),
            .I(N__25530));
    InMux I__5649 (
            .O(N__25530),
            .I(N__25527));
    LocalMux I__5648 (
            .O(N__25527),
            .I(N__25524));
    Span4Mux_h I__5647 (
            .O(N__25524),
            .I(N__25521));
    Span4Mux_h I__5646 (
            .O(N__25521),
            .I(N__25514));
    InMux I__5645 (
            .O(N__25520),
            .I(N__25509));
    InMux I__5644 (
            .O(N__25519),
            .I(N__25509));
    InMux I__5643 (
            .O(N__25518),
            .I(N__25506));
    InMux I__5642 (
            .O(N__25517),
            .I(N__25503));
    Span4Mux_h I__5641 (
            .O(N__25514),
            .I(N__25498));
    LocalMux I__5640 (
            .O(N__25509),
            .I(N__25491));
    LocalMux I__5639 (
            .O(N__25506),
            .I(N__25491));
    LocalMux I__5638 (
            .O(N__25503),
            .I(N__25491));
    InMux I__5637 (
            .O(N__25502),
            .I(N__25488));
    InMux I__5636 (
            .O(N__25501),
            .I(N__25485));
    Odrv4 I__5635 (
            .O(N__25498),
            .I(M_this_ppu_vram_addr_1));
    Odrv4 I__5634 (
            .O(N__25491),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__5633 (
            .O(N__25488),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__5632 (
            .O(N__25485),
            .I(M_this_ppu_vram_addr_1));
    CascadeMux I__5631 (
            .O(N__25476),
            .I(N__25473));
    InMux I__5630 (
            .O(N__25473),
            .I(N__25470));
    LocalMux I__5629 (
            .O(N__25470),
            .I(N__25465));
    InMux I__5628 (
            .O(N__25469),
            .I(N__25455));
    InMux I__5627 (
            .O(N__25468),
            .I(N__25455));
    Span12Mux_h I__5626 (
            .O(N__25465),
            .I(N__25452));
    InMux I__5625 (
            .O(N__25464),
            .I(N__25449));
    InMux I__5624 (
            .O(N__25463),
            .I(N__25444));
    InMux I__5623 (
            .O(N__25462),
            .I(N__25444));
    InMux I__5622 (
            .O(N__25461),
            .I(N__25441));
    InMux I__5621 (
            .O(N__25460),
            .I(N__25438));
    LocalMux I__5620 (
            .O(N__25455),
            .I(M_this_ppu_vram_addr_2));
    Odrv12 I__5619 (
            .O(N__25452),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__5618 (
            .O(N__25449),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__5617 (
            .O(N__25444),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__5616 (
            .O(N__25441),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__5615 (
            .O(N__25438),
            .I(M_this_ppu_vram_addr_2));
    CascadeMux I__5614 (
            .O(N__25425),
            .I(N__25422));
    InMux I__5613 (
            .O(N__25422),
            .I(N__25419));
    LocalMux I__5612 (
            .O(N__25419),
            .I(M_this_oam_ram_read_data_i_11));
    CascadeMux I__5611 (
            .O(N__25416),
            .I(N__25413));
    CascadeBuf I__5610 (
            .O(N__25413),
            .I(N__25409));
    CascadeMux I__5609 (
            .O(N__25412),
            .I(N__25406));
    CascadeMux I__5608 (
            .O(N__25409),
            .I(N__25403));
    InMux I__5607 (
            .O(N__25406),
            .I(N__25400));
    InMux I__5606 (
            .O(N__25403),
            .I(N__25397));
    LocalMux I__5605 (
            .O(N__25400),
            .I(N__25394));
    LocalMux I__5604 (
            .O(N__25397),
            .I(N__25391));
    Span4Mux_h I__5603 (
            .O(N__25394),
            .I(N__25388));
    Span4Mux_h I__5602 (
            .O(N__25391),
            .I(N__25385));
    Span4Mux_h I__5601 (
            .O(N__25388),
            .I(N__25378));
    Sp12to4 I__5600 (
            .O(N__25385),
            .I(N__25375));
    InMux I__5599 (
            .O(N__25384),
            .I(N__25370));
    InMux I__5598 (
            .O(N__25383),
            .I(N__25370));
    InMux I__5597 (
            .O(N__25382),
            .I(N__25367));
    InMux I__5596 (
            .O(N__25381),
            .I(N__25364));
    Span4Mux_h I__5595 (
            .O(N__25378),
            .I(N__25361));
    Span12Mux_v I__5594 (
            .O(N__25375),
            .I(N__25358));
    LocalMux I__5593 (
            .O(N__25370),
            .I(M_this_ppu_map_addr_0));
    LocalMux I__5592 (
            .O(N__25367),
            .I(M_this_ppu_map_addr_0));
    LocalMux I__5591 (
            .O(N__25364),
            .I(M_this_ppu_map_addr_0));
    Odrv4 I__5590 (
            .O(N__25361),
            .I(M_this_ppu_map_addr_0));
    Odrv12 I__5589 (
            .O(N__25358),
            .I(M_this_ppu_map_addr_0));
    CascadeMux I__5588 (
            .O(N__25347),
            .I(N__25344));
    InMux I__5587 (
            .O(N__25344),
            .I(N__25341));
    LocalMux I__5586 (
            .O(N__25341),
            .I(N__25338));
    Odrv4 I__5585 (
            .O(N__25338),
            .I(\this_ppu.un1_M_haddress_q_2_4 ));
    CascadeMux I__5584 (
            .O(N__25335),
            .I(N__25331));
    CascadeMux I__5583 (
            .O(N__25334),
            .I(N__25328));
    CascadeBuf I__5582 (
            .O(N__25331),
            .I(N__25325));
    InMux I__5581 (
            .O(N__25328),
            .I(N__25322));
    CascadeMux I__5580 (
            .O(N__25325),
            .I(N__25319));
    LocalMux I__5579 (
            .O(N__25322),
            .I(N__25316));
    InMux I__5578 (
            .O(N__25319),
            .I(N__25313));
    Sp12to4 I__5577 (
            .O(N__25316),
            .I(N__25309));
    LocalMux I__5576 (
            .O(N__25313),
            .I(N__25306));
    CascadeMux I__5575 (
            .O(N__25312),
            .I(N__25303));
    Span12Mux_v I__5574 (
            .O(N__25309),
            .I(N__25298));
    Span12Mux_s8_v I__5573 (
            .O(N__25306),
            .I(N__25295));
    InMux I__5572 (
            .O(N__25303),
            .I(N__25292));
    InMux I__5571 (
            .O(N__25302),
            .I(N__25289));
    InMux I__5570 (
            .O(N__25301),
            .I(N__25286));
    Span12Mux_h I__5569 (
            .O(N__25298),
            .I(N__25281));
    Span12Mux_h I__5568 (
            .O(N__25295),
            .I(N__25281));
    LocalMux I__5567 (
            .O(N__25292),
            .I(M_this_ppu_map_addr_1));
    LocalMux I__5566 (
            .O(N__25289),
            .I(M_this_ppu_map_addr_1));
    LocalMux I__5565 (
            .O(N__25286),
            .I(M_this_ppu_map_addr_1));
    Odrv12 I__5564 (
            .O(N__25281),
            .I(M_this_ppu_map_addr_1));
    CascadeMux I__5563 (
            .O(N__25272),
            .I(N__25269));
    CascadeBuf I__5562 (
            .O(N__25269),
            .I(N__25265));
    CascadeMux I__5561 (
            .O(N__25268),
            .I(N__25262));
    CascadeMux I__5560 (
            .O(N__25265),
            .I(N__25259));
    InMux I__5559 (
            .O(N__25262),
            .I(N__25253));
    InMux I__5558 (
            .O(N__25259),
            .I(N__25250));
    CascadeMux I__5557 (
            .O(N__25258),
            .I(N__25247));
    CascadeMux I__5556 (
            .O(N__25257),
            .I(N__25244));
    InMux I__5555 (
            .O(N__25256),
            .I(N__25240));
    LocalMux I__5554 (
            .O(N__25253),
            .I(N__25237));
    LocalMux I__5553 (
            .O(N__25250),
            .I(N__25234));
    InMux I__5552 (
            .O(N__25247),
            .I(N__25227));
    InMux I__5551 (
            .O(N__25244),
            .I(N__25227));
    InMux I__5550 (
            .O(N__25243),
            .I(N__25227));
    LocalMux I__5549 (
            .O(N__25240),
            .I(N__25222));
    Span12Mux_h I__5548 (
            .O(N__25237),
            .I(N__25222));
    Span12Mux_h I__5547 (
            .O(N__25234),
            .I(N__25219));
    LocalMux I__5546 (
            .O(N__25227),
            .I(M_this_ppu_map_addr_2));
    Odrv12 I__5545 (
            .O(N__25222),
            .I(M_this_ppu_map_addr_2));
    Odrv12 I__5544 (
            .O(N__25219),
            .I(M_this_ppu_map_addr_2));
    CascadeMux I__5543 (
            .O(N__25212),
            .I(N__25209));
    CascadeBuf I__5542 (
            .O(N__25209),
            .I(N__25206));
    CascadeMux I__5541 (
            .O(N__25206),
            .I(N__25203));
    InMux I__5540 (
            .O(N__25203),
            .I(N__25199));
    CascadeMux I__5539 (
            .O(N__25202),
            .I(N__25196));
    LocalMux I__5538 (
            .O(N__25199),
            .I(N__25193));
    InMux I__5537 (
            .O(N__25196),
            .I(N__25189));
    Span4Mux_v I__5536 (
            .O(N__25193),
            .I(N__25186));
    InMux I__5535 (
            .O(N__25192),
            .I(N__25181));
    LocalMux I__5534 (
            .O(N__25189),
            .I(N__25178));
    Sp12to4 I__5533 (
            .O(N__25186),
            .I(N__25175));
    InMux I__5532 (
            .O(N__25185),
            .I(N__25170));
    InMux I__5531 (
            .O(N__25184),
            .I(N__25170));
    LocalMux I__5530 (
            .O(N__25181),
            .I(N__25165));
    Span12Mux_s11_h I__5529 (
            .O(N__25178),
            .I(N__25165));
    Span12Mux_h I__5528 (
            .O(N__25175),
            .I(N__25162));
    LocalMux I__5527 (
            .O(N__25170),
            .I(M_this_ppu_map_addr_3));
    Odrv12 I__5526 (
            .O(N__25165),
            .I(M_this_ppu_map_addr_3));
    Odrv12 I__5525 (
            .O(N__25162),
            .I(M_this_ppu_map_addr_3));
    CascadeMux I__5524 (
            .O(N__25155),
            .I(N__25152));
    CascadeBuf I__5523 (
            .O(N__25152),
            .I(N__25149));
    CascadeMux I__5522 (
            .O(N__25149),
            .I(N__25146));
    InMux I__5521 (
            .O(N__25146),
            .I(N__25143));
    LocalMux I__5520 (
            .O(N__25143),
            .I(N__25140));
    Span4Mux_v I__5519 (
            .O(N__25140),
            .I(N__25136));
    InMux I__5518 (
            .O(N__25139),
            .I(N__25132));
    Sp12to4 I__5517 (
            .O(N__25136),
            .I(N__25129));
    InMux I__5516 (
            .O(N__25135),
            .I(N__25126));
    LocalMux I__5515 (
            .O(N__25132),
            .I(N__25123));
    Span12Mux_h I__5514 (
            .O(N__25129),
            .I(N__25120));
    LocalMux I__5513 (
            .O(N__25126),
            .I(M_this_ppu_map_addr_4));
    Odrv4 I__5512 (
            .O(N__25123),
            .I(M_this_ppu_map_addr_4));
    Odrv12 I__5511 (
            .O(N__25120),
            .I(M_this_ppu_map_addr_4));
    CascadeMux I__5510 (
            .O(N__25113),
            .I(N__25110));
    InMux I__5509 (
            .O(N__25110),
            .I(N__25107));
    LocalMux I__5508 (
            .O(N__25107),
            .I(\this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ));
    InMux I__5507 (
            .O(N__25104),
            .I(\this_ppu.un2_hscroll_cry_0 ));
    InMux I__5506 (
            .O(N__25101),
            .I(\this_ppu.un2_hscroll_cry_1 ));
    InMux I__5505 (
            .O(N__25098),
            .I(N__25095));
    LocalMux I__5504 (
            .O(N__25095),
            .I(\this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0 ));
    CEMux I__5503 (
            .O(N__25092),
            .I(N__25089));
    LocalMux I__5502 (
            .O(N__25089),
            .I(N__25085));
    CEMux I__5501 (
            .O(N__25088),
            .I(N__25082));
    Span4Mux_h I__5500 (
            .O(N__25085),
            .I(N__25077));
    LocalMux I__5499 (
            .O(N__25082),
            .I(N__25077));
    Span4Mux_v I__5498 (
            .O(N__25077),
            .I(N__25074));
    Span4Mux_h I__5497 (
            .O(N__25074),
            .I(N__25071));
    Odrv4 I__5496 (
            .O(N__25071),
            .I(\this_sprites_ram.mem_WE_12 ));
    InMux I__5495 (
            .O(N__25068),
            .I(N__25065));
    LocalMux I__5494 (
            .O(N__25065),
            .I(N__25062));
    Span4Mux_h I__5493 (
            .O(N__25062),
            .I(N__25059));
    Span4Mux_v I__5492 (
            .O(N__25059),
            .I(N__25056));
    Span4Mux_v I__5491 (
            .O(N__25056),
            .I(N__25053));
    Odrv4 I__5490 (
            .O(N__25053),
            .I(\this_sprites_ram.mem_out_bus6_2 ));
    InMux I__5489 (
            .O(N__25050),
            .I(N__25047));
    LocalMux I__5488 (
            .O(N__25047),
            .I(N__25044));
    Span4Mux_h I__5487 (
            .O(N__25044),
            .I(N__25041));
    Odrv4 I__5486 (
            .O(N__25041),
            .I(\this_sprites_ram.mem_out_bus2_2 ));
    InMux I__5485 (
            .O(N__25038),
            .I(N__25035));
    LocalMux I__5484 (
            .O(N__25035),
            .I(N__25032));
    Odrv12 I__5483 (
            .O(N__25032),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ));
    CascadeMux I__5482 (
            .O(N__25029),
            .I(N__25026));
    InMux I__5481 (
            .O(N__25026),
            .I(N__25023));
    LocalMux I__5480 (
            .O(N__25023),
            .I(M_this_oam_ram_read_data_i_9));
    InMux I__5479 (
            .O(N__25020),
            .I(N__25017));
    LocalMux I__5478 (
            .O(N__25017),
            .I(\this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0 ));
    CascadeMux I__5477 (
            .O(N__25014),
            .I(N__25009));
    CascadeMux I__5476 (
            .O(N__25013),
            .I(N__25006));
    InMux I__5475 (
            .O(N__25012),
            .I(N__24999));
    InMux I__5474 (
            .O(N__25009),
            .I(N__24990));
    InMux I__5473 (
            .O(N__25006),
            .I(N__24990));
    InMux I__5472 (
            .O(N__25005),
            .I(N__24987));
    InMux I__5471 (
            .O(N__25004),
            .I(N__24979));
    InMux I__5470 (
            .O(N__25003),
            .I(N__24979));
    InMux I__5469 (
            .O(N__25002),
            .I(N__24976));
    LocalMux I__5468 (
            .O(N__24999),
            .I(N__24973));
    InMux I__5467 (
            .O(N__24998),
            .I(N__24966));
    InMux I__5466 (
            .O(N__24997),
            .I(N__24966));
    InMux I__5465 (
            .O(N__24996),
            .I(N__24966));
    CascadeMux I__5464 (
            .O(N__24995),
            .I(N__24962));
    LocalMux I__5463 (
            .O(N__24990),
            .I(N__24957));
    LocalMux I__5462 (
            .O(N__24987),
            .I(N__24954));
    InMux I__5461 (
            .O(N__24986),
            .I(N__24949));
    InMux I__5460 (
            .O(N__24985),
            .I(N__24949));
    InMux I__5459 (
            .O(N__24984),
            .I(N__24946));
    LocalMux I__5458 (
            .O(N__24979),
            .I(N__24937));
    LocalMux I__5457 (
            .O(N__24976),
            .I(N__24937));
    Span4Mux_v I__5456 (
            .O(N__24973),
            .I(N__24937));
    LocalMux I__5455 (
            .O(N__24966),
            .I(N__24937));
    CascadeMux I__5454 (
            .O(N__24965),
            .I(N__24934));
    InMux I__5453 (
            .O(N__24962),
            .I(N__24930));
    InMux I__5452 (
            .O(N__24961),
            .I(N__24927));
    InMux I__5451 (
            .O(N__24960),
            .I(N__24924));
    Span4Mux_h I__5450 (
            .O(N__24957),
            .I(N__24919));
    Span4Mux_h I__5449 (
            .O(N__24954),
            .I(N__24919));
    LocalMux I__5448 (
            .O(N__24949),
            .I(N__24916));
    LocalMux I__5447 (
            .O(N__24946),
            .I(N__24911));
    Span4Mux_h I__5446 (
            .O(N__24937),
            .I(N__24911));
    InMux I__5445 (
            .O(N__24934),
            .I(N__24908));
    InMux I__5444 (
            .O(N__24933),
            .I(N__24905));
    LocalMux I__5443 (
            .O(N__24930),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__5442 (
            .O(N__24927),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__5441 (
            .O(N__24924),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__5440 (
            .O(N__24919),
            .I(M_this_state_qZ0Z_2));
    Odrv12 I__5439 (
            .O(N__24916),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__5438 (
            .O(N__24911),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__5437 (
            .O(N__24908),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__5436 (
            .O(N__24905),
            .I(M_this_state_qZ0Z_2));
    CascadeMux I__5435 (
            .O(N__24888),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_10_cascade_ ));
    InMux I__5434 (
            .O(N__24885),
            .I(N__24882));
    LocalMux I__5433 (
            .O(N__24882),
            .I(un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0));
    CascadeMux I__5432 (
            .O(N__24879),
            .I(N__24876));
    InMux I__5431 (
            .O(N__24876),
            .I(N__24871));
    CascadeMux I__5430 (
            .O(N__24875),
            .I(N__24868));
    CascadeMux I__5429 (
            .O(N__24874),
            .I(N__24865));
    LocalMux I__5428 (
            .O(N__24871),
            .I(N__24861));
    InMux I__5427 (
            .O(N__24868),
            .I(N__24858));
    InMux I__5426 (
            .O(N__24865),
            .I(N__24855));
    CascadeMux I__5425 (
            .O(N__24864),
            .I(N__24852));
    Span4Mux_h I__5424 (
            .O(N__24861),
            .I(N__24844));
    LocalMux I__5423 (
            .O(N__24858),
            .I(N__24844));
    LocalMux I__5422 (
            .O(N__24855),
            .I(N__24841));
    InMux I__5421 (
            .O(N__24852),
            .I(N__24838));
    CascadeMux I__5420 (
            .O(N__24851),
            .I(N__24835));
    CascadeMux I__5419 (
            .O(N__24850),
            .I(N__24832));
    CascadeMux I__5418 (
            .O(N__24849),
            .I(N__24827));
    Span4Mux_v I__5417 (
            .O(N__24844),
            .I(N__24818));
    Span4Mux_h I__5416 (
            .O(N__24841),
            .I(N__24818));
    LocalMux I__5415 (
            .O(N__24838),
            .I(N__24818));
    InMux I__5414 (
            .O(N__24835),
            .I(N__24815));
    InMux I__5413 (
            .O(N__24832),
            .I(N__24812));
    CascadeMux I__5412 (
            .O(N__24831),
            .I(N__24808));
    CascadeMux I__5411 (
            .O(N__24830),
            .I(N__24803));
    InMux I__5410 (
            .O(N__24827),
            .I(N__24800));
    CascadeMux I__5409 (
            .O(N__24826),
            .I(N__24797));
    CascadeMux I__5408 (
            .O(N__24825),
            .I(N__24794));
    Span4Mux_v I__5407 (
            .O(N__24818),
            .I(N__24788));
    LocalMux I__5406 (
            .O(N__24815),
            .I(N__24788));
    LocalMux I__5405 (
            .O(N__24812),
            .I(N__24785));
    CascadeMux I__5404 (
            .O(N__24811),
            .I(N__24782));
    InMux I__5403 (
            .O(N__24808),
            .I(N__24779));
    CascadeMux I__5402 (
            .O(N__24807),
            .I(N__24776));
    CascadeMux I__5401 (
            .O(N__24806),
            .I(N__24773));
    InMux I__5400 (
            .O(N__24803),
            .I(N__24770));
    LocalMux I__5399 (
            .O(N__24800),
            .I(N__24767));
    InMux I__5398 (
            .O(N__24797),
            .I(N__24764));
    InMux I__5397 (
            .O(N__24794),
            .I(N__24761));
    CascadeMux I__5396 (
            .O(N__24793),
            .I(N__24758));
    Span4Mux_v I__5395 (
            .O(N__24788),
            .I(N__24753));
    Span4Mux_h I__5394 (
            .O(N__24785),
            .I(N__24753));
    InMux I__5393 (
            .O(N__24782),
            .I(N__24750));
    LocalMux I__5392 (
            .O(N__24779),
            .I(N__24747));
    InMux I__5391 (
            .O(N__24776),
            .I(N__24744));
    InMux I__5390 (
            .O(N__24773),
            .I(N__24741));
    LocalMux I__5389 (
            .O(N__24770),
            .I(N__24737));
    Span4Mux_h I__5388 (
            .O(N__24767),
            .I(N__24732));
    LocalMux I__5387 (
            .O(N__24764),
            .I(N__24732));
    LocalMux I__5386 (
            .O(N__24761),
            .I(N__24729));
    InMux I__5385 (
            .O(N__24758),
            .I(N__24726));
    Span4Mux_v I__5384 (
            .O(N__24753),
            .I(N__24721));
    LocalMux I__5383 (
            .O(N__24750),
            .I(N__24721));
    Span4Mux_v I__5382 (
            .O(N__24747),
            .I(N__24714));
    LocalMux I__5381 (
            .O(N__24744),
            .I(N__24714));
    LocalMux I__5380 (
            .O(N__24741),
            .I(N__24714));
    CascadeMux I__5379 (
            .O(N__24740),
            .I(N__24711));
    Sp12to4 I__5378 (
            .O(N__24737),
            .I(N__24708));
    Span4Mux_v I__5377 (
            .O(N__24732),
            .I(N__24705));
    Span12Mux_h I__5376 (
            .O(N__24729),
            .I(N__24702));
    LocalMux I__5375 (
            .O(N__24726),
            .I(N__24699));
    Span4Mux_v I__5374 (
            .O(N__24721),
            .I(N__24694));
    Span4Mux_v I__5373 (
            .O(N__24714),
            .I(N__24694));
    InMux I__5372 (
            .O(N__24711),
            .I(N__24691));
    Span12Mux_v I__5371 (
            .O(N__24708),
            .I(N__24683));
    Sp12to4 I__5370 (
            .O(N__24705),
            .I(N__24683));
    Span12Mux_v I__5369 (
            .O(N__24702),
            .I(N__24674));
    Span12Mux_h I__5368 (
            .O(N__24699),
            .I(N__24674));
    Sp12to4 I__5367 (
            .O(N__24694),
            .I(N__24674));
    LocalMux I__5366 (
            .O(N__24691),
            .I(N__24674));
    InMux I__5365 (
            .O(N__24690),
            .I(N__24671));
    InMux I__5364 (
            .O(N__24689),
            .I(N__24668));
    InMux I__5363 (
            .O(N__24688),
            .I(N__24665));
    Odrv12 I__5362 (
            .O(N__24683),
            .I(M_this_sprites_address_qZ0Z_10));
    Odrv12 I__5361 (
            .O(N__24674),
            .I(M_this_sprites_address_qZ0Z_10));
    LocalMux I__5360 (
            .O(N__24671),
            .I(M_this_sprites_address_qZ0Z_10));
    LocalMux I__5359 (
            .O(N__24668),
            .I(M_this_sprites_address_qZ0Z_10));
    LocalMux I__5358 (
            .O(N__24665),
            .I(M_this_sprites_address_qZ0Z_10));
    InMux I__5357 (
            .O(N__24654),
            .I(N__24651));
    LocalMux I__5356 (
            .O(N__24651),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10 ));
    CascadeMux I__5355 (
            .O(N__24648),
            .I(N__24645));
    InMux I__5354 (
            .O(N__24645),
            .I(N__24642));
    LocalMux I__5353 (
            .O(N__24642),
            .I(N__24639));
    Odrv4 I__5352 (
            .O(N__24639),
            .I(M_this_substate_q_RNOZ0Z_3));
    InMux I__5351 (
            .O(N__24636),
            .I(N__24633));
    LocalMux I__5350 (
            .O(N__24633),
            .I(N__24630));
    Span12Mux_h I__5349 (
            .O(N__24630),
            .I(N__24627));
    Span12Mux_v I__5348 (
            .O(N__24627),
            .I(N__24624));
    Odrv12 I__5347 (
            .O(N__24624),
            .I(\this_sprites_ram.mem_out_bus0_1 ));
    InMux I__5346 (
            .O(N__24621),
            .I(N__24618));
    LocalMux I__5345 (
            .O(N__24618),
            .I(N__24615));
    Span4Mux_h I__5344 (
            .O(N__24615),
            .I(N__24612));
    Span4Mux_h I__5343 (
            .O(N__24612),
            .I(N__24609));
    Span4Mux_h I__5342 (
            .O(N__24609),
            .I(N__24606));
    Span4Mux_h I__5341 (
            .O(N__24606),
            .I(N__24603));
    Odrv4 I__5340 (
            .O(N__24603),
            .I(\this_sprites_ram.mem_out_bus4_1 ));
    CascadeMux I__5339 (
            .O(N__24600),
            .I(N__24596));
    CascadeMux I__5338 (
            .O(N__24599),
            .I(N__24590));
    InMux I__5337 (
            .O(N__24596),
            .I(N__24582));
    InMux I__5336 (
            .O(N__24595),
            .I(N__24582));
    InMux I__5335 (
            .O(N__24594),
            .I(N__24577));
    InMux I__5334 (
            .O(N__24593),
            .I(N__24577));
    InMux I__5333 (
            .O(N__24590),
            .I(N__24574));
    InMux I__5332 (
            .O(N__24589),
            .I(N__24569));
    InMux I__5331 (
            .O(N__24588),
            .I(N__24569));
    InMux I__5330 (
            .O(N__24587),
            .I(N__24566));
    LocalMux I__5329 (
            .O(N__24582),
            .I(N__24561));
    LocalMux I__5328 (
            .O(N__24577),
            .I(N__24561));
    LocalMux I__5327 (
            .O(N__24574),
            .I(N__24554));
    LocalMux I__5326 (
            .O(N__24569),
            .I(N__24554));
    LocalMux I__5325 (
            .O(N__24566),
            .I(N__24554));
    Odrv4 I__5324 (
            .O(N__24561),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    Odrv4 I__5323 (
            .O(N__24554),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    CascadeMux I__5322 (
            .O(N__24549),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_ ));
    InMux I__5321 (
            .O(N__24546),
            .I(N__24543));
    LocalMux I__5320 (
            .O(N__24543),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1 ));
    InMux I__5319 (
            .O(N__24540),
            .I(N__24537));
    LocalMux I__5318 (
            .O(N__24537),
            .I(N__24534));
    Span4Mux_h I__5317 (
            .O(N__24534),
            .I(N__24531));
    Span4Mux_v I__5316 (
            .O(N__24531),
            .I(N__24528));
    Odrv4 I__5315 (
            .O(N__24528),
            .I(\this_sprites_ram.mem_out_bus6_1 ));
    InMux I__5314 (
            .O(N__24525),
            .I(N__24522));
    LocalMux I__5313 (
            .O(N__24522),
            .I(N__24519));
    Span4Mux_v I__5312 (
            .O(N__24519),
            .I(N__24516));
    Odrv4 I__5311 (
            .O(N__24516),
            .I(\this_sprites_ram.mem_out_bus2_1 ));
    InMux I__5310 (
            .O(N__24513),
            .I(N__24510));
    LocalMux I__5309 (
            .O(N__24510),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ));
    InMux I__5308 (
            .O(N__24507),
            .I(N__24504));
    LocalMux I__5307 (
            .O(N__24504),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12 ));
    InMux I__5306 (
            .O(N__24501),
            .I(N__24498));
    LocalMux I__5305 (
            .O(N__24498),
            .I(un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0));
    InMux I__5304 (
            .O(N__24495),
            .I(N__24492));
    LocalMux I__5303 (
            .O(N__24492),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0 ));
    InMux I__5302 (
            .O(N__24489),
            .I(N__24486));
    LocalMux I__5301 (
            .O(N__24486),
            .I(M_this_sprites_address_q_RNIQ61C7Z0Z_0));
    CascadeMux I__5300 (
            .O(N__24483),
            .I(N__24480));
    InMux I__5299 (
            .O(N__24480),
            .I(N__24477));
    LocalMux I__5298 (
            .O(N__24477),
            .I(N__24474));
    Span4Mux_h I__5297 (
            .O(N__24474),
            .I(N__24471));
    Odrv4 I__5296 (
            .O(N__24471),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_0 ));
    CascadeMux I__5295 (
            .O(N__24468),
            .I(N__24464));
    CascadeMux I__5294 (
            .O(N__24467),
            .I(N__24461));
    InMux I__5293 (
            .O(N__24464),
            .I(N__24457));
    InMux I__5292 (
            .O(N__24461),
            .I(N__24454));
    CascadeMux I__5291 (
            .O(N__24460),
            .I(N__24451));
    LocalMux I__5290 (
            .O(N__24457),
            .I(N__24446));
    LocalMux I__5289 (
            .O(N__24454),
            .I(N__24443));
    InMux I__5288 (
            .O(N__24451),
            .I(N__24440));
    CascadeMux I__5287 (
            .O(N__24450),
            .I(N__24437));
    CascadeMux I__5286 (
            .O(N__24449),
            .I(N__24434));
    Span4Mux_v I__5285 (
            .O(N__24446),
            .I(N__24420));
    Span4Mux_h I__5284 (
            .O(N__24443),
            .I(N__24420));
    LocalMux I__5283 (
            .O(N__24440),
            .I(N__24420));
    InMux I__5282 (
            .O(N__24437),
            .I(N__24417));
    InMux I__5281 (
            .O(N__24434),
            .I(N__24414));
    CascadeMux I__5280 (
            .O(N__24433),
            .I(N__24411));
    CascadeMux I__5279 (
            .O(N__24432),
            .I(N__24408));
    CascadeMux I__5278 (
            .O(N__24431),
            .I(N__24405));
    CascadeMux I__5277 (
            .O(N__24430),
            .I(N__24400));
    CascadeMux I__5276 (
            .O(N__24429),
            .I(N__24397));
    CascadeMux I__5275 (
            .O(N__24428),
            .I(N__24394));
    CascadeMux I__5274 (
            .O(N__24427),
            .I(N__24391));
    Span4Mux_v I__5273 (
            .O(N__24420),
            .I(N__24385));
    LocalMux I__5272 (
            .O(N__24417),
            .I(N__24385));
    LocalMux I__5271 (
            .O(N__24414),
            .I(N__24382));
    InMux I__5270 (
            .O(N__24411),
            .I(N__24379));
    InMux I__5269 (
            .O(N__24408),
            .I(N__24376));
    InMux I__5268 (
            .O(N__24405),
            .I(N__24373));
    CascadeMux I__5267 (
            .O(N__24404),
            .I(N__24370));
    CascadeMux I__5266 (
            .O(N__24403),
            .I(N__24367));
    InMux I__5265 (
            .O(N__24400),
            .I(N__24364));
    InMux I__5264 (
            .O(N__24397),
            .I(N__24361));
    InMux I__5263 (
            .O(N__24394),
            .I(N__24358));
    InMux I__5262 (
            .O(N__24391),
            .I(N__24355));
    CascadeMux I__5261 (
            .O(N__24390),
            .I(N__24352));
    Span4Mux_v I__5260 (
            .O(N__24385),
            .I(N__24345));
    Span4Mux_h I__5259 (
            .O(N__24382),
            .I(N__24345));
    LocalMux I__5258 (
            .O(N__24379),
            .I(N__24345));
    LocalMux I__5257 (
            .O(N__24376),
            .I(N__24340));
    LocalMux I__5256 (
            .O(N__24373),
            .I(N__24340));
    InMux I__5255 (
            .O(N__24370),
            .I(N__24337));
    InMux I__5254 (
            .O(N__24367),
            .I(N__24334));
    LocalMux I__5253 (
            .O(N__24364),
            .I(N__24325));
    LocalMux I__5252 (
            .O(N__24361),
            .I(N__24325));
    LocalMux I__5251 (
            .O(N__24358),
            .I(N__24325));
    LocalMux I__5250 (
            .O(N__24355),
            .I(N__24322));
    InMux I__5249 (
            .O(N__24352),
            .I(N__24319));
    Span4Mux_v I__5248 (
            .O(N__24345),
            .I(N__24316));
    Span4Mux_v I__5247 (
            .O(N__24340),
            .I(N__24309));
    LocalMux I__5246 (
            .O(N__24337),
            .I(N__24309));
    LocalMux I__5245 (
            .O(N__24334),
            .I(N__24309));
    CascadeMux I__5244 (
            .O(N__24333),
            .I(N__24306));
    InMux I__5243 (
            .O(N__24332),
            .I(N__24303));
    Span12Mux_v I__5242 (
            .O(N__24325),
            .I(N__24300));
    Span12Mux_h I__5241 (
            .O(N__24322),
            .I(N__24297));
    LocalMux I__5240 (
            .O(N__24319),
            .I(N__24294));
    Span4Mux_v I__5239 (
            .O(N__24316),
            .I(N__24289));
    Span4Mux_v I__5238 (
            .O(N__24309),
            .I(N__24289));
    InMux I__5237 (
            .O(N__24306),
            .I(N__24286));
    LocalMux I__5236 (
            .O(N__24303),
            .I(N__24283));
    Span12Mux_h I__5235 (
            .O(N__24300),
            .I(N__24278));
    Span12Mux_v I__5234 (
            .O(N__24297),
            .I(N__24269));
    Span12Mux_h I__5233 (
            .O(N__24294),
            .I(N__24269));
    Sp12to4 I__5232 (
            .O(N__24289),
            .I(N__24269));
    LocalMux I__5231 (
            .O(N__24286),
            .I(N__24269));
    Span4Mux_h I__5230 (
            .O(N__24283),
            .I(N__24266));
    InMux I__5229 (
            .O(N__24282),
            .I(N__24263));
    InMux I__5228 (
            .O(N__24281),
            .I(N__24260));
    Odrv12 I__5227 (
            .O(N__24278),
            .I(M_this_sprites_address_qZ0Z_0));
    Odrv12 I__5226 (
            .O(N__24269),
            .I(M_this_sprites_address_qZ0Z_0));
    Odrv4 I__5225 (
            .O(N__24266),
            .I(M_this_sprites_address_qZ0Z_0));
    LocalMux I__5224 (
            .O(N__24263),
            .I(M_this_sprites_address_qZ0Z_0));
    LocalMux I__5223 (
            .O(N__24260),
            .I(M_this_sprites_address_qZ0Z_0));
    CascadeMux I__5222 (
            .O(N__24249),
            .I(N__24246));
    InMux I__5221 (
            .O(N__24246),
            .I(N__24243));
    LocalMux I__5220 (
            .O(N__24243),
            .I(N__24240));
    Odrv4 I__5219 (
            .O(N__24240),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_11 ));
    InMux I__5218 (
            .O(N__24237),
            .I(N__24234));
    LocalMux I__5217 (
            .O(N__24234),
            .I(N__24231));
    Odrv4 I__5216 (
            .O(N__24231),
            .I(M_this_substate_q_RNOZ0Z_1));
    InMux I__5215 (
            .O(N__24228),
            .I(N__24225));
    LocalMux I__5214 (
            .O(N__24225),
            .I(N__24222));
    Odrv12 I__5213 (
            .O(N__24222),
            .I(M_this_substate_q_s_1));
    InMux I__5212 (
            .O(N__24219),
            .I(N__24215));
    InMux I__5211 (
            .O(N__24218),
            .I(N__24212));
    LocalMux I__5210 (
            .O(N__24215),
            .I(N__24209));
    LocalMux I__5209 (
            .O(N__24212),
            .I(this_vga_signals_M_this_state_d_2_sqmuxa_0));
    Odrv4 I__5208 (
            .O(N__24209),
            .I(this_vga_signals_M_this_state_d_2_sqmuxa_0));
    InMux I__5207 (
            .O(N__24204),
            .I(N__24201));
    LocalMux I__5206 (
            .O(N__24201),
            .I(N__24196));
    InMux I__5205 (
            .O(N__24200),
            .I(N__24193));
    InMux I__5204 (
            .O(N__24199),
            .I(N__24190));
    Odrv4 I__5203 (
            .O(N__24196),
            .I(N_17_0));
    LocalMux I__5202 (
            .O(N__24193),
            .I(N_17_0));
    LocalMux I__5201 (
            .O(N__24190),
            .I(N_17_0));
    CascadeMux I__5200 (
            .O(N__24183),
            .I(N__24179));
    CascadeMux I__5199 (
            .O(N__24182),
            .I(N__24173));
    InMux I__5198 (
            .O(N__24179),
            .I(N__24170));
    CascadeMux I__5197 (
            .O(N__24178),
            .I(N__24167));
    CascadeMux I__5196 (
            .O(N__24177),
            .I(N__24160));
    CascadeMux I__5195 (
            .O(N__24176),
            .I(N__24156));
    InMux I__5194 (
            .O(N__24173),
            .I(N__24152));
    LocalMux I__5193 (
            .O(N__24170),
            .I(N__24149));
    InMux I__5192 (
            .O(N__24167),
            .I(N__24146));
    CascadeMux I__5191 (
            .O(N__24166),
            .I(N__24143));
    CascadeMux I__5190 (
            .O(N__24165),
            .I(N__24140));
    CascadeMux I__5189 (
            .O(N__24164),
            .I(N__24137));
    CascadeMux I__5188 (
            .O(N__24163),
            .I(N__24134));
    InMux I__5187 (
            .O(N__24160),
            .I(N__24127));
    CascadeMux I__5186 (
            .O(N__24159),
            .I(N__24124));
    InMux I__5185 (
            .O(N__24156),
            .I(N__24121));
    CascadeMux I__5184 (
            .O(N__24155),
            .I(N__24118));
    LocalMux I__5183 (
            .O(N__24152),
            .I(N__24111));
    Span4Mux_v I__5182 (
            .O(N__24149),
            .I(N__24111));
    LocalMux I__5181 (
            .O(N__24146),
            .I(N__24111));
    InMux I__5180 (
            .O(N__24143),
            .I(N__24108));
    InMux I__5179 (
            .O(N__24140),
            .I(N__24105));
    InMux I__5178 (
            .O(N__24137),
            .I(N__24102));
    InMux I__5177 (
            .O(N__24134),
            .I(N__24099));
    CascadeMux I__5176 (
            .O(N__24133),
            .I(N__24095));
    CascadeMux I__5175 (
            .O(N__24132),
            .I(N__24092));
    CascadeMux I__5174 (
            .O(N__24131),
            .I(N__24089));
    CascadeMux I__5173 (
            .O(N__24130),
            .I(N__24086));
    LocalMux I__5172 (
            .O(N__24127),
            .I(N__24083));
    InMux I__5171 (
            .O(N__24124),
            .I(N__24080));
    LocalMux I__5170 (
            .O(N__24121),
            .I(N__24077));
    InMux I__5169 (
            .O(N__24118),
            .I(N__24074));
    Span4Mux_v I__5168 (
            .O(N__24111),
            .I(N__24067));
    LocalMux I__5167 (
            .O(N__24108),
            .I(N__24067));
    LocalMux I__5166 (
            .O(N__24105),
            .I(N__24067));
    LocalMux I__5165 (
            .O(N__24102),
            .I(N__24062));
    LocalMux I__5164 (
            .O(N__24099),
            .I(N__24062));
    CascadeMux I__5163 (
            .O(N__24098),
            .I(N__24059));
    InMux I__5162 (
            .O(N__24095),
            .I(N__24056));
    InMux I__5161 (
            .O(N__24092),
            .I(N__24053));
    InMux I__5160 (
            .O(N__24089),
            .I(N__24050));
    InMux I__5159 (
            .O(N__24086),
            .I(N__24047));
    Span4Mux_v I__5158 (
            .O(N__24083),
            .I(N__24042));
    LocalMux I__5157 (
            .O(N__24080),
            .I(N__24042));
    Span4Mux_h I__5156 (
            .O(N__24077),
            .I(N__24039));
    LocalMux I__5155 (
            .O(N__24074),
            .I(N__24035));
    Span4Mux_v I__5154 (
            .O(N__24067),
            .I(N__24030));
    Span4Mux_v I__5153 (
            .O(N__24062),
            .I(N__24030));
    InMux I__5152 (
            .O(N__24059),
            .I(N__24026));
    LocalMux I__5151 (
            .O(N__24056),
            .I(N__24023));
    LocalMux I__5150 (
            .O(N__24053),
            .I(N__24020));
    LocalMux I__5149 (
            .O(N__24050),
            .I(N__24017));
    LocalMux I__5148 (
            .O(N__24047),
            .I(N__24014));
    Span4Mux_h I__5147 (
            .O(N__24042),
            .I(N__24009));
    Span4Mux_v I__5146 (
            .O(N__24039),
            .I(N__24009));
    CascadeMux I__5145 (
            .O(N__24038),
            .I(N__24006));
    Span4Mux_h I__5144 (
            .O(N__24035),
            .I(N__24003));
    Sp12to4 I__5143 (
            .O(N__24030),
            .I(N__24000));
    InMux I__5142 (
            .O(N__24029),
            .I(N__23996));
    LocalMux I__5141 (
            .O(N__24026),
            .I(N__23989));
    Span4Mux_v I__5140 (
            .O(N__24023),
            .I(N__23989));
    Span4Mux_v I__5139 (
            .O(N__24020),
            .I(N__23989));
    Span4Mux_h I__5138 (
            .O(N__24017),
            .I(N__23986));
    Span4Mux_h I__5137 (
            .O(N__24014),
            .I(N__23981));
    Span4Mux_v I__5136 (
            .O(N__24009),
            .I(N__23981));
    InMux I__5135 (
            .O(N__24006),
            .I(N__23978));
    Span4Mux_h I__5134 (
            .O(N__24003),
            .I(N__23975));
    Span12Mux_h I__5133 (
            .O(N__24000),
            .I(N__23972));
    InMux I__5132 (
            .O(N__23999),
            .I(N__23969));
    LocalMux I__5131 (
            .O(N__23996),
            .I(N__23962));
    Span4Mux_h I__5130 (
            .O(N__23989),
            .I(N__23962));
    Span4Mux_v I__5129 (
            .O(N__23986),
            .I(N__23962));
    Span4Mux_h I__5128 (
            .O(N__23981),
            .I(N__23959));
    LocalMux I__5127 (
            .O(N__23978),
            .I(N__23956));
    Sp12to4 I__5126 (
            .O(N__23975),
            .I(N__23951));
    Span12Mux_v I__5125 (
            .O(N__23972),
            .I(N__23951));
    LocalMux I__5124 (
            .O(N__23969),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv4 I__5123 (
            .O(N__23962),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv4 I__5122 (
            .O(N__23959),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv4 I__5121 (
            .O(N__23956),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv12 I__5120 (
            .O(N__23951),
            .I(M_this_sprites_address_qZ0Z_3));
    InMux I__5119 (
            .O(N__23940),
            .I(N__23937));
    LocalMux I__5118 (
            .O(N__23937),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_3 ));
    CascadeMux I__5117 (
            .O(N__23934),
            .I(N__23931));
    InMux I__5116 (
            .O(N__23931),
            .I(N__23928));
    LocalMux I__5115 (
            .O(N__23928),
            .I(N__23925));
    Odrv12 I__5114 (
            .O(N__23925),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_12 ));
    CascadeMux I__5113 (
            .O(N__23922),
            .I(N__23919));
    InMux I__5112 (
            .O(N__23919),
            .I(N__23916));
    LocalMux I__5111 (
            .O(N__23916),
            .I(N__23913));
    Odrv12 I__5110 (
            .O(N__23913),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_13 ));
    CascadeMux I__5109 (
            .O(N__23910),
            .I(N__23907));
    InMux I__5108 (
            .O(N__23907),
            .I(N__23901));
    InMux I__5107 (
            .O(N__23906),
            .I(N__23898));
    InMux I__5106 (
            .O(N__23905),
            .I(N__23893));
    InMux I__5105 (
            .O(N__23904),
            .I(N__23893));
    LocalMux I__5104 (
            .O(N__23901),
            .I(\this_ppu.N_1046_0 ));
    LocalMux I__5103 (
            .O(N__23898),
            .I(\this_ppu.N_1046_0 ));
    LocalMux I__5102 (
            .O(N__23893),
            .I(\this_ppu.N_1046_0 ));
    InMux I__5101 (
            .O(N__23886),
            .I(N__23882));
    InMux I__5100 (
            .O(N__23885),
            .I(N__23879));
    LocalMux I__5099 (
            .O(N__23882),
            .I(\this_ppu.un1_M_oam_idx_q_1_c1 ));
    LocalMux I__5098 (
            .O(N__23879),
            .I(\this_ppu.un1_M_oam_idx_q_1_c1 ));
    CascadeMux I__5097 (
            .O(N__23874),
            .I(N__23871));
    CascadeBuf I__5096 (
            .O(N__23871),
            .I(N__23868));
    CascadeMux I__5095 (
            .O(N__23868),
            .I(N__23865));
    InMux I__5094 (
            .O(N__23865),
            .I(N__23858));
    InMux I__5093 (
            .O(N__23864),
            .I(N__23855));
    InMux I__5092 (
            .O(N__23863),
            .I(N__23848));
    InMux I__5091 (
            .O(N__23862),
            .I(N__23848));
    InMux I__5090 (
            .O(N__23861),
            .I(N__23848));
    LocalMux I__5089 (
            .O(N__23858),
            .I(N__23845));
    LocalMux I__5088 (
            .O(N__23855),
            .I(M_this_ppu_oam_addr_1));
    LocalMux I__5087 (
            .O(N__23848),
            .I(M_this_ppu_oam_addr_1));
    Odrv12 I__5086 (
            .O(N__23845),
            .I(M_this_ppu_oam_addr_1));
    CascadeMux I__5085 (
            .O(N__23838),
            .I(N__23835));
    CascadeBuf I__5084 (
            .O(N__23835),
            .I(N__23832));
    CascadeMux I__5083 (
            .O(N__23832),
            .I(N__23829));
    InMux I__5082 (
            .O(N__23829),
            .I(N__23826));
    LocalMux I__5081 (
            .O(N__23826),
            .I(N__23822));
    InMux I__5080 (
            .O(N__23825),
            .I(N__23816));
    Span4Mux_h I__5079 (
            .O(N__23822),
            .I(N__23813));
    InMux I__5078 (
            .O(N__23821),
            .I(N__23810));
    InMux I__5077 (
            .O(N__23820),
            .I(N__23805));
    InMux I__5076 (
            .O(N__23819),
            .I(N__23805));
    LocalMux I__5075 (
            .O(N__23816),
            .I(N__23802));
    Span4Mux_h I__5074 (
            .O(N__23813),
            .I(N__23799));
    LocalMux I__5073 (
            .O(N__23810),
            .I(M_this_ppu_oam_addr_3));
    LocalMux I__5072 (
            .O(N__23805),
            .I(M_this_ppu_oam_addr_3));
    Odrv4 I__5071 (
            .O(N__23802),
            .I(M_this_ppu_oam_addr_3));
    Odrv4 I__5070 (
            .O(N__23799),
            .I(M_this_ppu_oam_addr_3));
    InMux I__5069 (
            .O(N__23790),
            .I(N__23787));
    LocalMux I__5068 (
            .O(N__23787),
            .I(\this_ppu.N_144_4 ));
    CascadeMux I__5067 (
            .O(N__23784),
            .I(N__23781));
    InMux I__5066 (
            .O(N__23781),
            .I(N__23778));
    LocalMux I__5065 (
            .O(N__23778),
            .I(N__23775));
    Span4Mux_h I__5064 (
            .O(N__23775),
            .I(N__23772));
    Odrv4 I__5063 (
            .O(N__23772),
            .I(\this_ppu.N_144 ));
    CascadeMux I__5062 (
            .O(N__23769),
            .I(N__23764));
    InMux I__5061 (
            .O(N__23768),
            .I(N__23760));
    CascadeMux I__5060 (
            .O(N__23767),
            .I(N__23757));
    InMux I__5059 (
            .O(N__23764),
            .I(N__23754));
    InMux I__5058 (
            .O(N__23763),
            .I(N__23751));
    LocalMux I__5057 (
            .O(N__23760),
            .I(N__23747));
    InMux I__5056 (
            .O(N__23757),
            .I(N__23744));
    LocalMux I__5055 (
            .O(N__23754),
            .I(N__23741));
    LocalMux I__5054 (
            .O(N__23751),
            .I(N__23738));
    CascadeMux I__5053 (
            .O(N__23750),
            .I(N__23735));
    Span4Mux_v I__5052 (
            .O(N__23747),
            .I(N__23730));
    LocalMux I__5051 (
            .O(N__23744),
            .I(N__23730));
    Span4Mux_v I__5050 (
            .O(N__23741),
            .I(N__23723));
    Span4Mux_v I__5049 (
            .O(N__23738),
            .I(N__23723));
    InMux I__5048 (
            .O(N__23735),
            .I(N__23720));
    Span4Mux_h I__5047 (
            .O(N__23730),
            .I(N__23717));
    InMux I__5046 (
            .O(N__23729),
            .I(N__23712));
    InMux I__5045 (
            .O(N__23728),
            .I(N__23712));
    Odrv4 I__5044 (
            .O(N__23723),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__5043 (
            .O(N__23720),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__5042 (
            .O(N__23717),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__5041 (
            .O(N__23712),
            .I(M_this_state_qZ0Z_8));
    InMux I__5040 (
            .O(N__23703),
            .I(N__23698));
    InMux I__5039 (
            .O(N__23702),
            .I(N__23694));
    InMux I__5038 (
            .O(N__23701),
            .I(N__23691));
    LocalMux I__5037 (
            .O(N__23698),
            .I(N__23687));
    InMux I__5036 (
            .O(N__23697),
            .I(N__23684));
    LocalMux I__5035 (
            .O(N__23694),
            .I(N__23681));
    LocalMux I__5034 (
            .O(N__23691),
            .I(N__23678));
    InMux I__5033 (
            .O(N__23690),
            .I(N__23674));
    Span4Mux_v I__5032 (
            .O(N__23687),
            .I(N__23670));
    LocalMux I__5031 (
            .O(N__23684),
            .I(N__23663));
    Span4Mux_v I__5030 (
            .O(N__23681),
            .I(N__23663));
    Span4Mux_v I__5029 (
            .O(N__23678),
            .I(N__23663));
    InMux I__5028 (
            .O(N__23677),
            .I(N__23660));
    LocalMux I__5027 (
            .O(N__23674),
            .I(N__23657));
    InMux I__5026 (
            .O(N__23673),
            .I(N__23654));
    Odrv4 I__5025 (
            .O(N__23670),
            .I(M_this_state_qZ0Z_7));
    Odrv4 I__5024 (
            .O(N__23663),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__5023 (
            .O(N__23660),
            .I(M_this_state_qZ0Z_7));
    Odrv4 I__5022 (
            .O(N__23657),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__5021 (
            .O(N__23654),
            .I(M_this_state_qZ0Z_7));
    InMux I__5020 (
            .O(N__23643),
            .I(N__23638));
    InMux I__5019 (
            .O(N__23642),
            .I(N__23633));
    InMux I__5018 (
            .O(N__23641),
            .I(N__23630));
    LocalMux I__5017 (
            .O(N__23638),
            .I(N__23626));
    InMux I__5016 (
            .O(N__23637),
            .I(N__23623));
    InMux I__5015 (
            .O(N__23636),
            .I(N__23620));
    LocalMux I__5014 (
            .O(N__23633),
            .I(N__23615));
    LocalMux I__5013 (
            .O(N__23630),
            .I(N__23612));
    InMux I__5012 (
            .O(N__23629),
            .I(N__23609));
    Span12Mux_s8_v I__5011 (
            .O(N__23626),
            .I(N__23602));
    LocalMux I__5010 (
            .O(N__23623),
            .I(N__23602));
    LocalMux I__5009 (
            .O(N__23620),
            .I(N__23602));
    InMux I__5008 (
            .O(N__23619),
            .I(N__23599));
    InMux I__5007 (
            .O(N__23618),
            .I(N__23596));
    Span12Mux_v I__5006 (
            .O(N__23615),
            .I(N__23591));
    Span12Mux_v I__5005 (
            .O(N__23612),
            .I(N__23591));
    LocalMux I__5004 (
            .O(N__23609),
            .I(N__23582));
    Span12Mux_v I__5003 (
            .O(N__23602),
            .I(N__23582));
    LocalMux I__5002 (
            .O(N__23599),
            .I(N__23582));
    LocalMux I__5001 (
            .O(N__23596),
            .I(N__23582));
    Span12Mux_h I__5000 (
            .O(N__23591),
            .I(N__23579));
    Span12Mux_s11_v I__4999 (
            .O(N__23582),
            .I(N__23576));
    Odrv12 I__4998 (
            .O(N__23579),
            .I(M_this_sprites_ram_write_data_2));
    Odrv12 I__4997 (
            .O(N__23576),
            .I(M_this_sprites_ram_write_data_2));
    CEMux I__4996 (
            .O(N__23571),
            .I(N__23567));
    CEMux I__4995 (
            .O(N__23570),
            .I(N__23564));
    LocalMux I__4994 (
            .O(N__23567),
            .I(N__23561));
    LocalMux I__4993 (
            .O(N__23564),
            .I(N__23558));
    Span4Mux_h I__4992 (
            .O(N__23561),
            .I(N__23555));
    Span4Mux_h I__4991 (
            .O(N__23558),
            .I(N__23552));
    Span4Mux_h I__4990 (
            .O(N__23555),
            .I(N__23549));
    Span4Mux_h I__4989 (
            .O(N__23552),
            .I(N__23546));
    Span4Mux_h I__4988 (
            .O(N__23549),
            .I(N__23543));
    Span4Mux_h I__4987 (
            .O(N__23546),
            .I(N__23540));
    Odrv4 I__4986 (
            .O(N__23543),
            .I(\this_sprites_ram.mem_WE_6 ));
    Odrv4 I__4985 (
            .O(N__23540),
            .I(\this_sprites_ram.mem_WE_6 ));
    InMux I__4984 (
            .O(N__23535),
            .I(N__23532));
    LocalMux I__4983 (
            .O(N__23532),
            .I(un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0));
    InMux I__4982 (
            .O(N__23529),
            .I(N__23526));
    LocalMux I__4981 (
            .O(N__23526),
            .I(N__23523));
    Span4Mux_v I__4980 (
            .O(N__23523),
            .I(N__23520));
    Odrv4 I__4979 (
            .O(N__23520),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13 ));
    InMux I__4978 (
            .O(N__23517),
            .I(N__23514));
    LocalMux I__4977 (
            .O(N__23514),
            .I(un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0));
    CascadeMux I__4976 (
            .O(N__23511),
            .I(\this_ppu.N_1046_0_cascade_ ));
    InMux I__4975 (
            .O(N__23508),
            .I(N__23501));
    InMux I__4974 (
            .O(N__23507),
            .I(N__23496));
    InMux I__4973 (
            .O(N__23506),
            .I(N__23496));
    InMux I__4972 (
            .O(N__23505),
            .I(N__23491));
    InMux I__4971 (
            .O(N__23504),
            .I(N__23491));
    LocalMux I__4970 (
            .O(N__23501),
            .I(N__23484));
    LocalMux I__4969 (
            .O(N__23496),
            .I(N__23484));
    LocalMux I__4968 (
            .O(N__23491),
            .I(N__23484));
    Odrv4 I__4967 (
            .O(N__23484),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    CascadeMux I__4966 (
            .O(N__23481),
            .I(\this_ppu.un1_M_oam_idx_q_1_c1_cascade_ ));
    InMux I__4965 (
            .O(N__23478),
            .I(N__23472));
    InMux I__4964 (
            .O(N__23477),
            .I(N__23472));
    LocalMux I__4963 (
            .O(N__23472),
            .I(\this_ppu.un1_M_oam_idx_q_1_c3 ));
    CascadeMux I__4962 (
            .O(N__23469),
            .I(N__23466));
    CascadeBuf I__4961 (
            .O(N__23466),
            .I(N__23463));
    CascadeMux I__4960 (
            .O(N__23463),
            .I(N__23460));
    InMux I__4959 (
            .O(N__23460),
            .I(N__23457));
    LocalMux I__4958 (
            .O(N__23457),
            .I(N__23453));
    CascadeMux I__4957 (
            .O(N__23456),
            .I(N__23450));
    Span4Mux_h I__4956 (
            .O(N__23453),
            .I(N__23445));
    InMux I__4955 (
            .O(N__23450),
            .I(N__23442));
    InMux I__4954 (
            .O(N__23449),
            .I(N__23437));
    InMux I__4953 (
            .O(N__23448),
            .I(N__23437));
    Span4Mux_h I__4952 (
            .O(N__23445),
            .I(N__23434));
    LocalMux I__4951 (
            .O(N__23442),
            .I(M_this_ppu_oam_addr_2));
    LocalMux I__4950 (
            .O(N__23437),
            .I(M_this_ppu_oam_addr_2));
    Odrv4 I__4949 (
            .O(N__23434),
            .I(M_this_ppu_oam_addr_2));
    CascadeMux I__4948 (
            .O(N__23427),
            .I(N__23424));
    CascadeBuf I__4947 (
            .O(N__23424),
            .I(N__23421));
    CascadeMux I__4946 (
            .O(N__23421),
            .I(N__23417));
    CascadeMux I__4945 (
            .O(N__23420),
            .I(N__23414));
    InMux I__4944 (
            .O(N__23417),
            .I(N__23409));
    InMux I__4943 (
            .O(N__23414),
            .I(N__23402));
    InMux I__4942 (
            .O(N__23413),
            .I(N__23402));
    InMux I__4941 (
            .O(N__23412),
            .I(N__23402));
    LocalMux I__4940 (
            .O(N__23409),
            .I(N__23399));
    LocalMux I__4939 (
            .O(N__23402),
            .I(M_this_ppu_oam_addr_0));
    Odrv12 I__4938 (
            .O(N__23399),
            .I(M_this_ppu_oam_addr_0));
    CascadeMux I__4937 (
            .O(N__23394),
            .I(N__23390));
    InMux I__4936 (
            .O(N__23393),
            .I(N__23387));
    InMux I__4935 (
            .O(N__23390),
            .I(N__23384));
    LocalMux I__4934 (
            .O(N__23387),
            .I(\this_ppu.M_oam_idx_qZ0Z_4 ));
    LocalMux I__4933 (
            .O(N__23384),
            .I(\this_ppu.M_oam_idx_qZ0Z_4 ));
    CascadeMux I__4932 (
            .O(N__23379),
            .I(\this_ppu.N_144_4_cascade_ ));
    InMux I__4931 (
            .O(N__23376),
            .I(N__23373));
    LocalMux I__4930 (
            .O(N__23373),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    InMux I__4929 (
            .O(N__23370),
            .I(N__23367));
    LocalMux I__4928 (
            .O(N__23367),
            .I(N__23362));
    InMux I__4927 (
            .O(N__23366),
            .I(N__23359));
    InMux I__4926 (
            .O(N__23365),
            .I(N__23356));
    Odrv4 I__4925 (
            .O(N__23362),
            .I(\this_ppu.N_156 ));
    LocalMux I__4924 (
            .O(N__23359),
            .I(\this_ppu.N_156 ));
    LocalMux I__4923 (
            .O(N__23356),
            .I(\this_ppu.N_156 ));
    CascadeMux I__4922 (
            .O(N__23349),
            .I(\this_ppu.un2_hscroll_axb_0_cascade_ ));
    CascadeMux I__4921 (
            .O(N__23346),
            .I(N__23340));
    CascadeMux I__4920 (
            .O(N__23345),
            .I(N__23335));
    CascadeMux I__4919 (
            .O(N__23344),
            .I(N__23329));
    CascadeMux I__4918 (
            .O(N__23343),
            .I(N__23326));
    InMux I__4917 (
            .O(N__23340),
            .I(N__23321));
    CascadeMux I__4916 (
            .O(N__23339),
            .I(N__23318));
    CascadeMux I__4915 (
            .O(N__23338),
            .I(N__23315));
    InMux I__4914 (
            .O(N__23335),
            .I(N__23310));
    CascadeMux I__4913 (
            .O(N__23334),
            .I(N__23307));
    CascadeMux I__4912 (
            .O(N__23333),
            .I(N__23304));
    CascadeMux I__4911 (
            .O(N__23332),
            .I(N__23301));
    InMux I__4910 (
            .O(N__23329),
            .I(N__23298));
    InMux I__4909 (
            .O(N__23326),
            .I(N__23295));
    CascadeMux I__4908 (
            .O(N__23325),
            .I(N__23292));
    CascadeMux I__4907 (
            .O(N__23324),
            .I(N__23289));
    LocalMux I__4906 (
            .O(N__23321),
            .I(N__23285));
    InMux I__4905 (
            .O(N__23318),
            .I(N__23282));
    InMux I__4904 (
            .O(N__23315),
            .I(N__23279));
    CascadeMux I__4903 (
            .O(N__23314),
            .I(N__23276));
    CascadeMux I__4902 (
            .O(N__23313),
            .I(N__23273));
    LocalMux I__4901 (
            .O(N__23310),
            .I(N__23268));
    InMux I__4900 (
            .O(N__23307),
            .I(N__23265));
    InMux I__4899 (
            .O(N__23304),
            .I(N__23262));
    InMux I__4898 (
            .O(N__23301),
            .I(N__23259));
    LocalMux I__4897 (
            .O(N__23298),
            .I(N__23254));
    LocalMux I__4896 (
            .O(N__23295),
            .I(N__23254));
    InMux I__4895 (
            .O(N__23292),
            .I(N__23251));
    InMux I__4894 (
            .O(N__23289),
            .I(N__23248));
    CascadeMux I__4893 (
            .O(N__23288),
            .I(N__23245));
    Span4Mux_s2_v I__4892 (
            .O(N__23285),
            .I(N__23240));
    LocalMux I__4891 (
            .O(N__23282),
            .I(N__23240));
    LocalMux I__4890 (
            .O(N__23279),
            .I(N__23237));
    InMux I__4889 (
            .O(N__23276),
            .I(N__23234));
    InMux I__4888 (
            .O(N__23273),
            .I(N__23231));
    CascadeMux I__4887 (
            .O(N__23272),
            .I(N__23228));
    CascadeMux I__4886 (
            .O(N__23271),
            .I(N__23225));
    Span4Mux_v I__4885 (
            .O(N__23268),
            .I(N__23220));
    LocalMux I__4884 (
            .O(N__23265),
            .I(N__23220));
    LocalMux I__4883 (
            .O(N__23262),
            .I(N__23217));
    LocalMux I__4882 (
            .O(N__23259),
            .I(N__23214));
    Span4Mux_v I__4881 (
            .O(N__23254),
            .I(N__23207));
    LocalMux I__4880 (
            .O(N__23251),
            .I(N__23207));
    LocalMux I__4879 (
            .O(N__23248),
            .I(N__23207));
    InMux I__4878 (
            .O(N__23245),
            .I(N__23204));
    Span4Mux_v I__4877 (
            .O(N__23240),
            .I(N__23197));
    Span4Mux_h I__4876 (
            .O(N__23237),
            .I(N__23197));
    LocalMux I__4875 (
            .O(N__23234),
            .I(N__23197));
    LocalMux I__4874 (
            .O(N__23231),
            .I(N__23194));
    InMux I__4873 (
            .O(N__23228),
            .I(N__23191));
    InMux I__4872 (
            .O(N__23225),
            .I(N__23188));
    Span4Mux_v I__4871 (
            .O(N__23220),
            .I(N__23181));
    Span4Mux_v I__4870 (
            .O(N__23217),
            .I(N__23181));
    Span4Mux_v I__4869 (
            .O(N__23214),
            .I(N__23181));
    Span4Mux_v I__4868 (
            .O(N__23207),
            .I(N__23176));
    LocalMux I__4867 (
            .O(N__23204),
            .I(N__23176));
    Span4Mux_v I__4866 (
            .O(N__23197),
            .I(N__23169));
    Span4Mux_h I__4865 (
            .O(N__23194),
            .I(N__23169));
    LocalMux I__4864 (
            .O(N__23191),
            .I(N__23169));
    LocalMux I__4863 (
            .O(N__23188),
            .I(N__23166));
    Span4Mux_h I__4862 (
            .O(N__23181),
            .I(N__23163));
    Span4Mux_h I__4861 (
            .O(N__23176),
            .I(N__23160));
    Span4Mux_v I__4860 (
            .O(N__23169),
            .I(N__23155));
    Span4Mux_h I__4859 (
            .O(N__23166),
            .I(N__23155));
    Span4Mux_h I__4858 (
            .O(N__23163),
            .I(N__23152));
    Span4Mux_v I__4857 (
            .O(N__23160),
            .I(N__23149));
    Span4Mux_h I__4856 (
            .O(N__23155),
            .I(N__23146));
    Odrv4 I__4855 (
            .O(N__23152),
            .I(M_this_ppu_sprites_addr_0));
    Odrv4 I__4854 (
            .O(N__23149),
            .I(M_this_ppu_sprites_addr_0));
    Odrv4 I__4853 (
            .O(N__23146),
            .I(M_this_ppu_sprites_addr_0));
    InMux I__4852 (
            .O(N__23139),
            .I(N__23133));
    InMux I__4851 (
            .O(N__23138),
            .I(N__23133));
    LocalMux I__4850 (
            .O(N__23133),
            .I(\this_ppu.un1_M_haddress_q_3_c2 ));
    SRMux I__4849 (
            .O(N__23130),
            .I(N__23126));
    SRMux I__4848 (
            .O(N__23129),
            .I(N__23123));
    LocalMux I__4847 (
            .O(N__23126),
            .I(\this_ppu.M_state_q_RNIGL6V4Z0Z_0 ));
    LocalMux I__4846 (
            .O(N__23123),
            .I(\this_ppu.M_state_q_RNIGL6V4Z0Z_0 ));
    CEMux I__4845 (
            .O(N__23118),
            .I(N__23115));
    LocalMux I__4844 (
            .O(N__23115),
            .I(N__23111));
    CEMux I__4843 (
            .O(N__23114),
            .I(N__23108));
    Span4Mux_h I__4842 (
            .O(N__23111),
            .I(N__23105));
    LocalMux I__4841 (
            .O(N__23108),
            .I(N__23102));
    Span4Mux_h I__4840 (
            .O(N__23105),
            .I(N__23099));
    Span4Mux_h I__4839 (
            .O(N__23102),
            .I(N__23096));
    Span4Mux_h I__4838 (
            .O(N__23099),
            .I(N__23093));
    Span4Mux_h I__4837 (
            .O(N__23096),
            .I(N__23090));
    Odrv4 I__4836 (
            .O(N__23093),
            .I(\this_sprites_ram.mem_WE_8 ));
    Odrv4 I__4835 (
            .O(N__23090),
            .I(\this_sprites_ram.mem_WE_8 ));
    CEMux I__4834 (
            .O(N__23085),
            .I(N__23081));
    CEMux I__4833 (
            .O(N__23084),
            .I(N__23078));
    LocalMux I__4832 (
            .O(N__23081),
            .I(N__23073));
    LocalMux I__4831 (
            .O(N__23078),
            .I(N__23073));
    Span4Mux_v I__4830 (
            .O(N__23073),
            .I(N__23070));
    Span4Mux_v I__4829 (
            .O(N__23070),
            .I(N__23067));
    Span4Mux_h I__4828 (
            .O(N__23067),
            .I(N__23064));
    Odrv4 I__4827 (
            .O(N__23064),
            .I(\this_sprites_ram.mem_WE_14 ));
    InMux I__4826 (
            .O(N__23061),
            .I(N__23058));
    LocalMux I__4825 (
            .O(N__23058),
            .I(N__23055));
    Span12Mux_h I__4824 (
            .O(N__23055),
            .I(N__23052));
    Span12Mux_v I__4823 (
            .O(N__23052),
            .I(N__23049));
    Odrv12 I__4822 (
            .O(N__23049),
            .I(\this_sprites_ram.mem_out_bus7_1 ));
    InMux I__4821 (
            .O(N__23046),
            .I(N__23043));
    LocalMux I__4820 (
            .O(N__23043),
            .I(N__23040));
    Span4Mux_h I__4819 (
            .O(N__23040),
            .I(N__23037));
    Odrv4 I__4818 (
            .O(N__23037),
            .I(\this_sprites_ram.mem_out_bus3_1 ));
    InMux I__4817 (
            .O(N__23034),
            .I(N__23031));
    LocalMux I__4816 (
            .O(N__23031),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ));
    InMux I__4815 (
            .O(N__23028),
            .I(N__23025));
    LocalMux I__4814 (
            .O(N__23025),
            .I(N__23022));
    Span12Mux_v I__4813 (
            .O(N__23022),
            .I(N__23019));
    Span12Mux_h I__4812 (
            .O(N__23019),
            .I(N__23016));
    Odrv12 I__4811 (
            .O(N__23016),
            .I(\this_sprites_ram.mem_out_bus4_3 ));
    InMux I__4810 (
            .O(N__23013),
            .I(N__23010));
    LocalMux I__4809 (
            .O(N__23010),
            .I(N__23007));
    Span4Mux_v I__4808 (
            .O(N__23007),
            .I(N__23004));
    Span4Mux_h I__4807 (
            .O(N__23004),
            .I(N__23001));
    Span4Mux_v I__4806 (
            .O(N__23001),
            .I(N__22998));
    Odrv4 I__4805 (
            .O(N__22998),
            .I(\this_sprites_ram.mem_out_bus0_3 ));
    InMux I__4804 (
            .O(N__22995),
            .I(N__22992));
    LocalMux I__4803 (
            .O(N__22992),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ));
    InMux I__4802 (
            .O(N__22989),
            .I(N__22985));
    InMux I__4801 (
            .O(N__22988),
            .I(N__22982));
    LocalMux I__4800 (
            .O(N__22985),
            .I(N__22979));
    LocalMux I__4799 (
            .O(N__22982),
            .I(N__22975));
    Span4Mux_h I__4798 (
            .O(N__22979),
            .I(N__22972));
    InMux I__4797 (
            .O(N__22978),
            .I(N__22969));
    Span4Mux_h I__4796 (
            .O(N__22975),
            .I(N__22966));
    Span4Mux_v I__4795 (
            .O(N__22972),
            .I(N__22963));
    LocalMux I__4794 (
            .O(N__22969),
            .I(N__22960));
    Span4Mux_v I__4793 (
            .O(N__22966),
            .I(N__22957));
    Sp12to4 I__4792 (
            .O(N__22963),
            .I(N__22949));
    Span12Mux_v I__4791 (
            .O(N__22960),
            .I(N__22949));
    Sp12to4 I__4790 (
            .O(N__22957),
            .I(N__22949));
    InMux I__4789 (
            .O(N__22956),
            .I(N__22946));
    Odrv12 I__4788 (
            .O(N__22949),
            .I(this_vga_signals_vvisibility));
    LocalMux I__4787 (
            .O(N__22946),
            .I(this_vga_signals_vvisibility));
    IoInMux I__4786 (
            .O(N__22941),
            .I(N__22938));
    LocalMux I__4785 (
            .O(N__22938),
            .I(N__22935));
    Span4Mux_s2_h I__4784 (
            .O(N__22935),
            .I(N__22932));
    Span4Mux_v I__4783 (
            .O(N__22932),
            .I(N__22927));
    InMux I__4782 (
            .O(N__22931),
            .I(N__22924));
    CascadeMux I__4781 (
            .O(N__22930),
            .I(N__22920));
    Sp12to4 I__4780 (
            .O(N__22927),
            .I(N__22917));
    LocalMux I__4779 (
            .O(N__22924),
            .I(N__22914));
    InMux I__4778 (
            .O(N__22923),
            .I(N__22911));
    InMux I__4777 (
            .O(N__22920),
            .I(N__22908));
    Span12Mux_h I__4776 (
            .O(N__22917),
            .I(N__22905));
    Span12Mux_v I__4775 (
            .O(N__22914),
            .I(N__22902));
    LocalMux I__4774 (
            .O(N__22911),
            .I(N__22898));
    LocalMux I__4773 (
            .O(N__22908),
            .I(N__22895));
    Span12Mux_v I__4772 (
            .O(N__22905),
            .I(N__22890));
    Span12Mux_h I__4771 (
            .O(N__22902),
            .I(N__22890));
    InMux I__4770 (
            .O(N__22901),
            .I(N__22887));
    Span12Mux_s7_h I__4769 (
            .O(N__22898),
            .I(N__22882));
    Span12Mux_v I__4768 (
            .O(N__22895),
            .I(N__22882));
    Odrv12 I__4767 (
            .O(N__22890),
            .I(dma_0));
    LocalMux I__4766 (
            .O(N__22887),
            .I(dma_0));
    Odrv12 I__4765 (
            .O(N__22882),
            .I(dma_0));
    CascadeMux I__4764 (
            .O(N__22875),
            .I(\this_ppu.N_150_cascade_ ));
    InMux I__4763 (
            .O(N__22872),
            .I(N__22867));
    InMux I__4762 (
            .O(N__22871),
            .I(N__22864));
    InMux I__4761 (
            .O(N__22870),
            .I(N__22855));
    LocalMux I__4760 (
            .O(N__22867),
            .I(N__22850));
    LocalMux I__4759 (
            .O(N__22864),
            .I(N__22850));
    InMux I__4758 (
            .O(N__22863),
            .I(N__22839));
    InMux I__4757 (
            .O(N__22862),
            .I(N__22839));
    InMux I__4756 (
            .O(N__22861),
            .I(N__22839));
    InMux I__4755 (
            .O(N__22860),
            .I(N__22839));
    InMux I__4754 (
            .O(N__22859),
            .I(N__22839));
    IoInMux I__4753 (
            .O(N__22858),
            .I(N__22836));
    LocalMux I__4752 (
            .O(N__22855),
            .I(N__22833));
    Span4Mux_v I__4751 (
            .O(N__22850),
            .I(N__22830));
    LocalMux I__4750 (
            .O(N__22839),
            .I(N__22827));
    LocalMux I__4749 (
            .O(N__22836),
            .I(N__22823));
    Span4Mux_h I__4748 (
            .O(N__22833),
            .I(N__22820));
    Span4Mux_h I__4747 (
            .O(N__22830),
            .I(N__22815));
    Span4Mux_h I__4746 (
            .O(N__22827),
            .I(N__22815));
    InMux I__4745 (
            .O(N__22826),
            .I(N__22812));
    Span12Mux_s5_v I__4744 (
            .O(N__22823),
            .I(N__22809));
    Odrv4 I__4743 (
            .O(N__22820),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__4742 (
            .O(N__22815),
            .I(M_this_reset_cond_out_0));
    LocalMux I__4741 (
            .O(N__22812),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__4740 (
            .O(N__22809),
            .I(M_this_reset_cond_out_0));
    CascadeMux I__4739 (
            .O(N__22800),
            .I(N__22795));
    CascadeMux I__4738 (
            .O(N__22799),
            .I(N__22790));
    CascadeMux I__4737 (
            .O(N__22798),
            .I(N__22787));
    InMux I__4736 (
            .O(N__22795),
            .I(N__22782));
    CascadeMux I__4735 (
            .O(N__22794),
            .I(N__22779));
    CascadeMux I__4734 (
            .O(N__22793),
            .I(N__22776));
    InMux I__4733 (
            .O(N__22790),
            .I(N__22767));
    InMux I__4732 (
            .O(N__22787),
            .I(N__22764));
    CascadeMux I__4731 (
            .O(N__22786),
            .I(N__22761));
    CascadeMux I__4730 (
            .O(N__22785),
            .I(N__22758));
    LocalMux I__4729 (
            .O(N__22782),
            .I(N__22754));
    InMux I__4728 (
            .O(N__22779),
            .I(N__22751));
    InMux I__4727 (
            .O(N__22776),
            .I(N__22748));
    CascadeMux I__4726 (
            .O(N__22775),
            .I(N__22745));
    CascadeMux I__4725 (
            .O(N__22774),
            .I(N__22742));
    CascadeMux I__4724 (
            .O(N__22773),
            .I(N__22737));
    CascadeMux I__4723 (
            .O(N__22772),
            .I(N__22734));
    CascadeMux I__4722 (
            .O(N__22771),
            .I(N__22731));
    CascadeMux I__4721 (
            .O(N__22770),
            .I(N__22728));
    LocalMux I__4720 (
            .O(N__22767),
            .I(N__22723));
    LocalMux I__4719 (
            .O(N__22764),
            .I(N__22723));
    InMux I__4718 (
            .O(N__22761),
            .I(N__22720));
    InMux I__4717 (
            .O(N__22758),
            .I(N__22717));
    CascadeMux I__4716 (
            .O(N__22757),
            .I(N__22714));
    Span4Mux_v I__4715 (
            .O(N__22754),
            .I(N__22707));
    LocalMux I__4714 (
            .O(N__22751),
            .I(N__22707));
    LocalMux I__4713 (
            .O(N__22748),
            .I(N__22707));
    InMux I__4712 (
            .O(N__22745),
            .I(N__22704));
    InMux I__4711 (
            .O(N__22742),
            .I(N__22701));
    CascadeMux I__4710 (
            .O(N__22741),
            .I(N__22698));
    CascadeMux I__4709 (
            .O(N__22740),
            .I(N__22695));
    InMux I__4708 (
            .O(N__22737),
            .I(N__22692));
    InMux I__4707 (
            .O(N__22734),
            .I(N__22689));
    InMux I__4706 (
            .O(N__22731),
            .I(N__22686));
    InMux I__4705 (
            .O(N__22728),
            .I(N__22683));
    Span4Mux_v I__4704 (
            .O(N__22723),
            .I(N__22676));
    LocalMux I__4703 (
            .O(N__22720),
            .I(N__22676));
    LocalMux I__4702 (
            .O(N__22717),
            .I(N__22676));
    InMux I__4701 (
            .O(N__22714),
            .I(N__22673));
    Span4Mux_v I__4700 (
            .O(N__22707),
            .I(N__22666));
    LocalMux I__4699 (
            .O(N__22704),
            .I(N__22666));
    LocalMux I__4698 (
            .O(N__22701),
            .I(N__22666));
    InMux I__4697 (
            .O(N__22698),
            .I(N__22663));
    InMux I__4696 (
            .O(N__22695),
            .I(N__22660));
    LocalMux I__4695 (
            .O(N__22692),
            .I(N__22653));
    LocalMux I__4694 (
            .O(N__22689),
            .I(N__22653));
    LocalMux I__4693 (
            .O(N__22686),
            .I(N__22653));
    LocalMux I__4692 (
            .O(N__22683),
            .I(N__22650));
    Span4Mux_v I__4691 (
            .O(N__22676),
            .I(N__22645));
    LocalMux I__4690 (
            .O(N__22673),
            .I(N__22645));
    Span4Mux_v I__4689 (
            .O(N__22666),
            .I(N__22640));
    LocalMux I__4688 (
            .O(N__22663),
            .I(N__22640));
    LocalMux I__4687 (
            .O(N__22660),
            .I(N__22637));
    Span12Mux_v I__4686 (
            .O(N__22653),
            .I(N__22632));
    Span12Mux_v I__4685 (
            .O(N__22650),
            .I(N__22632));
    Span4Mux_v I__4684 (
            .O(N__22645),
            .I(N__22627));
    Span4Mux_v I__4683 (
            .O(N__22640),
            .I(N__22627));
    Span12Mux_h I__4682 (
            .O(N__22637),
            .I(N__22622));
    Span12Mux_h I__4681 (
            .O(N__22632),
            .I(N__22622));
    Span4Mux_h I__4680 (
            .O(N__22627),
            .I(N__22619));
    Odrv12 I__4679 (
            .O(N__22622),
            .I(M_this_ppu_sprites_addr_2));
    Odrv4 I__4678 (
            .O(N__22619),
            .I(M_this_ppu_sprites_addr_2));
    CEMux I__4677 (
            .O(N__22614),
            .I(N__22611));
    LocalMux I__4676 (
            .O(N__22611),
            .I(N__22608));
    Span12Mux_h I__4675 (
            .O(N__22608),
            .I(N__22602));
    InMux I__4674 (
            .O(N__22607),
            .I(N__22597));
    InMux I__4673 (
            .O(N__22606),
            .I(N__22597));
    InMux I__4672 (
            .O(N__22605),
            .I(N__22594));
    Odrv12 I__4671 (
            .O(N__22602),
            .I(M_this_ppu_vram_en_0));
    LocalMux I__4670 (
            .O(N__22597),
            .I(M_this_ppu_vram_en_0));
    LocalMux I__4669 (
            .O(N__22594),
            .I(M_this_ppu_vram_en_0));
    InMux I__4668 (
            .O(N__22587),
            .I(N__22584));
    LocalMux I__4667 (
            .O(N__22584),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9 ));
    CascadeMux I__4666 (
            .O(N__22581),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_9_cascade_ ));
    InMux I__4665 (
            .O(N__22578),
            .I(N__22575));
    LocalMux I__4664 (
            .O(N__22575),
            .I(un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0));
    CascadeMux I__4663 (
            .O(N__22572),
            .I(N__22565));
    CascadeMux I__4662 (
            .O(N__22571),
            .I(N__22562));
    CascadeMux I__4661 (
            .O(N__22570),
            .I(N__22555));
    CascadeMux I__4660 (
            .O(N__22569),
            .I(N__22549));
    CascadeMux I__4659 (
            .O(N__22568),
            .I(N__22545));
    InMux I__4658 (
            .O(N__22565),
            .I(N__22542));
    InMux I__4657 (
            .O(N__22562),
            .I(N__22539));
    CascadeMux I__4656 (
            .O(N__22561),
            .I(N__22536));
    CascadeMux I__4655 (
            .O(N__22560),
            .I(N__22533));
    CascadeMux I__4654 (
            .O(N__22559),
            .I(N__22530));
    CascadeMux I__4653 (
            .O(N__22558),
            .I(N__22527));
    InMux I__4652 (
            .O(N__22555),
            .I(N__22524));
    CascadeMux I__4651 (
            .O(N__22554),
            .I(N__22521));
    CascadeMux I__4650 (
            .O(N__22553),
            .I(N__22517));
    CascadeMux I__4649 (
            .O(N__22552),
            .I(N__22514));
    InMux I__4648 (
            .O(N__22549),
            .I(N__22511));
    CascadeMux I__4647 (
            .O(N__22548),
            .I(N__22508));
    InMux I__4646 (
            .O(N__22545),
            .I(N__22505));
    LocalMux I__4645 (
            .O(N__22542),
            .I(N__22500));
    LocalMux I__4644 (
            .O(N__22539),
            .I(N__22500));
    InMux I__4643 (
            .O(N__22536),
            .I(N__22497));
    InMux I__4642 (
            .O(N__22533),
            .I(N__22494));
    InMux I__4641 (
            .O(N__22530),
            .I(N__22491));
    InMux I__4640 (
            .O(N__22527),
            .I(N__22488));
    LocalMux I__4639 (
            .O(N__22524),
            .I(N__22485));
    InMux I__4638 (
            .O(N__22521),
            .I(N__22482));
    CascadeMux I__4637 (
            .O(N__22520),
            .I(N__22479));
    InMux I__4636 (
            .O(N__22517),
            .I(N__22475));
    InMux I__4635 (
            .O(N__22514),
            .I(N__22472));
    LocalMux I__4634 (
            .O(N__22511),
            .I(N__22469));
    InMux I__4633 (
            .O(N__22508),
            .I(N__22466));
    LocalMux I__4632 (
            .O(N__22505),
            .I(N__22459));
    Span4Mux_v I__4631 (
            .O(N__22500),
            .I(N__22459));
    LocalMux I__4630 (
            .O(N__22497),
            .I(N__22459));
    LocalMux I__4629 (
            .O(N__22494),
            .I(N__22454));
    LocalMux I__4628 (
            .O(N__22491),
            .I(N__22454));
    LocalMux I__4627 (
            .O(N__22488),
            .I(N__22451));
    Span4Mux_v I__4626 (
            .O(N__22485),
            .I(N__22446));
    LocalMux I__4625 (
            .O(N__22482),
            .I(N__22446));
    InMux I__4624 (
            .O(N__22479),
            .I(N__22443));
    CascadeMux I__4623 (
            .O(N__22478),
            .I(N__22439));
    LocalMux I__4622 (
            .O(N__22475),
            .I(N__22436));
    LocalMux I__4621 (
            .O(N__22472),
            .I(N__22433));
    Span4Mux_h I__4620 (
            .O(N__22469),
            .I(N__22430));
    LocalMux I__4619 (
            .O(N__22466),
            .I(N__22427));
    Span4Mux_v I__4618 (
            .O(N__22459),
            .I(N__22422));
    Span4Mux_v I__4617 (
            .O(N__22454),
            .I(N__22422));
    Span4Mux_h I__4616 (
            .O(N__22451),
            .I(N__22419));
    Span4Mux_v I__4615 (
            .O(N__22446),
            .I(N__22413));
    LocalMux I__4614 (
            .O(N__22443),
            .I(N__22413));
    CascadeMux I__4613 (
            .O(N__22442),
            .I(N__22410));
    InMux I__4612 (
            .O(N__22439),
            .I(N__22407));
    Span4Mux_h I__4611 (
            .O(N__22436),
            .I(N__22404));
    Span4Mux_h I__4610 (
            .O(N__22433),
            .I(N__22399));
    Span4Mux_v I__4609 (
            .O(N__22430),
            .I(N__22399));
    Span4Mux_h I__4608 (
            .O(N__22427),
            .I(N__22396));
    Sp12to4 I__4607 (
            .O(N__22422),
            .I(N__22393));
    Span4Mux_h I__4606 (
            .O(N__22419),
            .I(N__22390));
    InMux I__4605 (
            .O(N__22418),
            .I(N__22387));
    Span4Mux_h I__4604 (
            .O(N__22413),
            .I(N__22384));
    InMux I__4603 (
            .O(N__22410),
            .I(N__22381));
    LocalMux I__4602 (
            .O(N__22407),
            .I(N__22378));
    Span4Mux_h I__4601 (
            .O(N__22404),
            .I(N__22374));
    Span4Mux_h I__4600 (
            .O(N__22399),
            .I(N__22370));
    Span4Mux_h I__4599 (
            .O(N__22396),
            .I(N__22367));
    Span12Mux_h I__4598 (
            .O(N__22393),
            .I(N__22364));
    Sp12to4 I__4597 (
            .O(N__22390),
            .I(N__22361));
    LocalMux I__4596 (
            .O(N__22387),
            .I(N__22356));
    Span4Mux_v I__4595 (
            .O(N__22384),
            .I(N__22356));
    LocalMux I__4594 (
            .O(N__22381),
            .I(N__22351));
    Span12Mux_h I__4593 (
            .O(N__22378),
            .I(N__22351));
    InMux I__4592 (
            .O(N__22377),
            .I(N__22348));
    Span4Mux_h I__4591 (
            .O(N__22374),
            .I(N__22345));
    InMux I__4590 (
            .O(N__22373),
            .I(N__22342));
    Span4Mux_h I__4589 (
            .O(N__22370),
            .I(N__22339));
    Sp12to4 I__4588 (
            .O(N__22367),
            .I(N__22334));
    Span12Mux_v I__4587 (
            .O(N__22364),
            .I(N__22334));
    Span12Mux_v I__4586 (
            .O(N__22361),
            .I(N__22331));
    Odrv4 I__4585 (
            .O(N__22356),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv12 I__4584 (
            .O(N__22351),
            .I(M_this_sprites_address_qZ0Z_9));
    LocalMux I__4583 (
            .O(N__22348),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv4 I__4582 (
            .O(N__22345),
            .I(M_this_sprites_address_qZ0Z_9));
    LocalMux I__4581 (
            .O(N__22342),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv4 I__4580 (
            .O(N__22339),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv12 I__4579 (
            .O(N__22334),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv12 I__4578 (
            .O(N__22331),
            .I(M_this_sprites_address_qZ0Z_9));
    InMux I__4577 (
            .O(N__22314),
            .I(N__22311));
    LocalMux I__4576 (
            .O(N__22311),
            .I(N__22308));
    Odrv12 I__4575 (
            .O(N__22308),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2 ));
    CascadeMux I__4574 (
            .O(N__22305),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_2_cascade_ ));
    InMux I__4573 (
            .O(N__22302),
            .I(N__22299));
    LocalMux I__4572 (
            .O(N__22299),
            .I(N__22296));
    Odrv4 I__4571 (
            .O(N__22296),
            .I(un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0));
    CascadeMux I__4570 (
            .O(N__22293),
            .I(N__22290));
    InMux I__4569 (
            .O(N__22290),
            .I(N__22286));
    CascadeMux I__4568 (
            .O(N__22289),
            .I(N__22283));
    LocalMux I__4567 (
            .O(N__22286),
            .I(N__22278));
    InMux I__4566 (
            .O(N__22283),
            .I(N__22275));
    CascadeMux I__4565 (
            .O(N__22282),
            .I(N__22272));
    CascadeMux I__4564 (
            .O(N__22281),
            .I(N__22268));
    Span4Mux_v I__4563 (
            .O(N__22278),
            .I(N__22260));
    LocalMux I__4562 (
            .O(N__22275),
            .I(N__22260));
    InMux I__4561 (
            .O(N__22272),
            .I(N__22257));
    CascadeMux I__4560 (
            .O(N__22271),
            .I(N__22254));
    InMux I__4559 (
            .O(N__22268),
            .I(N__22250));
    CascadeMux I__4558 (
            .O(N__22267),
            .I(N__22247));
    CascadeMux I__4557 (
            .O(N__22266),
            .I(N__22243));
    CascadeMux I__4556 (
            .O(N__22265),
            .I(N__22238));
    Span4Mux_h I__4555 (
            .O(N__22260),
            .I(N__22232));
    LocalMux I__4554 (
            .O(N__22257),
            .I(N__22232));
    InMux I__4553 (
            .O(N__22254),
            .I(N__22229));
    CascadeMux I__4552 (
            .O(N__22253),
            .I(N__22224));
    LocalMux I__4551 (
            .O(N__22250),
            .I(N__22221));
    InMux I__4550 (
            .O(N__22247),
            .I(N__22218));
    CascadeMux I__4549 (
            .O(N__22246),
            .I(N__22215));
    InMux I__4548 (
            .O(N__22243),
            .I(N__22212));
    CascadeMux I__4547 (
            .O(N__22242),
            .I(N__22209));
    CascadeMux I__4546 (
            .O(N__22241),
            .I(N__22206));
    InMux I__4545 (
            .O(N__22238),
            .I(N__22203));
    CascadeMux I__4544 (
            .O(N__22237),
            .I(N__22200));
    Span4Mux_v I__4543 (
            .O(N__22232),
            .I(N__22195));
    LocalMux I__4542 (
            .O(N__22229),
            .I(N__22195));
    CascadeMux I__4541 (
            .O(N__22228),
            .I(N__22192));
    CascadeMux I__4540 (
            .O(N__22227),
            .I(N__22189));
    InMux I__4539 (
            .O(N__22224),
            .I(N__22186));
    Span4Mux_h I__4538 (
            .O(N__22221),
            .I(N__22180));
    LocalMux I__4537 (
            .O(N__22218),
            .I(N__22180));
    InMux I__4536 (
            .O(N__22215),
            .I(N__22177));
    LocalMux I__4535 (
            .O(N__22212),
            .I(N__22174));
    InMux I__4534 (
            .O(N__22209),
            .I(N__22171));
    InMux I__4533 (
            .O(N__22206),
            .I(N__22168));
    LocalMux I__4532 (
            .O(N__22203),
            .I(N__22165));
    InMux I__4531 (
            .O(N__22200),
            .I(N__22162));
    Span4Mux_v I__4530 (
            .O(N__22195),
            .I(N__22159));
    InMux I__4529 (
            .O(N__22192),
            .I(N__22156));
    InMux I__4528 (
            .O(N__22189),
            .I(N__22153));
    LocalMux I__4527 (
            .O(N__22186),
            .I(N__22150));
    CascadeMux I__4526 (
            .O(N__22185),
            .I(N__22147));
    Span4Mux_v I__4525 (
            .O(N__22180),
            .I(N__22144));
    LocalMux I__4524 (
            .O(N__22177),
            .I(N__22141));
    Span4Mux_v I__4523 (
            .O(N__22174),
            .I(N__22134));
    LocalMux I__4522 (
            .O(N__22171),
            .I(N__22134));
    LocalMux I__4521 (
            .O(N__22168),
            .I(N__22134));
    Span12Mux_h I__4520 (
            .O(N__22165),
            .I(N__22129));
    LocalMux I__4519 (
            .O(N__22162),
            .I(N__22126));
    Sp12to4 I__4518 (
            .O(N__22159),
            .I(N__22121));
    LocalMux I__4517 (
            .O(N__22156),
            .I(N__22121));
    LocalMux I__4516 (
            .O(N__22153),
            .I(N__22118));
    Span12Mux_h I__4515 (
            .O(N__22150),
            .I(N__22115));
    InMux I__4514 (
            .O(N__22147),
            .I(N__22112));
    Span4Mux_h I__4513 (
            .O(N__22144),
            .I(N__22108));
    Span4Mux_v I__4512 (
            .O(N__22141),
            .I(N__22103));
    Span4Mux_v I__4511 (
            .O(N__22134),
            .I(N__22103));
    InMux I__4510 (
            .O(N__22133),
            .I(N__22100));
    InMux I__4509 (
            .O(N__22132),
            .I(N__22097));
    Span12Mux_v I__4508 (
            .O(N__22129),
            .I(N__22090));
    Span12Mux_h I__4507 (
            .O(N__22126),
            .I(N__22090));
    Span12Mux_h I__4506 (
            .O(N__22121),
            .I(N__22090));
    Span12Mux_s10_h I__4505 (
            .O(N__22118),
            .I(N__22087));
    Span12Mux_v I__4504 (
            .O(N__22115),
            .I(N__22082));
    LocalMux I__4503 (
            .O(N__22112),
            .I(N__22082));
    InMux I__4502 (
            .O(N__22111),
            .I(N__22079));
    Span4Mux_h I__4501 (
            .O(N__22108),
            .I(N__22072));
    Span4Mux_h I__4500 (
            .O(N__22103),
            .I(N__22072));
    LocalMux I__4499 (
            .O(N__22100),
            .I(N__22072));
    LocalMux I__4498 (
            .O(N__22097),
            .I(N__22069));
    Odrv12 I__4497 (
            .O(N__22090),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv12 I__4496 (
            .O(N__22087),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv12 I__4495 (
            .O(N__22082),
            .I(M_this_sprites_address_qZ0Z_2));
    LocalMux I__4494 (
            .O(N__22079),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv4 I__4493 (
            .O(N__22072),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv4 I__4492 (
            .O(N__22069),
            .I(M_this_sprites_address_qZ0Z_2));
    CascadeMux I__4491 (
            .O(N__22056),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3_cascade_ ));
    InMux I__4490 (
            .O(N__22053),
            .I(N__22050));
    LocalMux I__4489 (
            .O(N__22050),
            .I(N__22047));
    Odrv4 I__4488 (
            .O(N__22047),
            .I(un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0));
    CascadeMux I__4487 (
            .O(N__22044),
            .I(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_ ));
    InMux I__4486 (
            .O(N__22041),
            .I(N__22038));
    LocalMux I__4485 (
            .O(N__22038),
            .I(N__22035));
    Odrv4 I__4484 (
            .O(N__22035),
            .I(un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0));
    CascadeMux I__4483 (
            .O(N__22032),
            .I(N__22028));
    CascadeMux I__4482 (
            .O(N__22031),
            .I(N__22025));
    InMux I__4481 (
            .O(N__22028),
            .I(N__22018));
    InMux I__4480 (
            .O(N__22025),
            .I(N__22015));
    CascadeMux I__4479 (
            .O(N__22024),
            .I(N__22012));
    CascadeMux I__4478 (
            .O(N__22023),
            .I(N__22009));
    CascadeMux I__4477 (
            .O(N__22022),
            .I(N__22004));
    CascadeMux I__4476 (
            .O(N__22021),
            .I(N__22001));
    LocalMux I__4475 (
            .O(N__22018),
            .I(N__21995));
    LocalMux I__4474 (
            .O(N__22015),
            .I(N__21995));
    InMux I__4473 (
            .O(N__22012),
            .I(N__21992));
    InMux I__4472 (
            .O(N__22009),
            .I(N__21989));
    CascadeMux I__4471 (
            .O(N__22008),
            .I(N__21986));
    CascadeMux I__4470 (
            .O(N__22007),
            .I(N__21983));
    InMux I__4469 (
            .O(N__22004),
            .I(N__21979));
    InMux I__4468 (
            .O(N__22001),
            .I(N__21976));
    CascadeMux I__4467 (
            .O(N__22000),
            .I(N__21973));
    Span4Mux_v I__4466 (
            .O(N__21995),
            .I(N__21965));
    LocalMux I__4465 (
            .O(N__21992),
            .I(N__21965));
    LocalMux I__4464 (
            .O(N__21989),
            .I(N__21965));
    InMux I__4463 (
            .O(N__21986),
            .I(N__21962));
    InMux I__4462 (
            .O(N__21983),
            .I(N__21959));
    CascadeMux I__4461 (
            .O(N__21982),
            .I(N__21956));
    LocalMux I__4460 (
            .O(N__21979),
            .I(N__21949));
    LocalMux I__4459 (
            .O(N__21976),
            .I(N__21949));
    InMux I__4458 (
            .O(N__21973),
            .I(N__21946));
    CascadeMux I__4457 (
            .O(N__21972),
            .I(N__21943));
    Span4Mux_v I__4456 (
            .O(N__21965),
            .I(N__21936));
    LocalMux I__4455 (
            .O(N__21962),
            .I(N__21936));
    LocalMux I__4454 (
            .O(N__21959),
            .I(N__21936));
    InMux I__4453 (
            .O(N__21956),
            .I(N__21933));
    CascadeMux I__4452 (
            .O(N__21955),
            .I(N__21928));
    CascadeMux I__4451 (
            .O(N__21954),
            .I(N__21924));
    Span4Mux_v I__4450 (
            .O(N__21949),
            .I(N__21919));
    LocalMux I__4449 (
            .O(N__21946),
            .I(N__21919));
    InMux I__4448 (
            .O(N__21943),
            .I(N__21916));
    Span4Mux_v I__4447 (
            .O(N__21936),
            .I(N__21911));
    LocalMux I__4446 (
            .O(N__21933),
            .I(N__21911));
    CascadeMux I__4445 (
            .O(N__21932),
            .I(N__21908));
    CascadeMux I__4444 (
            .O(N__21931),
            .I(N__21905));
    InMux I__4443 (
            .O(N__21928),
            .I(N__21902));
    CascadeMux I__4442 (
            .O(N__21927),
            .I(N__21899));
    InMux I__4441 (
            .O(N__21924),
            .I(N__21896));
    Span4Mux_v I__4440 (
            .O(N__21919),
            .I(N__21891));
    LocalMux I__4439 (
            .O(N__21916),
            .I(N__21891));
    Span4Mux_v I__4438 (
            .O(N__21911),
            .I(N__21888));
    InMux I__4437 (
            .O(N__21908),
            .I(N__21885));
    InMux I__4436 (
            .O(N__21905),
            .I(N__21882));
    LocalMux I__4435 (
            .O(N__21902),
            .I(N__21879));
    InMux I__4434 (
            .O(N__21899),
            .I(N__21876));
    LocalMux I__4433 (
            .O(N__21896),
            .I(N__21873));
    Span4Mux_v I__4432 (
            .O(N__21891),
            .I(N__21870));
    Sp12to4 I__4431 (
            .O(N__21888),
            .I(N__21867));
    LocalMux I__4430 (
            .O(N__21885),
            .I(N__21864));
    LocalMux I__4429 (
            .O(N__21882),
            .I(N__21861));
    Span4Mux_v I__4428 (
            .O(N__21879),
            .I(N__21855));
    LocalMux I__4427 (
            .O(N__21876),
            .I(N__21855));
    Span4Mux_s3_v I__4426 (
            .O(N__21873),
            .I(N__21852));
    Sp12to4 I__4425 (
            .O(N__21870),
            .I(N__21849));
    Span12Mux_h I__4424 (
            .O(N__21867),
            .I(N__21846));
    Span4Mux_h I__4423 (
            .O(N__21864),
            .I(N__21843));
    Span4Mux_h I__4422 (
            .O(N__21861),
            .I(N__21840));
    InMux I__4421 (
            .O(N__21860),
            .I(N__21835));
    Span4Mux_v I__4420 (
            .O(N__21855),
            .I(N__21830));
    Span4Mux_v I__4419 (
            .O(N__21852),
            .I(N__21830));
    Span12Mux_h I__4418 (
            .O(N__21849),
            .I(N__21825));
    Span12Mux_v I__4417 (
            .O(N__21846),
            .I(N__21825));
    Span4Mux_h I__4416 (
            .O(N__21843),
            .I(N__21820));
    Span4Mux_h I__4415 (
            .O(N__21840),
            .I(N__21820));
    InMux I__4414 (
            .O(N__21839),
            .I(N__21815));
    InMux I__4413 (
            .O(N__21838),
            .I(N__21815));
    LocalMux I__4412 (
            .O(N__21835),
            .I(N__21812));
    Sp12to4 I__4411 (
            .O(N__21830),
            .I(N__21807));
    Span12Mux_v I__4410 (
            .O(N__21825),
            .I(N__21807));
    Odrv4 I__4409 (
            .O(N__21820),
            .I(M_this_sprites_address_qZ0Z_7));
    LocalMux I__4408 (
            .O(N__21815),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv4 I__4407 (
            .O(N__21812),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv12 I__4406 (
            .O(N__21807),
            .I(M_this_sprites_address_qZ0Z_7));
    InMux I__4405 (
            .O(N__21798),
            .I(N__21795));
    LocalMux I__4404 (
            .O(N__21795),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_7 ));
    InMux I__4403 (
            .O(N__21792),
            .I(N__21789));
    LocalMux I__4402 (
            .O(N__21789),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ));
    InMux I__4401 (
            .O(N__21786),
            .I(N__21783));
    LocalMux I__4400 (
            .O(N__21783),
            .I(N__21780));
    Span12Mux_v I__4399 (
            .O(N__21780),
            .I(N__21777));
    Span12Mux_h I__4398 (
            .O(N__21777),
            .I(N__21773));
    InMux I__4397 (
            .O(N__21776),
            .I(N__21770));
    Odrv12 I__4396 (
            .O(N__21773),
            .I(M_this_ppu_vram_data_1));
    LocalMux I__4395 (
            .O(N__21770),
            .I(M_this_ppu_vram_data_1));
    InMux I__4394 (
            .O(N__21765),
            .I(un1_M_this_sprites_address_q_cry_6));
    InMux I__4393 (
            .O(N__21762),
            .I(bfn_19_23_0_));
    InMux I__4392 (
            .O(N__21759),
            .I(un1_M_this_sprites_address_q_cry_8));
    InMux I__4391 (
            .O(N__21756),
            .I(un1_M_this_sprites_address_q_cry_9));
    InMux I__4390 (
            .O(N__21753),
            .I(un1_M_this_sprites_address_q_cry_10));
    InMux I__4389 (
            .O(N__21750),
            .I(un1_M_this_sprites_address_q_cry_11));
    InMux I__4388 (
            .O(N__21747),
            .I(un1_M_this_sprites_address_q_cry_12));
    InMux I__4387 (
            .O(N__21744),
            .I(N__21741));
    LocalMux I__4386 (
            .O(N__21741),
            .I(N__21738));
    Span4Mux_v I__4385 (
            .O(N__21738),
            .I(N__21735));
    Odrv4 I__4384 (
            .O(N__21735),
            .I(M_this_state_d25));
    InMux I__4383 (
            .O(N__21732),
            .I(N__21729));
    LocalMux I__4382 (
            .O(N__21729),
            .I(N__21724));
    InMux I__4381 (
            .O(N__21728),
            .I(N__21721));
    InMux I__4380 (
            .O(N__21727),
            .I(N__21718));
    Span12Mux_h I__4379 (
            .O(N__21724),
            .I(N__21711));
    LocalMux I__4378 (
            .O(N__21721),
            .I(N__21711));
    LocalMux I__4377 (
            .O(N__21718),
            .I(N__21711));
    Span12Mux_h I__4376 (
            .O(N__21711),
            .I(N__21707));
    InMux I__4375 (
            .O(N__21710),
            .I(N__21704));
    Odrv12 I__4374 (
            .O(N__21707),
            .I(port_rw_in));
    LocalMux I__4373 (
            .O(N__21704),
            .I(port_rw_in));
    IoInMux I__4372 (
            .O(N__21699),
            .I(N__21696));
    LocalMux I__4371 (
            .O(N__21696),
            .I(N__21693));
    Span4Mux_s3_h I__4370 (
            .O(N__21693),
            .I(N__21690));
    Sp12to4 I__4369 (
            .O(N__21690),
            .I(N__21686));
    InMux I__4368 (
            .O(N__21689),
            .I(N__21683));
    Span12Mux_v I__4367 (
            .O(N__21686),
            .I(N__21680));
    LocalMux I__4366 (
            .O(N__21683),
            .I(N__21675));
    Span12Mux_h I__4365 (
            .O(N__21680),
            .I(N__21672));
    InMux I__4364 (
            .O(N__21679),
            .I(N__21669));
    InMux I__4363 (
            .O(N__21678),
            .I(N__21666));
    Span4Mux_h I__4362 (
            .O(N__21675),
            .I(N__21663));
    Odrv12 I__4361 (
            .O(N__21672),
            .I(led_c_1));
    LocalMux I__4360 (
            .O(N__21669),
            .I(led_c_1));
    LocalMux I__4359 (
            .O(N__21666),
            .I(led_c_1));
    Odrv4 I__4358 (
            .O(N__21663),
            .I(led_c_1));
    CascadeMux I__4357 (
            .O(N__21654),
            .I(N__21651));
    InMux I__4356 (
            .O(N__21651),
            .I(N__21643));
    InMux I__4355 (
            .O(N__21650),
            .I(N__21643));
    InMux I__4354 (
            .O(N__21649),
            .I(N__21640));
    InMux I__4353 (
            .O(N__21648),
            .I(N__21636));
    LocalMux I__4352 (
            .O(N__21643),
            .I(N__21629));
    LocalMux I__4351 (
            .O(N__21640),
            .I(N__21629));
    InMux I__4350 (
            .O(N__21639),
            .I(N__21626));
    LocalMux I__4349 (
            .O(N__21636),
            .I(N__21623));
    InMux I__4348 (
            .O(N__21635),
            .I(N__21618));
    InMux I__4347 (
            .O(N__21634),
            .I(N__21618));
    Span4Mux_v I__4346 (
            .O(N__21629),
            .I(N__21613));
    LocalMux I__4345 (
            .O(N__21626),
            .I(N__21613));
    Odrv4 I__4344 (
            .O(N__21623),
            .I(N_459_0));
    LocalMux I__4343 (
            .O(N__21618),
            .I(N_459_0));
    Odrv4 I__4342 (
            .O(N__21613),
            .I(N_459_0));
    CascadeMux I__4341 (
            .O(N__21606),
            .I(N__21602));
    InMux I__4340 (
            .O(N__21605),
            .I(N__21599));
    InMux I__4339 (
            .O(N__21602),
            .I(N__21596));
    LocalMux I__4338 (
            .O(N__21599),
            .I(un1_M_this_state_q_12_0));
    LocalMux I__4337 (
            .O(N__21596),
            .I(un1_M_this_state_q_12_0));
    InMux I__4336 (
            .O(N__21591),
            .I(un1_M_this_sprites_address_q_cry_0));
    InMux I__4335 (
            .O(N__21588),
            .I(un1_M_this_sprites_address_q_cry_1));
    InMux I__4334 (
            .O(N__21585),
            .I(un1_M_this_sprites_address_q_cry_2));
    InMux I__4333 (
            .O(N__21582),
            .I(un1_M_this_sprites_address_q_cry_3));
    CascadeMux I__4332 (
            .O(N__21579),
            .I(N__21573));
    CascadeMux I__4331 (
            .O(N__21578),
            .I(N__21567));
    CascadeMux I__4330 (
            .O(N__21577),
            .I(N__21560));
    CascadeMux I__4329 (
            .O(N__21576),
            .I(N__21557));
    InMux I__4328 (
            .O(N__21573),
            .I(N__21554));
    CascadeMux I__4327 (
            .O(N__21572),
            .I(N__21551));
    CascadeMux I__4326 (
            .O(N__21571),
            .I(N__21545));
    CascadeMux I__4325 (
            .O(N__21570),
            .I(N__21542));
    InMux I__4324 (
            .O(N__21567),
            .I(N__21539));
    CascadeMux I__4323 (
            .O(N__21566),
            .I(N__21534));
    CascadeMux I__4322 (
            .O(N__21565),
            .I(N__21531));
    CascadeMux I__4321 (
            .O(N__21564),
            .I(N__21528));
    CascadeMux I__4320 (
            .O(N__21563),
            .I(N__21525));
    InMux I__4319 (
            .O(N__21560),
            .I(N__21522));
    InMux I__4318 (
            .O(N__21557),
            .I(N__21519));
    LocalMux I__4317 (
            .O(N__21554),
            .I(N__21516));
    InMux I__4316 (
            .O(N__21551),
            .I(N__21513));
    CascadeMux I__4315 (
            .O(N__21550),
            .I(N__21510));
    CascadeMux I__4314 (
            .O(N__21549),
            .I(N__21507));
    CascadeMux I__4313 (
            .O(N__21548),
            .I(N__21504));
    InMux I__4312 (
            .O(N__21545),
            .I(N__21501));
    InMux I__4311 (
            .O(N__21542),
            .I(N__21498));
    LocalMux I__4310 (
            .O(N__21539),
            .I(N__21495));
    CascadeMux I__4309 (
            .O(N__21538),
            .I(N__21492));
    CascadeMux I__4308 (
            .O(N__21537),
            .I(N__21489));
    InMux I__4307 (
            .O(N__21534),
            .I(N__21486));
    InMux I__4306 (
            .O(N__21531),
            .I(N__21483));
    InMux I__4305 (
            .O(N__21528),
            .I(N__21480));
    InMux I__4304 (
            .O(N__21525),
            .I(N__21477));
    LocalMux I__4303 (
            .O(N__21522),
            .I(N__21470));
    LocalMux I__4302 (
            .O(N__21519),
            .I(N__21470));
    Span4Mux_v I__4301 (
            .O(N__21516),
            .I(N__21470));
    LocalMux I__4300 (
            .O(N__21513),
            .I(N__21467));
    InMux I__4299 (
            .O(N__21510),
            .I(N__21464));
    InMux I__4298 (
            .O(N__21507),
            .I(N__21461));
    InMux I__4297 (
            .O(N__21504),
            .I(N__21458));
    LocalMux I__4296 (
            .O(N__21501),
            .I(N__21453));
    LocalMux I__4295 (
            .O(N__21498),
            .I(N__21453));
    Span4Mux_v I__4294 (
            .O(N__21495),
            .I(N__21450));
    InMux I__4293 (
            .O(N__21492),
            .I(N__21447));
    InMux I__4292 (
            .O(N__21489),
            .I(N__21444));
    LocalMux I__4291 (
            .O(N__21486),
            .I(N__21441));
    LocalMux I__4290 (
            .O(N__21483),
            .I(N__21434));
    LocalMux I__4289 (
            .O(N__21480),
            .I(N__21434));
    LocalMux I__4288 (
            .O(N__21477),
            .I(N__21434));
    Span4Mux_v I__4287 (
            .O(N__21470),
            .I(N__21429));
    Span4Mux_v I__4286 (
            .O(N__21467),
            .I(N__21429));
    LocalMux I__4285 (
            .O(N__21464),
            .I(N__21424));
    LocalMux I__4284 (
            .O(N__21461),
            .I(N__21419));
    LocalMux I__4283 (
            .O(N__21458),
            .I(N__21419));
    Span4Mux_v I__4282 (
            .O(N__21453),
            .I(N__21414));
    Span4Mux_v I__4281 (
            .O(N__21450),
            .I(N__21414));
    LocalMux I__4280 (
            .O(N__21447),
            .I(N__21405));
    LocalMux I__4279 (
            .O(N__21444),
            .I(N__21405));
    Span12Mux_s7_h I__4278 (
            .O(N__21441),
            .I(N__21405));
    Span12Mux_s9_v I__4277 (
            .O(N__21434),
            .I(N__21405));
    Sp12to4 I__4276 (
            .O(N__21429),
            .I(N__21402));
    InMux I__4275 (
            .O(N__21428),
            .I(N__21398));
    InMux I__4274 (
            .O(N__21427),
            .I(N__21395));
    Span12Mux_s7_h I__4273 (
            .O(N__21424),
            .I(N__21386));
    Span12Mux_s10_v I__4272 (
            .O(N__21419),
            .I(N__21386));
    Sp12to4 I__4271 (
            .O(N__21414),
            .I(N__21386));
    Span12Mux_v I__4270 (
            .O(N__21405),
            .I(N__21386));
    Span12Mux_h I__4269 (
            .O(N__21402),
            .I(N__21383));
    InMux I__4268 (
            .O(N__21401),
            .I(N__21380));
    LocalMux I__4267 (
            .O(N__21398),
            .I(M_this_sprites_address_qZ0Z_5));
    LocalMux I__4266 (
            .O(N__21395),
            .I(M_this_sprites_address_qZ0Z_5));
    Odrv12 I__4265 (
            .O(N__21386),
            .I(M_this_sprites_address_qZ0Z_5));
    Odrv12 I__4264 (
            .O(N__21383),
            .I(M_this_sprites_address_qZ0Z_5));
    LocalMux I__4263 (
            .O(N__21380),
            .I(M_this_sprites_address_qZ0Z_5));
    InMux I__4262 (
            .O(N__21369),
            .I(N__21366));
    LocalMux I__4261 (
            .O(N__21366),
            .I(un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0));
    InMux I__4260 (
            .O(N__21363),
            .I(un1_M_this_sprites_address_q_cry_4));
    CascadeMux I__4259 (
            .O(N__21360),
            .I(N__21356));
    CascadeMux I__4258 (
            .O(N__21359),
            .I(N__21353));
    InMux I__4257 (
            .O(N__21356),
            .I(N__21348));
    InMux I__4256 (
            .O(N__21353),
            .I(N__21345));
    CascadeMux I__4255 (
            .O(N__21352),
            .I(N__21342));
    CascadeMux I__4254 (
            .O(N__21351),
            .I(N__21339));
    LocalMux I__4253 (
            .O(N__21348),
            .I(N__21334));
    LocalMux I__4252 (
            .O(N__21345),
            .I(N__21331));
    InMux I__4251 (
            .O(N__21342),
            .I(N__21328));
    InMux I__4250 (
            .O(N__21339),
            .I(N__21325));
    CascadeMux I__4249 (
            .O(N__21338),
            .I(N__21322));
    CascadeMux I__4248 (
            .O(N__21337),
            .I(N__21319));
    Span4Mux_v I__4247 (
            .O(N__21334),
            .I(N__21310));
    Span4Mux_h I__4246 (
            .O(N__21331),
            .I(N__21310));
    LocalMux I__4245 (
            .O(N__21328),
            .I(N__21310));
    LocalMux I__4244 (
            .O(N__21325),
            .I(N__21307));
    InMux I__4243 (
            .O(N__21322),
            .I(N__21304));
    InMux I__4242 (
            .O(N__21319),
            .I(N__21301));
    CascadeMux I__4241 (
            .O(N__21318),
            .I(N__21298));
    CascadeMux I__4240 (
            .O(N__21317),
            .I(N__21293));
    Span4Mux_v I__4239 (
            .O(N__21310),
            .I(N__21284));
    Span4Mux_h I__4238 (
            .O(N__21307),
            .I(N__21284));
    LocalMux I__4237 (
            .O(N__21304),
            .I(N__21284));
    LocalMux I__4236 (
            .O(N__21301),
            .I(N__21281));
    InMux I__4235 (
            .O(N__21298),
            .I(N__21278));
    CascadeMux I__4234 (
            .O(N__21297),
            .I(N__21275));
    CascadeMux I__4233 (
            .O(N__21296),
            .I(N__21272));
    InMux I__4232 (
            .O(N__21293),
            .I(N__21267));
    CascadeMux I__4231 (
            .O(N__21292),
            .I(N__21264));
    CascadeMux I__4230 (
            .O(N__21291),
            .I(N__21261));
    Span4Mux_v I__4229 (
            .O(N__21284),
            .I(N__21253));
    Span4Mux_h I__4228 (
            .O(N__21281),
            .I(N__21253));
    LocalMux I__4227 (
            .O(N__21278),
            .I(N__21253));
    InMux I__4226 (
            .O(N__21275),
            .I(N__21250));
    InMux I__4225 (
            .O(N__21272),
            .I(N__21247));
    CascadeMux I__4224 (
            .O(N__21271),
            .I(N__21244));
    CascadeMux I__4223 (
            .O(N__21270),
            .I(N__21241));
    LocalMux I__4222 (
            .O(N__21267),
            .I(N__21238));
    InMux I__4221 (
            .O(N__21264),
            .I(N__21235));
    InMux I__4220 (
            .O(N__21261),
            .I(N__21232));
    CascadeMux I__4219 (
            .O(N__21260),
            .I(N__21229));
    Span4Mux_v I__4218 (
            .O(N__21253),
            .I(N__21226));
    LocalMux I__4217 (
            .O(N__21250),
            .I(N__21221));
    LocalMux I__4216 (
            .O(N__21247),
            .I(N__21221));
    InMux I__4215 (
            .O(N__21244),
            .I(N__21218));
    InMux I__4214 (
            .O(N__21241),
            .I(N__21215));
    Span4Mux_v I__4213 (
            .O(N__21238),
            .I(N__21208));
    LocalMux I__4212 (
            .O(N__21235),
            .I(N__21208));
    LocalMux I__4211 (
            .O(N__21232),
            .I(N__21205));
    InMux I__4210 (
            .O(N__21229),
            .I(N__21202));
    Span4Mux_v I__4209 (
            .O(N__21226),
            .I(N__21193));
    Span4Mux_v I__4208 (
            .O(N__21221),
            .I(N__21193));
    LocalMux I__4207 (
            .O(N__21218),
            .I(N__21193));
    LocalMux I__4206 (
            .O(N__21215),
            .I(N__21193));
    CascadeMux I__4205 (
            .O(N__21214),
            .I(N__21190));
    InMux I__4204 (
            .O(N__21213),
            .I(N__21187));
    Span4Mux_v I__4203 (
            .O(N__21208),
            .I(N__21181));
    Span4Mux_v I__4202 (
            .O(N__21205),
            .I(N__21181));
    LocalMux I__4201 (
            .O(N__21202),
            .I(N__21178));
    Span4Mux_v I__4200 (
            .O(N__21193),
            .I(N__21175));
    InMux I__4199 (
            .O(N__21190),
            .I(N__21172));
    LocalMux I__4198 (
            .O(N__21187),
            .I(N__21169));
    CascadeMux I__4197 (
            .O(N__21186),
            .I(N__21165));
    Sp12to4 I__4196 (
            .O(N__21181),
            .I(N__21162));
    Span12Mux_h I__4195 (
            .O(N__21178),
            .I(N__21155));
    Sp12to4 I__4194 (
            .O(N__21175),
            .I(N__21155));
    LocalMux I__4193 (
            .O(N__21172),
            .I(N__21155));
    Span4Mux_h I__4192 (
            .O(N__21169),
            .I(N__21152));
    InMux I__4191 (
            .O(N__21168),
            .I(N__21149));
    InMux I__4190 (
            .O(N__21165),
            .I(N__21146));
    Odrv12 I__4189 (
            .O(N__21162),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv12 I__4188 (
            .O(N__21155),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv4 I__4187 (
            .O(N__21152),
            .I(M_this_sprites_address_qZ0Z_6));
    LocalMux I__4186 (
            .O(N__21149),
            .I(M_this_sprites_address_qZ0Z_6));
    LocalMux I__4185 (
            .O(N__21146),
            .I(M_this_sprites_address_qZ0Z_6));
    InMux I__4184 (
            .O(N__21135),
            .I(N__21132));
    LocalMux I__4183 (
            .O(N__21132),
            .I(un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0));
    InMux I__4182 (
            .O(N__21129),
            .I(un1_M_this_sprites_address_q_cry_5));
    InMux I__4181 (
            .O(N__21126),
            .I(N__21123));
    LocalMux I__4180 (
            .O(N__21123),
            .I(N__21120));
    Span4Mux_h I__4179 (
            .O(N__21120),
            .I(N__21117));
    Span4Mux_v I__4178 (
            .O(N__21117),
            .I(N__21114));
    Span4Mux_h I__4177 (
            .O(N__21114),
            .I(N__21111));
    Odrv4 I__4176 (
            .O(N__21111),
            .I(\this_sprites_ram.mem_out_bus6_3 ));
    InMux I__4175 (
            .O(N__21108),
            .I(N__21105));
    LocalMux I__4174 (
            .O(N__21105),
            .I(N__21102));
    Span4Mux_h I__4173 (
            .O(N__21102),
            .I(N__21099));
    Span4Mux_v I__4172 (
            .O(N__21099),
            .I(N__21096));
    Odrv4 I__4171 (
            .O(N__21096),
            .I(\this_sprites_ram.mem_out_bus2_3 ));
    InMux I__4170 (
            .O(N__21093),
            .I(N__21090));
    LocalMux I__4169 (
            .O(N__21090),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ));
    InMux I__4168 (
            .O(N__21087),
            .I(N__21084));
    LocalMux I__4167 (
            .O(N__21084),
            .I(N__21081));
    Span4Mux_h I__4166 (
            .O(N__21081),
            .I(N__21078));
    Span4Mux_v I__4165 (
            .O(N__21078),
            .I(N__21075));
    Span4Mux_v I__4164 (
            .O(N__21075),
            .I(N__21072));
    Span4Mux_h I__4163 (
            .O(N__21072),
            .I(N__21069));
    Odrv4 I__4162 (
            .O(N__21069),
            .I(\this_sprites_ram.mem_out_bus7_3 ));
    InMux I__4161 (
            .O(N__21066),
            .I(N__21063));
    LocalMux I__4160 (
            .O(N__21063),
            .I(N__21060));
    Span4Mux_h I__4159 (
            .O(N__21060),
            .I(N__21057));
    Span4Mux_h I__4158 (
            .O(N__21057),
            .I(N__21054));
    Span4Mux_h I__4157 (
            .O(N__21054),
            .I(N__21051));
    Odrv4 I__4156 (
            .O(N__21051),
            .I(\this_sprites_ram.mem_out_bus3_3 ));
    InMux I__4155 (
            .O(N__21048),
            .I(N__21045));
    LocalMux I__4154 (
            .O(N__21045),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ));
    InMux I__4153 (
            .O(N__21042),
            .I(N__21039));
    LocalMux I__4152 (
            .O(N__21039),
            .I(N__21036));
    Span4Mux_h I__4151 (
            .O(N__21036),
            .I(N__21033));
    Odrv4 I__4150 (
            .O(N__21033),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__4149 (
            .O(N__21030),
            .I(N__21024));
    InMux I__4148 (
            .O(N__21029),
            .I(N__21024));
    LocalMux I__4147 (
            .O(N__21024),
            .I(N__21018));
    InMux I__4146 (
            .O(N__21023),
            .I(N__21015));
    InMux I__4145 (
            .O(N__21022),
            .I(N__21010));
    InMux I__4144 (
            .O(N__21021),
            .I(N__21010));
    Span4Mux_v I__4143 (
            .O(N__21018),
            .I(N__21007));
    LocalMux I__4142 (
            .O(N__21015),
            .I(N__21004));
    LocalMux I__4141 (
            .O(N__21010),
            .I(N__21001));
    Span4Mux_v I__4140 (
            .O(N__21007),
            .I(N__20998));
    Span4Mux_v I__4139 (
            .O(N__21004),
            .I(N__20993));
    Span4Mux_h I__4138 (
            .O(N__21001),
            .I(N__20993));
    Span4Mux_v I__4137 (
            .O(N__20998),
            .I(N__20985));
    Span4Mux_v I__4136 (
            .O(N__20993),
            .I(N__20982));
    InMux I__4135 (
            .O(N__20992),
            .I(N__20973));
    InMux I__4134 (
            .O(N__20991),
            .I(N__20973));
    InMux I__4133 (
            .O(N__20990),
            .I(N__20973));
    InMux I__4132 (
            .O(N__20989),
            .I(N__20973));
    InMux I__4131 (
            .O(N__20988),
            .I(N__20970));
    Span4Mux_v I__4130 (
            .O(N__20985),
            .I(N__20967));
    Span4Mux_v I__4129 (
            .O(N__20982),
            .I(N__20964));
    LocalMux I__4128 (
            .O(N__20973),
            .I(N__20959));
    LocalMux I__4127 (
            .O(N__20970),
            .I(N__20959));
    IoSpan4Mux I__4126 (
            .O(N__20967),
            .I(N__20956));
    Span4Mux_v I__4125 (
            .O(N__20964),
            .I(N__20953));
    Span12Mux_v I__4124 (
            .O(N__20959),
            .I(N__20950));
    Odrv4 I__4123 (
            .O(N__20956),
            .I(rst_n_c));
    Odrv4 I__4122 (
            .O(N__20953),
            .I(rst_n_c));
    Odrv12 I__4121 (
            .O(N__20950),
            .I(rst_n_c));
    InMux I__4120 (
            .O(N__20943),
            .I(N__20940));
    LocalMux I__4119 (
            .O(N__20940),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    CascadeMux I__4118 (
            .O(N__20937),
            .I(N__20931));
    InMux I__4117 (
            .O(N__20936),
            .I(N__20928));
    InMux I__4116 (
            .O(N__20935),
            .I(N__20925));
    CascadeMux I__4115 (
            .O(N__20934),
            .I(N__20921));
    InMux I__4114 (
            .O(N__20931),
            .I(N__20917));
    LocalMux I__4113 (
            .O(N__20928),
            .I(N__20914));
    LocalMux I__4112 (
            .O(N__20925),
            .I(N__20911));
    InMux I__4111 (
            .O(N__20924),
            .I(N__20904));
    InMux I__4110 (
            .O(N__20921),
            .I(N__20904));
    InMux I__4109 (
            .O(N__20920),
            .I(N__20904));
    LocalMux I__4108 (
            .O(N__20917),
            .I(this_start_data_delay_M_last_q));
    Odrv4 I__4107 (
            .O(N__20914),
            .I(this_start_data_delay_M_last_q));
    Odrv4 I__4106 (
            .O(N__20911),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__4105 (
            .O(N__20904),
            .I(this_start_data_delay_M_last_q));
    CascadeMux I__4104 (
            .O(N__20895),
            .I(N__20890));
    CascadeMux I__4103 (
            .O(N__20894),
            .I(N__20887));
    CascadeMux I__4102 (
            .O(N__20893),
            .I(N__20882));
    InMux I__4101 (
            .O(N__20890),
            .I(N__20878));
    InMux I__4100 (
            .O(N__20887),
            .I(N__20875));
    InMux I__4099 (
            .O(N__20886),
            .I(N__20866));
    InMux I__4098 (
            .O(N__20885),
            .I(N__20866));
    InMux I__4097 (
            .O(N__20882),
            .I(N__20866));
    InMux I__4096 (
            .O(N__20881),
            .I(N__20866));
    LocalMux I__4095 (
            .O(N__20878),
            .I(N__20862));
    LocalMux I__4094 (
            .O(N__20875),
            .I(N__20859));
    LocalMux I__4093 (
            .O(N__20866),
            .I(N__20856));
    InMux I__4092 (
            .O(N__20865),
            .I(N__20853));
    Span4Mux_v I__4091 (
            .O(N__20862),
            .I(N__20850));
    Span4Mux_v I__4090 (
            .O(N__20859),
            .I(N__20847));
    Span4Mux_v I__4089 (
            .O(N__20856),
            .I(N__20842));
    LocalMux I__4088 (
            .O(N__20853),
            .I(N__20842));
    Span4Mux_h I__4087 (
            .O(N__20850),
            .I(N__20837));
    Span4Mux_h I__4086 (
            .O(N__20847),
            .I(N__20837));
    Span4Mux_h I__4085 (
            .O(N__20842),
            .I(N__20834));
    Span4Mux_v I__4084 (
            .O(N__20837),
            .I(N__20831));
    Sp12to4 I__4083 (
            .O(N__20834),
            .I(N__20828));
    Sp12to4 I__4082 (
            .O(N__20831),
            .I(N__20823));
    Span12Mux_v I__4081 (
            .O(N__20828),
            .I(N__20823));
    Span12Mux_h I__4080 (
            .O(N__20823),
            .I(N__20820));
    Odrv12 I__4079 (
            .O(N__20820),
            .I(port_enb_c));
    InMux I__4078 (
            .O(N__20817),
            .I(N__20813));
    InMux I__4077 (
            .O(N__20816),
            .I(N__20810));
    LocalMux I__4076 (
            .O(N__20813),
            .I(N__20806));
    LocalMux I__4075 (
            .O(N__20810),
            .I(N__20803));
    InMux I__4074 (
            .O(N__20809),
            .I(N__20796));
    Span4Mux_h I__4073 (
            .O(N__20806),
            .I(N__20791));
    Span4Mux_v I__4072 (
            .O(N__20803),
            .I(N__20791));
    InMux I__4071 (
            .O(N__20802),
            .I(N__20782));
    InMux I__4070 (
            .O(N__20801),
            .I(N__20782));
    InMux I__4069 (
            .O(N__20800),
            .I(N__20782));
    InMux I__4068 (
            .O(N__20799),
            .I(N__20782));
    LocalMux I__4067 (
            .O(N__20796),
            .I(M_this_delay_clk_out_0));
    Odrv4 I__4066 (
            .O(N__20791),
            .I(M_this_delay_clk_out_0));
    LocalMux I__4065 (
            .O(N__20782),
            .I(M_this_delay_clk_out_0));
    CascadeMux I__4064 (
            .O(N__20775),
            .I(N_156_0_cascade_));
    InMux I__4063 (
            .O(N__20772),
            .I(N__20769));
    LocalMux I__4062 (
            .O(N__20769),
            .I(N__20766));
    Span12Mux_h I__4061 (
            .O(N__20766),
            .I(N__20763));
    Odrv12 I__4060 (
            .O(N__20763),
            .I(N_35_0));
    CascadeMux I__4059 (
            .O(N__20760),
            .I(N__20757));
    InMux I__4058 (
            .O(N__20757),
            .I(N__20754));
    LocalMux I__4057 (
            .O(N__20754),
            .I(N__20751));
    Span4Mux_v I__4056 (
            .O(N__20751),
            .I(N__20748));
    Sp12to4 I__4055 (
            .O(N__20748),
            .I(N__20745));
    Span12Mux_h I__4054 (
            .O(N__20745),
            .I(N__20742));
    Odrv12 I__4053 (
            .O(N__20742),
            .I(M_this_map_ram_read_data_5));
    InMux I__4052 (
            .O(N__20739),
            .I(N__20736));
    LocalMux I__4051 (
            .O(N__20736),
            .I(N__20733));
    Span4Mux_v I__4050 (
            .O(N__20733),
            .I(N__20730));
    Sp12to4 I__4049 (
            .O(N__20730),
            .I(N__20727));
    Span12Mux_h I__4048 (
            .O(N__20727),
            .I(N__20724));
    Odrv12 I__4047 (
            .O(N__20724),
            .I(M_this_ppu_vram_data_3));
    InMux I__4046 (
            .O(N__20721),
            .I(N__20718));
    LocalMux I__4045 (
            .O(N__20718),
            .I(N__20715));
    Span4Mux_h I__4044 (
            .O(N__20715),
            .I(N__20712));
    Span4Mux_h I__4043 (
            .O(N__20712),
            .I(N__20709));
    Span4Mux_h I__4042 (
            .O(N__20709),
            .I(N__20705));
    InMux I__4041 (
            .O(N__20708),
            .I(N__20702));
    Odrv4 I__4040 (
            .O(N__20705),
            .I(M_this_ppu_vram_data_2));
    LocalMux I__4039 (
            .O(N__20702),
            .I(M_this_ppu_vram_data_2));
    CascadeMux I__4038 (
            .O(N__20697),
            .I(M_this_ppu_vram_data_3_cascade_));
    InMux I__4037 (
            .O(N__20694),
            .I(N__20691));
    LocalMux I__4036 (
            .O(N__20691),
            .I(N__20688));
    Span12Mux_v I__4035 (
            .O(N__20688),
            .I(N__20684));
    InMux I__4034 (
            .O(N__20687),
            .I(N__20681));
    Odrv12 I__4033 (
            .O(N__20684),
            .I(M_this_ppu_vram_data_0));
    LocalMux I__4032 (
            .O(N__20681),
            .I(M_this_ppu_vram_data_0));
    CascadeMux I__4031 (
            .O(N__20676),
            .I(\this_ppu.N_156_cascade_ ));
    InMux I__4030 (
            .O(N__20673),
            .I(N__20670));
    LocalMux I__4029 (
            .O(N__20670),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3 ));
    InMux I__4028 (
            .O(N__20667),
            .I(N__20664));
    LocalMux I__4027 (
            .O(N__20664),
            .I(N__20661));
    Span4Mux_h I__4026 (
            .O(N__20661),
            .I(N__20658));
    Span4Mux_v I__4025 (
            .O(N__20658),
            .I(N__20655));
    Span4Mux_h I__4024 (
            .O(N__20655),
            .I(N__20652));
    Odrv4 I__4023 (
            .O(N__20652),
            .I(\this_sprites_ram.mem_out_bus5_2 ));
    InMux I__4022 (
            .O(N__20649),
            .I(N__20646));
    LocalMux I__4021 (
            .O(N__20646),
            .I(N__20643));
    Span4Mux_h I__4020 (
            .O(N__20643),
            .I(N__20640));
    Span4Mux_h I__4019 (
            .O(N__20640),
            .I(N__20637));
    Span4Mux_v I__4018 (
            .O(N__20637),
            .I(N__20634));
    Odrv4 I__4017 (
            .O(N__20634),
            .I(\this_sprites_ram.mem_out_bus1_2 ));
    InMux I__4016 (
            .O(N__20631),
            .I(N__20628));
    LocalMux I__4015 (
            .O(N__20628),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ));
    CascadeMux I__4014 (
            .O(N__20625),
            .I(\this_ppu.un1_M_haddress_q_3_c2_cascade_ ));
    InMux I__4013 (
            .O(N__20622),
            .I(N__20613));
    InMux I__4012 (
            .O(N__20621),
            .I(N__20613));
    InMux I__4011 (
            .O(N__20620),
            .I(N__20613));
    LocalMux I__4010 (
            .O(N__20613),
            .I(\this_ppu.un1_M_haddress_q_3_c5 ));
    InMux I__4009 (
            .O(N__20610),
            .I(N__20604));
    InMux I__4008 (
            .O(N__20609),
            .I(N__20601));
    InMux I__4007 (
            .O(N__20608),
            .I(N__20597));
    InMux I__4006 (
            .O(N__20607),
            .I(N__20594));
    LocalMux I__4005 (
            .O(N__20604),
            .I(N__20591));
    LocalMux I__4004 (
            .O(N__20601),
            .I(N__20588));
    InMux I__4003 (
            .O(N__20600),
            .I(N__20585));
    LocalMux I__4002 (
            .O(N__20597),
            .I(N__20580));
    LocalMux I__4001 (
            .O(N__20594),
            .I(N__20580));
    Span4Mux_v I__4000 (
            .O(N__20591),
            .I(N__20574));
    Span4Mux_v I__3999 (
            .O(N__20588),
            .I(N__20574));
    LocalMux I__3998 (
            .O(N__20585),
            .I(N__20571));
    Span4Mux_h I__3997 (
            .O(N__20580),
            .I(N__20568));
    InMux I__3996 (
            .O(N__20579),
            .I(N__20565));
    Odrv4 I__3995 (
            .O(N__20574),
            .I(M_this_state_d55));
    Odrv4 I__3994 (
            .O(N__20571),
            .I(M_this_state_d55));
    Odrv4 I__3993 (
            .O(N__20568),
            .I(M_this_state_d55));
    LocalMux I__3992 (
            .O(N__20565),
            .I(M_this_state_d55));
    CascadeMux I__3991 (
            .O(N__20556),
            .I(this_vga_signals_M_this_state_q_ns_i_o3_0_7_cascade_));
    CascadeMux I__3990 (
            .O(N__20553),
            .I(N__20548));
    InMux I__3989 (
            .O(N__20552),
            .I(N__20545));
    InMux I__3988 (
            .O(N__20551),
            .I(N__20542));
    InMux I__3987 (
            .O(N__20548),
            .I(N__20539));
    LocalMux I__3986 (
            .O(N__20545),
            .I(N__20536));
    LocalMux I__3985 (
            .O(N__20542),
            .I(N__20533));
    LocalMux I__3984 (
            .O(N__20539),
            .I(N__20530));
    Odrv12 I__3983 (
            .O(N__20536),
            .I(\this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3Z0Z_0 ));
    Odrv4 I__3982 (
            .O(N__20533),
            .I(\this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3Z0Z_0 ));
    Odrv4 I__3981 (
            .O(N__20530),
            .I(\this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3Z0Z_0 ));
    InMux I__3980 (
            .O(N__20523),
            .I(N__20520));
    LocalMux I__3979 (
            .O(N__20520),
            .I(N__20516));
    InMux I__3978 (
            .O(N__20519),
            .I(N__20513));
    Span4Mux_v I__3977 (
            .O(N__20516),
            .I(N__20509));
    LocalMux I__3976 (
            .O(N__20513),
            .I(N__20506));
    InMux I__3975 (
            .O(N__20512),
            .I(N__20503));
    Odrv4 I__3974 (
            .O(N__20509),
            .I(\this_vga_signals.N_279 ));
    Odrv4 I__3973 (
            .O(N__20506),
            .I(\this_vga_signals.N_279 ));
    LocalMux I__3972 (
            .O(N__20503),
            .I(\this_vga_signals.N_279 ));
    CascadeMux I__3971 (
            .O(N__20496),
            .I(N__20493));
    InMux I__3970 (
            .O(N__20493),
            .I(N__20489));
    InMux I__3969 (
            .O(N__20492),
            .I(N__20484));
    LocalMux I__3968 (
            .O(N__20489),
            .I(N__20481));
    InMux I__3967 (
            .O(N__20488),
            .I(N__20476));
    InMux I__3966 (
            .O(N__20487),
            .I(N__20476));
    LocalMux I__3965 (
            .O(N__20484),
            .I(N__20473));
    Span4Mux_h I__3964 (
            .O(N__20481),
            .I(N__20470));
    LocalMux I__3963 (
            .O(N__20476),
            .I(M_this_state_qZ0Z_6));
    Odrv4 I__3962 (
            .O(N__20473),
            .I(M_this_state_qZ0Z_6));
    Odrv4 I__3961 (
            .O(N__20470),
            .I(M_this_state_qZ0Z_6));
    InMux I__3960 (
            .O(N__20463),
            .I(N__20460));
    LocalMux I__3959 (
            .O(N__20460),
            .I(N__20455));
    InMux I__3958 (
            .O(N__20459),
            .I(N__20452));
    InMux I__3957 (
            .O(N__20458),
            .I(N__20449));
    Span4Mux_h I__3956 (
            .O(N__20455),
            .I(N__20446));
    LocalMux I__3955 (
            .O(N__20452),
            .I(N__20441));
    LocalMux I__3954 (
            .O(N__20449),
            .I(N__20441));
    Odrv4 I__3953 (
            .O(N__20446),
            .I(N_210));
    Odrv12 I__3952 (
            .O(N__20441),
            .I(N_210));
    InMux I__3951 (
            .O(N__20436),
            .I(N__20430));
    InMux I__3950 (
            .O(N__20435),
            .I(N__20426));
    InMux I__3949 (
            .O(N__20434),
            .I(N__20421));
    InMux I__3948 (
            .O(N__20433),
            .I(N__20421));
    LocalMux I__3947 (
            .O(N__20430),
            .I(N__20417));
    InMux I__3946 (
            .O(N__20429),
            .I(N__20411));
    LocalMux I__3945 (
            .O(N__20426),
            .I(N__20404));
    LocalMux I__3944 (
            .O(N__20421),
            .I(N__20404));
    InMux I__3943 (
            .O(N__20420),
            .I(N__20401));
    Span4Mux_v I__3942 (
            .O(N__20417),
            .I(N__20398));
    InMux I__3941 (
            .O(N__20416),
            .I(N__20395));
    InMux I__3940 (
            .O(N__20415),
            .I(N__20392));
    InMux I__3939 (
            .O(N__20414),
            .I(N__20389));
    LocalMux I__3938 (
            .O(N__20411),
            .I(N__20386));
    InMux I__3937 (
            .O(N__20410),
            .I(N__20383));
    InMux I__3936 (
            .O(N__20409),
            .I(N__20380));
    Span4Mux_h I__3935 (
            .O(N__20404),
            .I(N__20377));
    LocalMux I__3934 (
            .O(N__20401),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3933 (
            .O(N__20398),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__3932 (
            .O(N__20395),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__3931 (
            .O(N__20392),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__3930 (
            .O(N__20389),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3929 (
            .O(N__20386),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__3928 (
            .O(N__20383),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__3927 (
            .O(N__20380),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3926 (
            .O(N__20377),
            .I(M_this_state_qZ0Z_5));
    InMux I__3925 (
            .O(N__20358),
            .I(N__20355));
    LocalMux I__3924 (
            .O(N__20355),
            .I(N__20351));
    InMux I__3923 (
            .O(N__20354),
            .I(N__20348));
    Odrv4 I__3922 (
            .O(N__20351),
            .I(\this_vga_signals.N_166 ));
    LocalMux I__3921 (
            .O(N__20348),
            .I(\this_vga_signals.N_166 ));
    InMux I__3920 (
            .O(N__20343),
            .I(N__20339));
    InMux I__3919 (
            .O(N__20342),
            .I(N__20336));
    LocalMux I__3918 (
            .O(N__20339),
            .I(N__20330));
    LocalMux I__3917 (
            .O(N__20336),
            .I(N__20327));
    InMux I__3916 (
            .O(N__20335),
            .I(N__20320));
    InMux I__3915 (
            .O(N__20334),
            .I(N__20320));
    InMux I__3914 (
            .O(N__20333),
            .I(N__20320));
    Odrv4 I__3913 (
            .O(N__20330),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__3912 (
            .O(N__20327),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__3911 (
            .O(N__20320),
            .I(M_this_state_qZ0Z_3));
    InMux I__3910 (
            .O(N__20313),
            .I(N__20310));
    LocalMux I__3909 (
            .O(N__20310),
            .I(N__20307));
    Span4Mux_h I__3908 (
            .O(N__20307),
            .I(N__20304));
    Span4Mux_v I__3907 (
            .O(N__20304),
            .I(N__20301));
    Span4Mux_h I__3906 (
            .O(N__20301),
            .I(N__20298));
    Span4Mux_h I__3905 (
            .O(N__20298),
            .I(N__20295));
    Odrv4 I__3904 (
            .O(N__20295),
            .I(\this_sprites_ram.mem_out_bus5_1 ));
    InMux I__3903 (
            .O(N__20292),
            .I(N__20289));
    LocalMux I__3902 (
            .O(N__20289),
            .I(N__20286));
    Span4Mux_h I__3901 (
            .O(N__20286),
            .I(N__20283));
    Span4Mux_v I__3900 (
            .O(N__20283),
            .I(N__20280));
    Span4Mux_v I__3899 (
            .O(N__20280),
            .I(N__20277));
    Odrv4 I__3898 (
            .O(N__20277),
            .I(\this_sprites_ram.mem_out_bus1_1 ));
    CascadeMux I__3897 (
            .O(N__20274),
            .I(N_210_cascade_));
    InMux I__3896 (
            .O(N__20271),
            .I(N__20267));
    InMux I__3895 (
            .O(N__20270),
            .I(N__20264));
    LocalMux I__3894 (
            .O(N__20267),
            .I(\this_vga_signals.N_159_0 ));
    LocalMux I__3893 (
            .O(N__20264),
            .I(\this_vga_signals.N_159_0 ));
    CascadeMux I__3892 (
            .O(N__20259),
            .I(\this_vga_signals.N_167_0_cascade_ ));
    InMux I__3891 (
            .O(N__20256),
            .I(N__20253));
    LocalMux I__3890 (
            .O(N__20253),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5 ));
    CascadeMux I__3889 (
            .O(N__20250),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_5_cascade_ ));
    InMux I__3888 (
            .O(N__20247),
            .I(N__20244));
    LocalMux I__3887 (
            .O(N__20244),
            .I(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6 ));
    CascadeMux I__3886 (
            .O(N__20241),
            .I(N__20238));
    InMux I__3885 (
            .O(N__20238),
            .I(N__20235));
    LocalMux I__3884 (
            .O(N__20235),
            .I(N__20232));
    Span4Mux_v I__3883 (
            .O(N__20232),
            .I(N__20229));
    Span4Mux_v I__3882 (
            .O(N__20229),
            .I(N__20226));
    Odrv4 I__3881 (
            .O(N__20226),
            .I(\this_vga_signals.M_this_sprites_address_q_mZ0Z_6 ));
    CascadeMux I__3880 (
            .O(N__20223),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ));
    CascadeMux I__3879 (
            .O(N__20220),
            .I(N__20217));
    InMux I__3878 (
            .O(N__20217),
            .I(N__20214));
    LocalMux I__3877 (
            .O(N__20214),
            .I(N__20211));
    Span4Mux_v I__3876 (
            .O(N__20211),
            .I(N__20208));
    Span4Mux_v I__3875 (
            .O(N__20208),
            .I(N__20205));
    Span4Mux_v I__3874 (
            .O(N__20205),
            .I(N__20202));
    Span4Mux_h I__3873 (
            .O(N__20202),
            .I(N__20199));
    Span4Mux_h I__3872 (
            .O(N__20199),
            .I(N__20196));
    Odrv4 I__3871 (
            .O(N__20196),
            .I(M_this_map_ram_read_data_7));
    InMux I__3870 (
            .O(N__20193),
            .I(N__20190));
    LocalMux I__3869 (
            .O(N__20190),
            .I(N__20187));
    Span4Mux_v I__3868 (
            .O(N__20187),
            .I(N__20184));
    Sp12to4 I__3867 (
            .O(N__20184),
            .I(N__20181));
    Span12Mux_h I__3866 (
            .O(N__20181),
            .I(N__20178));
    Span12Mux_v I__3865 (
            .O(N__20178),
            .I(N__20175));
    Odrv12 I__3864 (
            .O(N__20175),
            .I(\this_sprites_ram.mem_out_bus7_2 ));
    InMux I__3863 (
            .O(N__20172),
            .I(N__20169));
    LocalMux I__3862 (
            .O(N__20169),
            .I(N__20166));
    Span4Mux_v I__3861 (
            .O(N__20166),
            .I(N__20163));
    Span4Mux_h I__3860 (
            .O(N__20163),
            .I(N__20160));
    Span4Mux_h I__3859 (
            .O(N__20160),
            .I(N__20157));
    Odrv4 I__3858 (
            .O(N__20157),
            .I(\this_sprites_ram.mem_out_bus3_2 ));
    InMux I__3857 (
            .O(N__20154),
            .I(N__20151));
    LocalMux I__3856 (
            .O(N__20151),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ));
    InMux I__3855 (
            .O(N__20148),
            .I(N__20141));
    InMux I__3854 (
            .O(N__20147),
            .I(N__20141));
    InMux I__3853 (
            .O(N__20146),
            .I(N__20138));
    LocalMux I__3852 (
            .O(N__20141),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    LocalMux I__3851 (
            .O(N__20138),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    InMux I__3850 (
            .O(N__20133),
            .I(N__20128));
    InMux I__3849 (
            .O(N__20132),
            .I(N__20125));
    InMux I__3848 (
            .O(N__20131),
            .I(N__20122));
    LocalMux I__3847 (
            .O(N__20128),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    LocalMux I__3846 (
            .O(N__20125),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    LocalMux I__3845 (
            .O(N__20122),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    CascadeMux I__3844 (
            .O(N__20115),
            .I(N__20111));
    CascadeMux I__3843 (
            .O(N__20114),
            .I(N__20105));
    InMux I__3842 (
            .O(N__20111),
            .I(N__20099));
    InMux I__3841 (
            .O(N__20110),
            .I(N__20096));
    InMux I__3840 (
            .O(N__20109),
            .I(N__20093));
    InMux I__3839 (
            .O(N__20108),
            .I(N__20087));
    InMux I__3838 (
            .O(N__20105),
            .I(N__20082));
    InMux I__3837 (
            .O(N__20104),
            .I(N__20082));
    InMux I__3836 (
            .O(N__20103),
            .I(N__20079));
    InMux I__3835 (
            .O(N__20102),
            .I(N__20075));
    LocalMux I__3834 (
            .O(N__20099),
            .I(N__20072));
    LocalMux I__3833 (
            .O(N__20096),
            .I(N__20069));
    LocalMux I__3832 (
            .O(N__20093),
            .I(N__20066));
    CascadeMux I__3831 (
            .O(N__20092),
            .I(N__20063));
    CascadeMux I__3830 (
            .O(N__20091),
            .I(N__20060));
    CascadeMux I__3829 (
            .O(N__20090),
            .I(N__20057));
    LocalMux I__3828 (
            .O(N__20087),
            .I(N__20054));
    LocalMux I__3827 (
            .O(N__20082),
            .I(N__20051));
    LocalMux I__3826 (
            .O(N__20079),
            .I(N__20048));
    CascadeMux I__3825 (
            .O(N__20078),
            .I(N__20045));
    LocalMux I__3824 (
            .O(N__20075),
            .I(N__20036));
    Span4Mux_v I__3823 (
            .O(N__20072),
            .I(N__20036));
    Span4Mux_v I__3822 (
            .O(N__20069),
            .I(N__20036));
    Span4Mux_h I__3821 (
            .O(N__20066),
            .I(N__20036));
    InMux I__3820 (
            .O(N__20063),
            .I(N__20031));
    InMux I__3819 (
            .O(N__20060),
            .I(N__20031));
    InMux I__3818 (
            .O(N__20057),
            .I(N__20028));
    Span4Mux_v I__3817 (
            .O(N__20054),
            .I(N__20021));
    Span4Mux_v I__3816 (
            .O(N__20051),
            .I(N__20021));
    Span4Mux_v I__3815 (
            .O(N__20048),
            .I(N__20021));
    InMux I__3814 (
            .O(N__20045),
            .I(N__20018));
    Span4Mux_h I__3813 (
            .O(N__20036),
            .I(N__20015));
    LocalMux I__3812 (
            .O(N__20031),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__3811 (
            .O(N__20028),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__3810 (
            .O(N__20021),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__3809 (
            .O(N__20018),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__3808 (
            .O(N__20015),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    CascadeMux I__3807 (
            .O(N__20004),
            .I(N__20001));
    InMux I__3806 (
            .O(N__20001),
            .I(N__19997));
    CascadeMux I__3805 (
            .O(N__20000),
            .I(N__19994));
    LocalMux I__3804 (
            .O(N__19997),
            .I(N__19991));
    InMux I__3803 (
            .O(N__19994),
            .I(N__19988));
    Span4Mux_v I__3802 (
            .O(N__19991),
            .I(N__19983));
    LocalMux I__3801 (
            .O(N__19988),
            .I(N__19983));
    Odrv4 I__3800 (
            .O(N__19983),
            .I(\this_vga_signals.line_clk_1 ));
    InMux I__3799 (
            .O(N__19980),
            .I(N__19977));
    LocalMux I__3798 (
            .O(N__19977),
            .I(N__19971));
    InMux I__3797 (
            .O(N__19976),
            .I(N__19968));
    InMux I__3796 (
            .O(N__19975),
            .I(N__19964));
    InMux I__3795 (
            .O(N__19974),
            .I(N__19961));
    Span4Mux_h I__3794 (
            .O(N__19971),
            .I(N__19958));
    LocalMux I__3793 (
            .O(N__19968),
            .I(N__19955));
    InMux I__3792 (
            .O(N__19967),
            .I(N__19952));
    LocalMux I__3791 (
            .O(N__19964),
            .I(N__19949));
    LocalMux I__3790 (
            .O(N__19961),
            .I(N__19945));
    Span4Mux_v I__3789 (
            .O(N__19958),
            .I(N__19939));
    Span4Mux_h I__3788 (
            .O(N__19955),
            .I(N__19939));
    LocalMux I__3787 (
            .O(N__19952),
            .I(N__19935));
    Span4Mux_v I__3786 (
            .O(N__19949),
            .I(N__19932));
    InMux I__3785 (
            .O(N__19948),
            .I(N__19929));
    Span4Mux_h I__3784 (
            .O(N__19945),
            .I(N__19926));
    InMux I__3783 (
            .O(N__19944),
            .I(N__19923));
    Span4Mux_v I__3782 (
            .O(N__19939),
            .I(N__19920));
    InMux I__3781 (
            .O(N__19938),
            .I(N__19917));
    Span4Mux_h I__3780 (
            .O(N__19935),
            .I(N__19914));
    Span4Mux_v I__3779 (
            .O(N__19932),
            .I(N__19909));
    LocalMux I__3778 (
            .O(N__19929),
            .I(N__19909));
    Span4Mux_v I__3777 (
            .O(N__19926),
            .I(N__19906));
    LocalMux I__3776 (
            .O(N__19923),
            .I(N__19903));
    Sp12to4 I__3775 (
            .O(N__19920),
            .I(N__19898));
    LocalMux I__3774 (
            .O(N__19917),
            .I(N__19898));
    Span4Mux_h I__3773 (
            .O(N__19914),
            .I(N__19895));
    Span4Mux_h I__3772 (
            .O(N__19909),
            .I(N__19892));
    Span4Mux_h I__3771 (
            .O(N__19906),
            .I(N__19889));
    Span12Mux_h I__3770 (
            .O(N__19903),
            .I(N__19884));
    Span12Mux_h I__3769 (
            .O(N__19898),
            .I(N__19884));
    Span4Mux_h I__3768 (
            .O(N__19895),
            .I(N__19879));
    Span4Mux_h I__3767 (
            .O(N__19892),
            .I(N__19879));
    Odrv4 I__3766 (
            .O(N__19889),
            .I(M_this_sprites_ram_write_data_3));
    Odrv12 I__3765 (
            .O(N__19884),
            .I(M_this_sprites_ram_write_data_3));
    Odrv4 I__3764 (
            .O(N__19879),
            .I(M_this_sprites_ram_write_data_3));
    InMux I__3763 (
            .O(N__19872),
            .I(N__19866));
    InMux I__3762 (
            .O(N__19871),
            .I(N__19866));
    LocalMux I__3761 (
            .O(N__19866),
            .I(N__19863));
    Span4Mux_h I__3760 (
            .O(N__19863),
            .I(N__19859));
    InMux I__3759 (
            .O(N__19862),
            .I(N__19856));
    Odrv4 I__3758 (
            .O(N__19859),
            .I(\this_vga_signals.N_169_0 ));
    LocalMux I__3757 (
            .O(N__19856),
            .I(\this_vga_signals.N_169_0 ));
    InMux I__3756 (
            .O(N__19851),
            .I(N__19848));
    LocalMux I__3755 (
            .O(N__19848),
            .I(N__19845));
    Span4Mux_v I__3754 (
            .O(N__19845),
            .I(N__19842));
    Sp12to4 I__3753 (
            .O(N__19842),
            .I(N__19839));
    Span12Mux_h I__3752 (
            .O(N__19839),
            .I(N__19836));
    Odrv12 I__3751 (
            .O(N__19836),
            .I(\this_sprites_ram.mem_out_bus5_0 ));
    InMux I__3750 (
            .O(N__19833),
            .I(N__19830));
    LocalMux I__3749 (
            .O(N__19830),
            .I(N__19827));
    Span4Mux_h I__3748 (
            .O(N__19827),
            .I(N__19824));
    Span4Mux_h I__3747 (
            .O(N__19824),
            .I(N__19821));
    Span4Mux_v I__3746 (
            .O(N__19821),
            .I(N__19818));
    Odrv4 I__3745 (
            .O(N__19818),
            .I(\this_sprites_ram.mem_out_bus1_0 ));
    InMux I__3744 (
            .O(N__19815),
            .I(N__19812));
    LocalMux I__3743 (
            .O(N__19812),
            .I(N__19809));
    Span4Mux_v I__3742 (
            .O(N__19809),
            .I(N__19806));
    Span4Mux_v I__3741 (
            .O(N__19806),
            .I(N__19803));
    Sp12to4 I__3740 (
            .O(N__19803),
            .I(N__19800));
    Odrv12 I__3739 (
            .O(N__19800),
            .I(\this_sprites_ram.mem_out_bus4_0 ));
    InMux I__3738 (
            .O(N__19797),
            .I(N__19794));
    LocalMux I__3737 (
            .O(N__19794),
            .I(N__19791));
    Span4Mux_h I__3736 (
            .O(N__19791),
            .I(N__19788));
    Span4Mux_h I__3735 (
            .O(N__19788),
            .I(N__19785));
    Span4Mux_v I__3734 (
            .O(N__19785),
            .I(N__19782));
    Span4Mux_v I__3733 (
            .O(N__19782),
            .I(N__19779));
    Odrv4 I__3732 (
            .O(N__19779),
            .I(\this_sprites_ram.mem_out_bus0_0 ));
    CascadeMux I__3731 (
            .O(N__19776),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_ ));
    InMux I__3730 (
            .O(N__19773),
            .I(N__19770));
    LocalMux I__3729 (
            .O(N__19770),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ));
    InMux I__3728 (
            .O(N__19767),
            .I(N__19764));
    LocalMux I__3727 (
            .O(N__19764),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ));
    CascadeMux I__3726 (
            .O(N__19761),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_ ));
    InMux I__3725 (
            .O(N__19758),
            .I(N__19755));
    LocalMux I__3724 (
            .O(N__19755),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ));
    InMux I__3723 (
            .O(N__19752),
            .I(N__19749));
    LocalMux I__3722 (
            .O(N__19749),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    InMux I__3721 (
            .O(N__19746),
            .I(N__19743));
    LocalMux I__3720 (
            .O(N__19743),
            .I(\this_reset_cond.M_stage_qZ0Z_3 ));
    InMux I__3719 (
            .O(N__19740),
            .I(N__19737));
    LocalMux I__3718 (
            .O(N__19737),
            .I(\this_reset_cond.M_stage_qZ0Z_4 ));
    InMux I__3717 (
            .O(N__19734),
            .I(N__19731));
    LocalMux I__3716 (
            .O(N__19731),
            .I(N__19728));
    Span4Mux_v I__3715 (
            .O(N__19728),
            .I(N__19725));
    Span4Mux_v I__3714 (
            .O(N__19725),
            .I(N__19722));
    Sp12to4 I__3713 (
            .O(N__19722),
            .I(N__19719));
    Odrv12 I__3712 (
            .O(N__19719),
            .I(\this_sprites_ram.mem_out_bus4_2 ));
    InMux I__3711 (
            .O(N__19716),
            .I(N__19713));
    LocalMux I__3710 (
            .O(N__19713),
            .I(N__19710));
    Span4Mux_h I__3709 (
            .O(N__19710),
            .I(N__19707));
    Span4Mux_h I__3708 (
            .O(N__19707),
            .I(N__19704));
    Span4Mux_v I__3707 (
            .O(N__19704),
            .I(N__19701));
    Span4Mux_v I__3706 (
            .O(N__19701),
            .I(N__19698));
    Odrv4 I__3705 (
            .O(N__19698),
            .I(\this_sprites_ram.mem_out_bus0_2 ));
    CascadeMux I__3704 (
            .O(N__19695),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ));
    CascadeMux I__3703 (
            .O(N__19692),
            .I(N__19686));
    InMux I__3702 (
            .O(N__19691),
            .I(N__19683));
    InMux I__3701 (
            .O(N__19690),
            .I(N__19678));
    InMux I__3700 (
            .O(N__19689),
            .I(N__19678));
    InMux I__3699 (
            .O(N__19686),
            .I(N__19675));
    LocalMux I__3698 (
            .O(N__19683),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__3697 (
            .O(N__19678),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__3696 (
            .O(N__19675),
            .I(M_this_state_qZ0Z_11));
    InMux I__3695 (
            .O(N__19668),
            .I(N__19662));
    InMux I__3694 (
            .O(N__19667),
            .I(N__19662));
    LocalMux I__3693 (
            .O(N__19662),
            .I(N_456_0_1));
    InMux I__3692 (
            .O(N__19659),
            .I(N__19656));
    LocalMux I__3691 (
            .O(N__19656),
            .I(N_500));
    InMux I__3690 (
            .O(N__19653),
            .I(N__19648));
    InMux I__3689 (
            .O(N__19652),
            .I(N__19644));
    InMux I__3688 (
            .O(N__19651),
            .I(N__19637));
    LocalMux I__3687 (
            .O(N__19648),
            .I(N__19634));
    InMux I__3686 (
            .O(N__19647),
            .I(N__19631));
    LocalMux I__3685 (
            .O(N__19644),
            .I(N__19628));
    InMux I__3684 (
            .O(N__19643),
            .I(N__19625));
    InMux I__3683 (
            .O(N__19642),
            .I(N__19622));
    InMux I__3682 (
            .O(N__19641),
            .I(N__19619));
    InMux I__3681 (
            .O(N__19640),
            .I(N__19616));
    LocalMux I__3680 (
            .O(N__19637),
            .I(N__19613));
    Span12Mux_h I__3679 (
            .O(N__19634),
            .I(N__19610));
    LocalMux I__3678 (
            .O(N__19631),
            .I(N__19607));
    Span12Mux_s11_v I__3677 (
            .O(N__19628),
            .I(N__19602));
    LocalMux I__3676 (
            .O(N__19625),
            .I(N__19602));
    LocalMux I__3675 (
            .O(N__19622),
            .I(N__19599));
    LocalMux I__3674 (
            .O(N__19619),
            .I(N__19596));
    LocalMux I__3673 (
            .O(N__19616),
            .I(N__19593));
    Span12Mux_h I__3672 (
            .O(N__19613),
            .I(N__19590));
    Span12Mux_v I__3671 (
            .O(N__19610),
            .I(N__19585));
    Span12Mux_h I__3670 (
            .O(N__19607),
            .I(N__19585));
    Span12Mux_v I__3669 (
            .O(N__19602),
            .I(N__19576));
    Span12Mux_s8_v I__3668 (
            .O(N__19599),
            .I(N__19576));
    Span12Mux_h I__3667 (
            .O(N__19596),
            .I(N__19576));
    Span12Mux_s7_h I__3666 (
            .O(N__19593),
            .I(N__19576));
    Odrv12 I__3665 (
            .O(N__19590),
            .I(M_this_sprites_ram_write_data_0));
    Odrv12 I__3664 (
            .O(N__19585),
            .I(M_this_sprites_ram_write_data_0));
    Odrv12 I__3663 (
            .O(N__19576),
            .I(M_this_sprites_ram_write_data_0));
    CascadeMux I__3662 (
            .O(N__19569),
            .I(N__19566));
    InMux I__3661 (
            .O(N__19566),
            .I(N__19563));
    LocalMux I__3660 (
            .O(N__19563),
            .I(N__19559));
    InMux I__3659 (
            .O(N__19562),
            .I(N__19556));
    Span4Mux_v I__3658 (
            .O(N__19559),
            .I(N__19553));
    LocalMux I__3657 (
            .O(N__19556),
            .I(N__19550));
    Odrv4 I__3656 (
            .O(N__19553),
            .I(M_this_state_d_2_sqmuxa));
    Odrv4 I__3655 (
            .O(N__19550),
            .I(M_this_state_d_2_sqmuxa));
    InMux I__3654 (
            .O(N__19545),
            .I(N__19540));
    InMux I__3653 (
            .O(N__19544),
            .I(N__19537));
    InMux I__3652 (
            .O(N__19543),
            .I(N__19534));
    LocalMux I__3651 (
            .O(N__19540),
            .I(M_this_substate_qZ0));
    LocalMux I__3650 (
            .O(N__19537),
            .I(M_this_substate_qZ0));
    LocalMux I__3649 (
            .O(N__19534),
            .I(M_this_substate_qZ0));
    CascadeMux I__3648 (
            .O(N__19527),
            .I(N__19523));
    InMux I__3647 (
            .O(N__19526),
            .I(N__19518));
    InMux I__3646 (
            .O(N__19523),
            .I(N__19518));
    LocalMux I__3645 (
            .O(N__19518),
            .I(N__19515));
    Odrv4 I__3644 (
            .O(N__19515),
            .I(this_vga_signals_M_this_state_q_ns_0_a3_0_0_1));
    InMux I__3643 (
            .O(N__19512),
            .I(N__19509));
    LocalMux I__3642 (
            .O(N__19509),
            .I(N__19506));
    Span4Mux_v I__3641 (
            .O(N__19506),
            .I(N__19503));
    Sp12to4 I__3640 (
            .O(N__19503),
            .I(N__19500));
    Span12Mux_h I__3639 (
            .O(N__19500),
            .I(N__19497));
    Span12Mux_v I__3638 (
            .O(N__19497),
            .I(N__19494));
    Odrv12 I__3637 (
            .O(N__19494),
            .I(\this_sprites_ram.mem_out_bus7_0 ));
    InMux I__3636 (
            .O(N__19491),
            .I(N__19488));
    LocalMux I__3635 (
            .O(N__19488),
            .I(N__19485));
    Span4Mux_h I__3634 (
            .O(N__19485),
            .I(N__19482));
    Span4Mux_h I__3633 (
            .O(N__19482),
            .I(N__19479));
    Odrv4 I__3632 (
            .O(N__19479),
            .I(\this_sprites_ram.mem_out_bus3_0 ));
    InMux I__3631 (
            .O(N__19476),
            .I(N__19473));
    LocalMux I__3630 (
            .O(N__19473),
            .I(N__19470));
    Span4Mux_h I__3629 (
            .O(N__19470),
            .I(N__19467));
    Span4Mux_v I__3628 (
            .O(N__19467),
            .I(N__19464));
    Span4Mux_v I__3627 (
            .O(N__19464),
            .I(N__19461));
    Span4Mux_h I__3626 (
            .O(N__19461),
            .I(N__19458));
    Odrv4 I__3625 (
            .O(N__19458),
            .I(\this_sprites_ram.mem_out_bus6_0 ));
    InMux I__3624 (
            .O(N__19455),
            .I(N__19452));
    LocalMux I__3623 (
            .O(N__19452),
            .I(N__19449));
    Span4Mux_h I__3622 (
            .O(N__19449),
            .I(N__19446));
    Span4Mux_h I__3621 (
            .O(N__19446),
            .I(N__19443));
    Odrv4 I__3620 (
            .O(N__19443),
            .I(\this_sprites_ram.mem_out_bus2_0 ));
    InMux I__3619 (
            .O(N__19440),
            .I(N__19437));
    LocalMux I__3618 (
            .O(N__19437),
            .I(N__19433));
    CascadeMux I__3617 (
            .O(N__19436),
            .I(N__19430));
    Span4Mux_v I__3616 (
            .O(N__19433),
            .I(N__19427));
    InMux I__3615 (
            .O(N__19430),
            .I(N__19424));
    Span4Mux_h I__3614 (
            .O(N__19427),
            .I(N__19421));
    LocalMux I__3613 (
            .O(N__19424),
            .I(N__19418));
    Odrv4 I__3612 (
            .O(N__19421),
            .I(this_vga_signals_N_419_i_i_0_a3_1_0));
    Odrv4 I__3611 (
            .O(N__19418),
            .I(this_vga_signals_N_419_i_i_0_a3_1_0));
    CascadeMux I__3610 (
            .O(N__19413),
            .I(N_496_0_cascade_));
    InMux I__3609 (
            .O(N__19410),
            .I(N__19406));
    InMux I__3608 (
            .O(N__19409),
            .I(N__19403));
    LocalMux I__3607 (
            .O(N__19406),
            .I(N__19400));
    LocalMux I__3606 (
            .O(N__19403),
            .I(N__19397));
    Span4Mux_h I__3605 (
            .O(N__19400),
            .I(N__19390));
    Span4Mux_h I__3604 (
            .O(N__19397),
            .I(N__19390));
    InMux I__3603 (
            .O(N__19396),
            .I(N__19385));
    InMux I__3602 (
            .O(N__19395),
            .I(N__19385));
    Odrv4 I__3601 (
            .O(N__19390),
            .I(N_278));
    LocalMux I__3600 (
            .O(N__19385),
            .I(N_278));
    CascadeMux I__3599 (
            .O(N__19380),
            .I(M_this_state_qsr_0_cascade_));
    InMux I__3598 (
            .O(N__19377),
            .I(N__19374));
    LocalMux I__3597 (
            .O(N__19374),
            .I(N_462_0));
    CascadeMux I__3596 (
            .O(N__19371),
            .I(M_this_state_qsr_2_cascade_));
    InMux I__3595 (
            .O(N__19368),
            .I(N__19365));
    LocalMux I__3594 (
            .O(N__19365),
            .I(N__19362));
    Span4Mux_h I__3593 (
            .O(N__19362),
            .I(N__19357));
    InMux I__3592 (
            .O(N__19361),
            .I(N__19352));
    InMux I__3591 (
            .O(N__19360),
            .I(N__19352));
    Odrv4 I__3590 (
            .O(N__19357),
            .I(N_484_0));
    LocalMux I__3589 (
            .O(N__19352),
            .I(N_484_0));
    CascadeMux I__3588 (
            .O(N__19347),
            .I(\this_vga_signals.N_159_0_cascade_ ));
    InMux I__3587 (
            .O(N__19344),
            .I(N__19340));
    InMux I__3586 (
            .O(N__19343),
            .I(N__19335));
    LocalMux I__3585 (
            .O(N__19340),
            .I(N__19332));
    InMux I__3584 (
            .O(N__19339),
            .I(N__19329));
    InMux I__3583 (
            .O(N__19338),
            .I(N__19326));
    LocalMux I__3582 (
            .O(N__19335),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__3581 (
            .O(N__19332),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__3580 (
            .O(N__19329),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__3579 (
            .O(N__19326),
            .I(M_this_state_qZ0Z_9));
    InMux I__3578 (
            .O(N__19317),
            .I(N__19314));
    LocalMux I__3577 (
            .O(N__19314),
            .I(N__19310));
    InMux I__3576 (
            .O(N__19313),
            .I(N__19307));
    Span4Mux_v I__3575 (
            .O(N__19310),
            .I(N__19302));
    LocalMux I__3574 (
            .O(N__19307),
            .I(N__19302));
    Odrv4 I__3573 (
            .O(N__19302),
            .I(N_168_0));
    CascadeMux I__3572 (
            .O(N__19299),
            .I(N_168_0_cascade_));
    InMux I__3571 (
            .O(N__19296),
            .I(N__19293));
    LocalMux I__3570 (
            .O(N__19293),
            .I(\this_vga_signals.M_this_external_address_d_0_sqmuxa_1Z0Z_2 ));
    CascadeMux I__3569 (
            .O(N__19290),
            .I(N__19285));
    InMux I__3568 (
            .O(N__19289),
            .I(N__19278));
    InMux I__3567 (
            .O(N__19288),
            .I(N__19278));
    InMux I__3566 (
            .O(N__19285),
            .I(N__19273));
    InMux I__3565 (
            .O(N__19284),
            .I(N__19273));
    InMux I__3564 (
            .O(N__19283),
            .I(N__19270));
    LocalMux I__3563 (
            .O(N__19278),
            .I(\this_ppu.un16_0 ));
    LocalMux I__3562 (
            .O(N__19273),
            .I(\this_ppu.un16_0 ));
    LocalMux I__3561 (
            .O(N__19270),
            .I(\this_ppu.un16_0 ));
    InMux I__3560 (
            .O(N__19263),
            .I(N__19260));
    LocalMux I__3559 (
            .O(N__19260),
            .I(\this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ));
    CascadeMux I__3558 (
            .O(N__19257),
            .I(\this_ppu.un16_0_cascade_ ));
    InMux I__3557 (
            .O(N__19254),
            .I(N__19240));
    InMux I__3556 (
            .O(N__19253),
            .I(N__19240));
    InMux I__3555 (
            .O(N__19252),
            .I(N__19240));
    InMux I__3554 (
            .O(N__19251),
            .I(N__19240));
    InMux I__3553 (
            .O(N__19250),
            .I(N__19237));
    InMux I__3552 (
            .O(N__19249),
            .I(N__19234));
    LocalMux I__3551 (
            .O(N__19240),
            .I(\this_ppu.N_1157_0 ));
    LocalMux I__3550 (
            .O(N__19237),
            .I(\this_ppu.N_1157_0 ));
    LocalMux I__3549 (
            .O(N__19234),
            .I(\this_ppu.N_1157_0 ));
    CascadeMux I__3548 (
            .O(N__19227),
            .I(N__19224));
    InMux I__3547 (
            .O(N__19224),
            .I(N__19221));
    LocalMux I__3546 (
            .O(N__19221),
            .I(N__19216));
    InMux I__3545 (
            .O(N__19220),
            .I(N__19213));
    InMux I__3544 (
            .O(N__19219),
            .I(N__19210));
    Span4Mux_h I__3543 (
            .O(N__19216),
            .I(N__19207));
    LocalMux I__3542 (
            .O(N__19213),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    LocalMux I__3541 (
            .O(N__19210),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    Odrv4 I__3540 (
            .O(N__19207),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    CascadeMux I__3539 (
            .O(N__19200),
            .I(N_459_0_cascade_));
    CascadeMux I__3538 (
            .O(N__19197),
            .I(N_458_0_cascade_));
    CascadeMux I__3537 (
            .O(N__19194),
            .I(\this_ppu.N_132_0_cascade_ ));
    InMux I__3536 (
            .O(N__19191),
            .I(N__19186));
    InMux I__3535 (
            .O(N__19190),
            .I(N__19181));
    InMux I__3534 (
            .O(N__19189),
            .I(N__19181));
    LocalMux I__3533 (
            .O(N__19186),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    LocalMux I__3532 (
            .O(N__19181),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    InMux I__3531 (
            .O(N__19176),
            .I(N__19173));
    LocalMux I__3530 (
            .O(N__19173),
            .I(N__19170));
    Span4Mux_h I__3529 (
            .O(N__19170),
            .I(N__19167));
    Odrv4 I__3528 (
            .O(N__19167),
            .I(\this_vga_signals.M_vcounter_d8 ));
    CascadeMux I__3527 (
            .O(N__19164),
            .I(\this_vga_signals.un1_M_hcounter_d7_1_0_cascade_ ));
    CascadeMux I__3526 (
            .O(N__19161),
            .I(N__19158));
    InMux I__3525 (
            .O(N__19158),
            .I(N__19155));
    LocalMux I__3524 (
            .O(N__19155),
            .I(\this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ));
    InMux I__3523 (
            .O(N__19152),
            .I(N__19147));
    InMux I__3522 (
            .O(N__19151),
            .I(N__19144));
    InMux I__3521 (
            .O(N__19150),
            .I(N__19141));
    LocalMux I__3520 (
            .O(N__19147),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    LocalMux I__3519 (
            .O(N__19144),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    LocalMux I__3518 (
            .O(N__19141),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    InMux I__3517 (
            .O(N__19134),
            .I(N__19124));
    InMux I__3516 (
            .O(N__19133),
            .I(N__19124));
    InMux I__3515 (
            .O(N__19132),
            .I(N__19124));
    CascadeMux I__3514 (
            .O(N__19131),
            .I(N__19120));
    LocalMux I__3513 (
            .O(N__19124),
            .I(N__19116));
    InMux I__3512 (
            .O(N__19123),
            .I(N__19109));
    InMux I__3511 (
            .O(N__19120),
            .I(N__19106));
    InMux I__3510 (
            .O(N__19119),
            .I(N__19103));
    Span4Mux_v I__3509 (
            .O(N__19116),
            .I(N__19099));
    InMux I__3508 (
            .O(N__19115),
            .I(N__19090));
    InMux I__3507 (
            .O(N__19114),
            .I(N__19090));
    InMux I__3506 (
            .O(N__19113),
            .I(N__19090));
    InMux I__3505 (
            .O(N__19112),
            .I(N__19090));
    LocalMux I__3504 (
            .O(N__19109),
            .I(N__19083));
    LocalMux I__3503 (
            .O(N__19106),
            .I(N__19083));
    LocalMux I__3502 (
            .O(N__19103),
            .I(N__19083));
    InMux I__3501 (
            .O(N__19102),
            .I(N__19080));
    Span4Mux_h I__3500 (
            .O(N__19099),
            .I(N__19075));
    LocalMux I__3499 (
            .O(N__19090),
            .I(N__19075));
    Span4Mux_h I__3498 (
            .O(N__19083),
            .I(N__19072));
    LocalMux I__3497 (
            .O(N__19080),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__3496 (
            .O(N__19075),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__3495 (
            .O(N__19072),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    InMux I__3494 (
            .O(N__19065),
            .I(N__19048));
    InMux I__3493 (
            .O(N__19064),
            .I(N__19048));
    InMux I__3492 (
            .O(N__19063),
            .I(N__19039));
    InMux I__3491 (
            .O(N__19062),
            .I(N__19039));
    InMux I__3490 (
            .O(N__19061),
            .I(N__19039));
    InMux I__3489 (
            .O(N__19060),
            .I(N__19039));
    InMux I__3488 (
            .O(N__19059),
            .I(N__19032));
    InMux I__3487 (
            .O(N__19058),
            .I(N__19032));
    InMux I__3486 (
            .O(N__19057),
            .I(N__19032));
    InMux I__3485 (
            .O(N__19056),
            .I(N__19029));
    InMux I__3484 (
            .O(N__19055),
            .I(N__19026));
    InMux I__3483 (
            .O(N__19054),
            .I(N__19020));
    InMux I__3482 (
            .O(N__19053),
            .I(N__19020));
    LocalMux I__3481 (
            .O(N__19048),
            .I(N__19013));
    LocalMux I__3480 (
            .O(N__19039),
            .I(N__19013));
    LocalMux I__3479 (
            .O(N__19032),
            .I(N__19013));
    LocalMux I__3478 (
            .O(N__19029),
            .I(N__19010));
    LocalMux I__3477 (
            .O(N__19026),
            .I(N__19004));
    InMux I__3476 (
            .O(N__19025),
            .I(N__19001));
    LocalMux I__3475 (
            .O(N__19020),
            .I(N__18994));
    Span4Mux_v I__3474 (
            .O(N__19013),
            .I(N__18991));
    Span12Mux_s1_h I__3473 (
            .O(N__19010),
            .I(N__18988));
    CEMux I__3472 (
            .O(N__19009),
            .I(N__18985));
    InMux I__3471 (
            .O(N__19008),
            .I(N__18980));
    InMux I__3470 (
            .O(N__19007),
            .I(N__18980));
    Span4Mux_v I__3469 (
            .O(N__19004),
            .I(N__18975));
    LocalMux I__3468 (
            .O(N__19001),
            .I(N__18975));
    InMux I__3467 (
            .O(N__19000),
            .I(N__18969));
    InMux I__3466 (
            .O(N__18999),
            .I(N__18969));
    InMux I__3465 (
            .O(N__18998),
            .I(N__18964));
    InMux I__3464 (
            .O(N__18997),
            .I(N__18964));
    Span4Mux_h I__3463 (
            .O(N__18994),
            .I(N__18961));
    Span4Mux_h I__3462 (
            .O(N__18991),
            .I(N__18958));
    Span12Mux_h I__3461 (
            .O(N__18988),
            .I(N__18955));
    LocalMux I__3460 (
            .O(N__18985),
            .I(N__18948));
    LocalMux I__3459 (
            .O(N__18980),
            .I(N__18948));
    Span4Mux_h I__3458 (
            .O(N__18975),
            .I(N__18948));
    InMux I__3457 (
            .O(N__18974),
            .I(N__18945));
    LocalMux I__3456 (
            .O(N__18969),
            .I(\this_vga_signals.GZ0Z_330 ));
    LocalMux I__3455 (
            .O(N__18964),
            .I(\this_vga_signals.GZ0Z_330 ));
    Odrv4 I__3454 (
            .O(N__18961),
            .I(\this_vga_signals.GZ0Z_330 ));
    Odrv4 I__3453 (
            .O(N__18958),
            .I(\this_vga_signals.GZ0Z_330 ));
    Odrv12 I__3452 (
            .O(N__18955),
            .I(\this_vga_signals.GZ0Z_330 ));
    Odrv4 I__3451 (
            .O(N__18948),
            .I(\this_vga_signals.GZ0Z_330 ));
    LocalMux I__3450 (
            .O(N__18945),
            .I(\this_vga_signals.GZ0Z_330 ));
    InMux I__3449 (
            .O(N__18930),
            .I(N__18927));
    LocalMux I__3448 (
            .O(N__18927),
            .I(\this_vga_signals.un1_M_hcounter_d7_1_0 ));
    CascadeMux I__3447 (
            .O(N__18924),
            .I(\this_vga_signals.CO0_cascade_ ));
    InMux I__3446 (
            .O(N__18921),
            .I(N__18914));
    InMux I__3445 (
            .O(N__18920),
            .I(N__18914));
    InMux I__3444 (
            .O(N__18919),
            .I(N__18911));
    LocalMux I__3443 (
            .O(N__18914),
            .I(\this_ppu.N_1157_0_1 ));
    LocalMux I__3442 (
            .O(N__18911),
            .I(\this_ppu.N_1157_0_1 ));
    InMux I__3441 (
            .O(N__18906),
            .I(N__18903));
    LocalMux I__3440 (
            .O(N__18903),
            .I(\this_vga_signals.M_this_state_d55Z0Z_9 ));
    InMux I__3439 (
            .O(N__18900),
            .I(N__18897));
    LocalMux I__3438 (
            .O(N__18897),
            .I(\this_vga_signals.M_this_state_d55Z0Z_8 ));
    CascadeMux I__3437 (
            .O(N__18894),
            .I(\this_vga_signals.M_this_state_d55Z0Z_7_cascade_ ));
    InMux I__3436 (
            .O(N__18891),
            .I(N__18888));
    LocalMux I__3435 (
            .O(N__18888),
            .I(\this_vga_signals.M_this_state_d55Z0Z_6 ));
    InMux I__3434 (
            .O(N__18885),
            .I(N__18880));
    InMux I__3433 (
            .O(N__18884),
            .I(N__18875));
    InMux I__3432 (
            .O(N__18883),
            .I(N__18875));
    LocalMux I__3431 (
            .O(N__18880),
            .I(N__18872));
    LocalMux I__3430 (
            .O(N__18875),
            .I(N__18868));
    Span4Mux_v I__3429 (
            .O(N__18872),
            .I(N__18865));
    InMux I__3428 (
            .O(N__18871),
            .I(N__18862));
    Span4Mux_v I__3427 (
            .O(N__18868),
            .I(N__18859));
    Sp12to4 I__3426 (
            .O(N__18865),
            .I(N__18853));
    LocalMux I__3425 (
            .O(N__18862),
            .I(N__18853));
    Span4Mux_h I__3424 (
            .O(N__18859),
            .I(N__18850));
    InMux I__3423 (
            .O(N__18858),
            .I(N__18847));
    Odrv12 I__3422 (
            .O(N__18853),
            .I(M_this_vram_read_data_2));
    Odrv4 I__3421 (
            .O(N__18850),
            .I(M_this_vram_read_data_2));
    LocalMux I__3420 (
            .O(N__18847),
            .I(M_this_vram_read_data_2));
    CascadeMux I__3419 (
            .O(N__18840),
            .I(N__18836));
    CascadeMux I__3418 (
            .O(N__18839),
            .I(N__18833));
    InMux I__3417 (
            .O(N__18836),
            .I(N__18824));
    InMux I__3416 (
            .O(N__18833),
            .I(N__18824));
    InMux I__3415 (
            .O(N__18832),
            .I(N__18824));
    InMux I__3414 (
            .O(N__18831),
            .I(N__18821));
    LocalMux I__3413 (
            .O(N__18824),
            .I(N__18817));
    LocalMux I__3412 (
            .O(N__18821),
            .I(N__18814));
    InMux I__3411 (
            .O(N__18820),
            .I(N__18810));
    Span4Mux_v I__3410 (
            .O(N__18817),
            .I(N__18807));
    Span4Mux_v I__3409 (
            .O(N__18814),
            .I(N__18804));
    InMux I__3408 (
            .O(N__18813),
            .I(N__18801));
    LocalMux I__3407 (
            .O(N__18810),
            .I(N__18794));
    Sp12to4 I__3406 (
            .O(N__18807),
            .I(N__18794));
    Sp12to4 I__3405 (
            .O(N__18804),
            .I(N__18794));
    LocalMux I__3404 (
            .O(N__18801),
            .I(M_this_vram_read_data_1));
    Odrv12 I__3403 (
            .O(N__18794),
            .I(M_this_vram_read_data_1));
    CascadeMux I__3402 (
            .O(N__18789),
            .I(N__18786));
    InMux I__3401 (
            .O(N__18786),
            .I(N__18781));
    CascadeMux I__3400 (
            .O(N__18785),
            .I(N__18778));
    CascadeMux I__3399 (
            .O(N__18784),
            .I(N__18774));
    LocalMux I__3398 (
            .O(N__18781),
            .I(N__18770));
    InMux I__3397 (
            .O(N__18778),
            .I(N__18767));
    InMux I__3396 (
            .O(N__18777),
            .I(N__18760));
    InMux I__3395 (
            .O(N__18774),
            .I(N__18760));
    InMux I__3394 (
            .O(N__18773),
            .I(N__18760));
    Span4Mux_v I__3393 (
            .O(N__18770),
            .I(N__18756));
    LocalMux I__3392 (
            .O(N__18767),
            .I(N__18751));
    LocalMux I__3391 (
            .O(N__18760),
            .I(N__18751));
    CascadeMux I__3390 (
            .O(N__18759),
            .I(N__18748));
    Span4Mux_h I__3389 (
            .O(N__18756),
            .I(N__18743));
    Span4Mux_v I__3388 (
            .O(N__18751),
            .I(N__18743));
    InMux I__3387 (
            .O(N__18748),
            .I(N__18740));
    Span4Mux_h I__3386 (
            .O(N__18743),
            .I(N__18737));
    LocalMux I__3385 (
            .O(N__18740),
            .I(M_this_vram_read_data_3));
    Odrv4 I__3384 (
            .O(N__18737),
            .I(M_this_vram_read_data_3));
    InMux I__3383 (
            .O(N__18732),
            .I(N__18726));
    InMux I__3382 (
            .O(N__18731),
            .I(N__18719));
    InMux I__3381 (
            .O(N__18730),
            .I(N__18719));
    InMux I__3380 (
            .O(N__18729),
            .I(N__18719));
    LocalMux I__3379 (
            .O(N__18726),
            .I(N__18716));
    LocalMux I__3378 (
            .O(N__18719),
            .I(N__18712));
    Span4Mux_v I__3377 (
            .O(N__18716),
            .I(N__18709));
    InMux I__3376 (
            .O(N__18715),
            .I(N__18706));
    Span4Mux_h I__3375 (
            .O(N__18712),
            .I(N__18703));
    Sp12to4 I__3374 (
            .O(N__18709),
            .I(N__18697));
    LocalMux I__3373 (
            .O(N__18706),
            .I(N__18697));
    Span4Mux_h I__3372 (
            .O(N__18703),
            .I(N__18694));
    InMux I__3371 (
            .O(N__18702),
            .I(N__18691));
    Odrv12 I__3370 (
            .O(N__18697),
            .I(M_this_vram_read_data_0));
    Odrv4 I__3369 (
            .O(N__18694),
            .I(M_this_vram_read_data_0));
    LocalMux I__3368 (
            .O(N__18691),
            .I(M_this_vram_read_data_0));
    InMux I__3367 (
            .O(N__18684),
            .I(N__18681));
    LocalMux I__3366 (
            .O(N__18681),
            .I(N__18678));
    Span4Mux_h I__3365 (
            .O(N__18678),
            .I(N__18675));
    Odrv4 I__3364 (
            .O(N__18675),
            .I(\this_vga_ramdac.m16 ));
    InMux I__3363 (
            .O(N__18672),
            .I(N__18669));
    LocalMux I__3362 (
            .O(N__18669),
            .I(\this_reset_cond.M_stage_qZ0Z_5 ));
    InMux I__3361 (
            .O(N__18666),
            .I(N__18663));
    LocalMux I__3360 (
            .O(N__18663),
            .I(N__18660));
    Odrv4 I__3359 (
            .O(N__18660),
            .I(\this_reset_cond.M_stage_qZ0Z_8 ));
    InMux I__3358 (
            .O(N__18657),
            .I(N__18654));
    LocalMux I__3357 (
            .O(N__18654),
            .I(\this_reset_cond.M_stage_qZ0Z_6 ));
    InMux I__3356 (
            .O(N__18651),
            .I(N__18648));
    LocalMux I__3355 (
            .O(N__18648),
            .I(\this_reset_cond.M_stage_qZ0Z_7 ));
    InMux I__3354 (
            .O(N__18645),
            .I(N__18641));
    InMux I__3353 (
            .O(N__18644),
            .I(N__18638));
    LocalMux I__3352 (
            .O(N__18641),
            .I(\this_ppu.M_count_qZ0Z_7 ));
    LocalMux I__3351 (
            .O(N__18638),
            .I(\this_ppu.M_count_qZ0Z_7 ));
    InMux I__3350 (
            .O(N__18633),
            .I(N__18630));
    LocalMux I__3349 (
            .O(N__18630),
            .I(\this_ppu.M_count_d_1_sqmuxa_1_i_a2_3 ));
    InMux I__3348 (
            .O(N__18627),
            .I(N__18624));
    LocalMux I__3347 (
            .O(N__18624),
            .I(N__18621));
    Odrv4 I__3346 (
            .O(N__18621),
            .I(M_this_state_qc_3_1));
    CascadeMux I__3345 (
            .O(N__18618),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_4_cascade_ ));
    CascadeMux I__3344 (
            .O(N__18615),
            .I(N__18612));
    InMux I__3343 (
            .O(N__18612),
            .I(N__18606));
    InMux I__3342 (
            .O(N__18611),
            .I(N__18599));
    InMux I__3341 (
            .O(N__18610),
            .I(N__18599));
    InMux I__3340 (
            .O(N__18609),
            .I(N__18599));
    LocalMux I__3339 (
            .O(N__18606),
            .I(N__18596));
    LocalMux I__3338 (
            .O(N__18599),
            .I(N__18593));
    Odrv4 I__3337 (
            .O(N__18596),
            .I(N_465_0));
    Odrv12 I__3336 (
            .O(N__18593),
            .I(N_465_0));
    InMux I__3335 (
            .O(N__18588),
            .I(N__18580));
    InMux I__3334 (
            .O(N__18587),
            .I(N__18580));
    InMux I__3333 (
            .O(N__18586),
            .I(N__18576));
    InMux I__3332 (
            .O(N__18585),
            .I(N__18573));
    LocalMux I__3331 (
            .O(N__18580),
            .I(N__18570));
    CascadeMux I__3330 (
            .O(N__18579),
            .I(N__18561));
    LocalMux I__3329 (
            .O(N__18576),
            .I(N__18555));
    LocalMux I__3328 (
            .O(N__18573),
            .I(N__18552));
    Span4Mux_h I__3327 (
            .O(N__18570),
            .I(N__18549));
    InMux I__3326 (
            .O(N__18569),
            .I(N__18546));
    InMux I__3325 (
            .O(N__18568),
            .I(N__18539));
    InMux I__3324 (
            .O(N__18567),
            .I(N__18539));
    InMux I__3323 (
            .O(N__18566),
            .I(N__18539));
    InMux I__3322 (
            .O(N__18565),
            .I(N__18534));
    InMux I__3321 (
            .O(N__18564),
            .I(N__18534));
    InMux I__3320 (
            .O(N__18561),
            .I(N__18525));
    InMux I__3319 (
            .O(N__18560),
            .I(N__18525));
    InMux I__3318 (
            .O(N__18559),
            .I(N__18525));
    InMux I__3317 (
            .O(N__18558),
            .I(N__18525));
    Odrv12 I__3316 (
            .O(N__18555),
            .I(N_610_0_i));
    Odrv4 I__3315 (
            .O(N__18552),
            .I(N_610_0_i));
    Odrv4 I__3314 (
            .O(N__18549),
            .I(N_610_0_i));
    LocalMux I__3313 (
            .O(N__18546),
            .I(N_610_0_i));
    LocalMux I__3312 (
            .O(N__18539),
            .I(N_610_0_i));
    LocalMux I__3311 (
            .O(N__18534),
            .I(N_610_0_i));
    LocalMux I__3310 (
            .O(N__18525),
            .I(N_610_0_i));
    CascadeMux I__3309 (
            .O(N__18510),
            .I(N__18507));
    InMux I__3308 (
            .O(N__18507),
            .I(N__18504));
    LocalMux I__3307 (
            .O(N__18504),
            .I(N__18501));
    Odrv4 I__3306 (
            .O(N__18501),
            .I(M_this_data_count_q_cry_0_THRU_CO));
    CEMux I__3305 (
            .O(N__18498),
            .I(N__18495));
    LocalMux I__3304 (
            .O(N__18495),
            .I(N__18492));
    Span4Mux_v I__3303 (
            .O(N__18492),
            .I(N__18488));
    CEMux I__3302 (
            .O(N__18491),
            .I(N__18485));
    Span4Mux_v I__3301 (
            .O(N__18488),
            .I(N__18478));
    LocalMux I__3300 (
            .O(N__18485),
            .I(N__18478));
    CEMux I__3299 (
            .O(N__18484),
            .I(N__18473));
    CEMux I__3298 (
            .O(N__18483),
            .I(N__18470));
    Span4Mux_v I__3297 (
            .O(N__18478),
            .I(N__18467));
    CEMux I__3296 (
            .O(N__18477),
            .I(N__18464));
    CEMux I__3295 (
            .O(N__18476),
            .I(N__18461));
    LocalMux I__3294 (
            .O(N__18473),
            .I(M_this_data_count_qe_0_i));
    LocalMux I__3293 (
            .O(N__18470),
            .I(M_this_data_count_qe_0_i));
    Odrv4 I__3292 (
            .O(N__18467),
            .I(M_this_data_count_qe_0_i));
    LocalMux I__3291 (
            .O(N__18464),
            .I(M_this_data_count_qe_0_i));
    LocalMux I__3290 (
            .O(N__18461),
            .I(M_this_data_count_qe_0_i));
    CascadeMux I__3289 (
            .O(N__18450),
            .I(N__18446));
    InMux I__3288 (
            .O(N__18449),
            .I(N__18442));
    InMux I__3287 (
            .O(N__18446),
            .I(N__18439));
    InMux I__3286 (
            .O(N__18445),
            .I(N__18436));
    LocalMux I__3285 (
            .O(N__18442),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__3284 (
            .O(N__18439),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__3283 (
            .O(N__18436),
            .I(M_this_data_count_qZ0Z_3));
    InMux I__3282 (
            .O(N__18429),
            .I(N__18424));
    InMux I__3281 (
            .O(N__18428),
            .I(N__18421));
    InMux I__3280 (
            .O(N__18427),
            .I(N__18418));
    LocalMux I__3279 (
            .O(N__18424),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__3278 (
            .O(N__18421),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__3277 (
            .O(N__18418),
            .I(M_this_data_count_qZ0Z_2));
    CascadeMux I__3276 (
            .O(N__18411),
            .I(N__18408));
    InMux I__3275 (
            .O(N__18408),
            .I(N__18404));
    InMux I__3274 (
            .O(N__18407),
            .I(N__18400));
    LocalMux I__3273 (
            .O(N__18404),
            .I(N__18397));
    InMux I__3272 (
            .O(N__18403),
            .I(N__18394));
    LocalMux I__3271 (
            .O(N__18400),
            .I(M_this_data_count_qZ0Z_1));
    Odrv4 I__3270 (
            .O(N__18397),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__3269 (
            .O(N__18394),
            .I(M_this_data_count_qZ0Z_1));
    InMux I__3268 (
            .O(N__18387),
            .I(N__18383));
    InMux I__3267 (
            .O(N__18386),
            .I(N__18380));
    LocalMux I__3266 (
            .O(N__18383),
            .I(N__18377));
    LocalMux I__3265 (
            .O(N__18380),
            .I(N__18374));
    Span4Mux_v I__3264 (
            .O(N__18377),
            .I(N__18371));
    Odrv4 I__3263 (
            .O(N__18374),
            .I(M_this_data_count_qZ0Z_10));
    Odrv4 I__3262 (
            .O(N__18371),
            .I(M_this_data_count_qZ0Z_10));
    InMux I__3261 (
            .O(N__18366),
            .I(N__18361));
    CascadeMux I__3260 (
            .O(N__18365),
            .I(N__18358));
    CascadeMux I__3259 (
            .O(N__18364),
            .I(N__18355));
    LocalMux I__3258 (
            .O(N__18361),
            .I(N__18352));
    InMux I__3257 (
            .O(N__18358),
            .I(N__18349));
    InMux I__3256 (
            .O(N__18355),
            .I(N__18346));
    Odrv4 I__3255 (
            .O(N__18352),
            .I(M_this_data_count_qZ0Z_11));
    LocalMux I__3254 (
            .O(N__18349),
            .I(M_this_data_count_qZ0Z_11));
    LocalMux I__3253 (
            .O(N__18346),
            .I(M_this_data_count_qZ0Z_11));
    InMux I__3252 (
            .O(N__18339),
            .I(N__18335));
    InMux I__3251 (
            .O(N__18338),
            .I(N__18331));
    LocalMux I__3250 (
            .O(N__18335),
            .I(N__18328));
    InMux I__3249 (
            .O(N__18334),
            .I(N__18325));
    LocalMux I__3248 (
            .O(N__18331),
            .I(M_this_data_count_qZ0Z_0));
    Odrv4 I__3247 (
            .O(N__18328),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__3246 (
            .O(N__18325),
            .I(M_this_data_count_qZ0Z_0));
    CascadeMux I__3245 (
            .O(N__18318),
            .I(\this_vga_signals.N_322_cascade_ ));
    CascadeMux I__3244 (
            .O(N__18315),
            .I(N__18312));
    InMux I__3243 (
            .O(N__18312),
            .I(N__18309));
    LocalMux I__3242 (
            .O(N__18309),
            .I(this_vga_signals_M_this_state_q_ns_i_o3_0_10));
    InMux I__3241 (
            .O(N__18306),
            .I(N__18299));
    InMux I__3240 (
            .O(N__18305),
            .I(N__18294));
    InMux I__3239 (
            .O(N__18304),
            .I(N__18294));
    InMux I__3238 (
            .O(N__18303),
            .I(N__18289));
    InMux I__3237 (
            .O(N__18302),
            .I(N__18289));
    LocalMux I__3236 (
            .O(N__18299),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__3235 (
            .O(N__18294),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__3234 (
            .O(N__18289),
            .I(M_this_state_qZ0Z_10));
    InMux I__3233 (
            .O(N__18282),
            .I(N__18277));
    InMux I__3232 (
            .O(N__18281),
            .I(N__18274));
    InMux I__3231 (
            .O(N__18280),
            .I(N__18271));
    LocalMux I__3230 (
            .O(N__18277),
            .I(N__18268));
    LocalMux I__3229 (
            .O(N__18274),
            .I(N_212));
    LocalMux I__3228 (
            .O(N__18271),
            .I(N_212));
    Odrv12 I__3227 (
            .O(N__18268),
            .I(N_212));
    CEMux I__3226 (
            .O(N__18261),
            .I(N__18257));
    CascadeMux I__3225 (
            .O(N__18260),
            .I(N__18252));
    LocalMux I__3224 (
            .O(N__18257),
            .I(N__18245));
    InMux I__3223 (
            .O(N__18256),
            .I(N__18242));
    InMux I__3222 (
            .O(N__18255),
            .I(N__18234));
    InMux I__3221 (
            .O(N__18252),
            .I(N__18231));
    CascadeMux I__3220 (
            .O(N__18251),
            .I(N__18228));
    CEMux I__3219 (
            .O(N__18250),
            .I(N__18225));
    InMux I__3218 (
            .O(N__18249),
            .I(N__18220));
    InMux I__3217 (
            .O(N__18248),
            .I(N__18220));
    Span4Mux_v I__3216 (
            .O(N__18245),
            .I(N__18217));
    LocalMux I__3215 (
            .O(N__18242),
            .I(N__18214));
    InMux I__3214 (
            .O(N__18241),
            .I(N__18209));
    InMux I__3213 (
            .O(N__18240),
            .I(N__18209));
    InMux I__3212 (
            .O(N__18239),
            .I(N__18206));
    InMux I__3211 (
            .O(N__18238),
            .I(N__18201));
    InMux I__3210 (
            .O(N__18237),
            .I(N__18201));
    LocalMux I__3209 (
            .O(N__18234),
            .I(N__18196));
    LocalMux I__3208 (
            .O(N__18231),
            .I(N__18196));
    InMux I__3207 (
            .O(N__18228),
            .I(N__18193));
    LocalMux I__3206 (
            .O(N__18225),
            .I(N__18188));
    LocalMux I__3205 (
            .O(N__18220),
            .I(N__18188));
    Span4Mux_v I__3204 (
            .O(N__18217),
            .I(N__18185));
    Span4Mux_h I__3203 (
            .O(N__18214),
            .I(N__18178));
    LocalMux I__3202 (
            .O(N__18209),
            .I(N__18178));
    LocalMux I__3201 (
            .O(N__18206),
            .I(N__18178));
    LocalMux I__3200 (
            .O(N__18201),
            .I(N__18175));
    Span4Mux_h I__3199 (
            .O(N__18196),
            .I(N__18172));
    LocalMux I__3198 (
            .O(N__18193),
            .I(N__18169));
    Span12Mux_h I__3197 (
            .O(N__18188),
            .I(N__18166));
    Span4Mux_h I__3196 (
            .O(N__18185),
            .I(N__18161));
    Span4Mux_v I__3195 (
            .O(N__18178),
            .I(N__18161));
    Span4Mux_v I__3194 (
            .O(N__18175),
            .I(N__18156));
    Span4Mux_h I__3193 (
            .O(N__18172),
            .I(N__18156));
    Odrv4 I__3192 (
            .O(N__18169),
            .I(N_160_0));
    Odrv12 I__3191 (
            .O(N__18166),
            .I(N_160_0));
    Odrv4 I__3190 (
            .O(N__18161),
            .I(N_160_0));
    Odrv4 I__3189 (
            .O(N__18156),
            .I(N_160_0));
    CascadeMux I__3188 (
            .O(N__18147),
            .I(N__18144));
    InMux I__3187 (
            .O(N__18144),
            .I(N__18141));
    LocalMux I__3186 (
            .O(N__18141),
            .I(\this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ));
    CascadeMux I__3185 (
            .O(N__18138),
            .I(N__18134));
    InMux I__3184 (
            .O(N__18137),
            .I(N__18130));
    InMux I__3183 (
            .O(N__18134),
            .I(N__18125));
    InMux I__3182 (
            .O(N__18133),
            .I(N__18125));
    LocalMux I__3181 (
            .O(N__18130),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    LocalMux I__3180 (
            .O(N__18125),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    CascadeMux I__3179 (
            .O(N__18120),
            .I(N__18117));
    InMux I__3178 (
            .O(N__18117),
            .I(N__18112));
    InMux I__3177 (
            .O(N__18116),
            .I(N__18107));
    InMux I__3176 (
            .O(N__18115),
            .I(N__18107));
    LocalMux I__3175 (
            .O(N__18112),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    LocalMux I__3174 (
            .O(N__18107),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    CascadeMux I__3173 (
            .O(N__18102),
            .I(N__18099));
    InMux I__3172 (
            .O(N__18099),
            .I(N__18094));
    CascadeMux I__3171 (
            .O(N__18098),
            .I(N__18091));
    CascadeMux I__3170 (
            .O(N__18097),
            .I(N__18088));
    LocalMux I__3169 (
            .O(N__18094),
            .I(N__18085));
    InMux I__3168 (
            .O(N__18091),
            .I(N__18080));
    InMux I__3167 (
            .O(N__18088),
            .I(N__18080));
    Odrv4 I__3166 (
            .O(N__18085),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    LocalMux I__3165 (
            .O(N__18080),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    CascadeMux I__3164 (
            .O(N__18075),
            .I(N__18072));
    InMux I__3163 (
            .O(N__18072),
            .I(N__18067));
    InMux I__3162 (
            .O(N__18071),
            .I(N__18062));
    InMux I__3161 (
            .O(N__18070),
            .I(N__18062));
    LocalMux I__3160 (
            .O(N__18067),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    LocalMux I__3159 (
            .O(N__18062),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    InMux I__3158 (
            .O(N__18057),
            .I(N__18054));
    LocalMux I__3157 (
            .O(N__18054),
            .I(N__18051));
    Odrv4 I__3156 (
            .O(N__18051),
            .I(\this_ppu.M_count_d_1_sqmuxa_1_i_a2_4 ));
    InMux I__3155 (
            .O(N__18048),
            .I(N__18045));
    LocalMux I__3154 (
            .O(N__18045),
            .I(N__18042));
    Span4Mux_h I__3153 (
            .O(N__18042),
            .I(N__18039));
    Odrv4 I__3152 (
            .O(N__18039),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    CascadeMux I__3151 (
            .O(N__18036),
            .I(\this_vga_signals.un20_i_a2_sxZ0Z_3_cascade_ ));
    InMux I__3150 (
            .O(N__18033),
            .I(\this_ppu.un1_M_count_q_1_cry_1_s1 ));
    InMux I__3149 (
            .O(N__18030),
            .I(\this_ppu.un1_M_count_q_1_cry_2_s1 ));
    InMux I__3148 (
            .O(N__18027),
            .I(\this_ppu.un1_M_count_q_1_cry_3_s1 ));
    InMux I__3147 (
            .O(N__18024),
            .I(\this_ppu.un1_M_count_q_1_cry_4_s1 ));
    SRMux I__3146 (
            .O(N__18021),
            .I(N__18016));
    SRMux I__3145 (
            .O(N__18020),
            .I(N__18013));
    SRMux I__3144 (
            .O(N__18019),
            .I(N__18007));
    LocalMux I__3143 (
            .O(N__18016),
            .I(N__18001));
    LocalMux I__3142 (
            .O(N__18013),
            .I(N__18001));
    SRMux I__3141 (
            .O(N__18012),
            .I(N__17998));
    IoInMux I__3140 (
            .O(N__18011),
            .I(N__17993));
    SRMux I__3139 (
            .O(N__18010),
            .I(N__17986));
    LocalMux I__3138 (
            .O(N__18007),
            .I(N__17983));
    SRMux I__3137 (
            .O(N__18006),
            .I(N__17980));
    Span4Mux_v I__3136 (
            .O(N__18001),
            .I(N__17975));
    LocalMux I__3135 (
            .O(N__17998),
            .I(N__17975));
    SRMux I__3134 (
            .O(N__17997),
            .I(N__17972));
    SRMux I__3133 (
            .O(N__17996),
            .I(N__17969));
    LocalMux I__3132 (
            .O(N__17993),
            .I(N__17965));
    SRMux I__3131 (
            .O(N__17992),
            .I(N__17960));
    SRMux I__3130 (
            .O(N__17991),
            .I(N__17953));
    IoInMux I__3129 (
            .O(N__17990),
            .I(N__17949));
    SRMux I__3128 (
            .O(N__17989),
            .I(N__17944));
    LocalMux I__3127 (
            .O(N__17986),
            .I(N__17935));
    Span4Mux_h I__3126 (
            .O(N__17983),
            .I(N__17935));
    LocalMux I__3125 (
            .O(N__17980),
            .I(N__17935));
    Span4Mux_h I__3124 (
            .O(N__17975),
            .I(N__17927));
    LocalMux I__3123 (
            .O(N__17972),
            .I(N__17927));
    LocalMux I__3122 (
            .O(N__17969),
            .I(N__17927));
    SRMux I__3121 (
            .O(N__17968),
            .I(N__17924));
    IoSpan4Mux I__3120 (
            .O(N__17965),
            .I(N__17919));
    SRMux I__3119 (
            .O(N__17964),
            .I(N__17916));
    SRMux I__3118 (
            .O(N__17963),
            .I(N__17913));
    LocalMux I__3117 (
            .O(N__17960),
            .I(N__17910));
    SRMux I__3116 (
            .O(N__17959),
            .I(N__17907));
    SRMux I__3115 (
            .O(N__17958),
            .I(N__17902));
    SRMux I__3114 (
            .O(N__17957),
            .I(N__17899));
    SRMux I__3113 (
            .O(N__17956),
            .I(N__17891));
    LocalMux I__3112 (
            .O(N__17953),
            .I(N__17888));
    SRMux I__3111 (
            .O(N__17952),
            .I(N__17885));
    LocalMux I__3110 (
            .O(N__17949),
            .I(N__17881));
    SRMux I__3109 (
            .O(N__17948),
            .I(N__17878));
    SRMux I__3108 (
            .O(N__17947),
            .I(N__17875));
    LocalMux I__3107 (
            .O(N__17944),
            .I(N__17872));
    SRMux I__3106 (
            .O(N__17943),
            .I(N__17869));
    SRMux I__3105 (
            .O(N__17942),
            .I(N__17866));
    Span4Mux_v I__3104 (
            .O(N__17935),
            .I(N__17861));
    SRMux I__3103 (
            .O(N__17934),
            .I(N__17858));
    Span4Mux_v I__3102 (
            .O(N__17927),
            .I(N__17853));
    LocalMux I__3101 (
            .O(N__17924),
            .I(N__17853));
    SRMux I__3100 (
            .O(N__17923),
            .I(N__17850));
    SRMux I__3099 (
            .O(N__17922),
            .I(N__17846));
    Span4Mux_s3_h I__3098 (
            .O(N__17919),
            .I(N__17843));
    LocalMux I__3097 (
            .O(N__17916),
            .I(N__17838));
    LocalMux I__3096 (
            .O(N__17913),
            .I(N__17838));
    Span4Mux_v I__3095 (
            .O(N__17910),
            .I(N__17833));
    LocalMux I__3094 (
            .O(N__17907),
            .I(N__17833));
    SRMux I__3093 (
            .O(N__17906),
            .I(N__17830));
    SRMux I__3092 (
            .O(N__17905),
            .I(N__17827));
    LocalMux I__3091 (
            .O(N__17902),
            .I(N__17824));
    LocalMux I__3090 (
            .O(N__17899),
            .I(N__17821));
    SRMux I__3089 (
            .O(N__17898),
            .I(N__17818));
    CascadeMux I__3088 (
            .O(N__17897),
            .I(N__17814));
    CascadeMux I__3087 (
            .O(N__17896),
            .I(N__17811));
    CascadeMux I__3086 (
            .O(N__17895),
            .I(N__17807));
    SRMux I__3085 (
            .O(N__17894),
            .I(N__17800));
    LocalMux I__3084 (
            .O(N__17891),
            .I(N__17793));
    Span4Mux_h I__3083 (
            .O(N__17888),
            .I(N__17793));
    LocalMux I__3082 (
            .O(N__17885),
            .I(N__17793));
    SRMux I__3081 (
            .O(N__17884),
            .I(N__17790));
    IoSpan4Mux I__3080 (
            .O(N__17881),
            .I(N__17787));
    LocalMux I__3079 (
            .O(N__17878),
            .I(N__17782));
    LocalMux I__3078 (
            .O(N__17875),
            .I(N__17782));
    Span4Mux_v I__3077 (
            .O(N__17872),
            .I(N__17775));
    LocalMux I__3076 (
            .O(N__17869),
            .I(N__17775));
    LocalMux I__3075 (
            .O(N__17866),
            .I(N__17775));
    SRMux I__3074 (
            .O(N__17865),
            .I(N__17772));
    SRMux I__3073 (
            .O(N__17864),
            .I(N__17769));
    Span4Mux_h I__3072 (
            .O(N__17861),
            .I(N__17756));
    LocalMux I__3071 (
            .O(N__17858),
            .I(N__17756));
    Span4Mux_v I__3070 (
            .O(N__17853),
            .I(N__17756));
    LocalMux I__3069 (
            .O(N__17850),
            .I(N__17756));
    SRMux I__3068 (
            .O(N__17849),
            .I(N__17753));
    LocalMux I__3067 (
            .O(N__17846),
            .I(N__17749));
    Span4Mux_h I__3066 (
            .O(N__17843),
            .I(N__17740));
    Span4Mux_v I__3065 (
            .O(N__17838),
            .I(N__17740));
    Span4Mux_v I__3064 (
            .O(N__17833),
            .I(N__17740));
    LocalMux I__3063 (
            .O(N__17830),
            .I(N__17740));
    LocalMux I__3062 (
            .O(N__17827),
            .I(N__17735));
    Span4Mux_h I__3061 (
            .O(N__17824),
            .I(N__17732));
    Span4Mux_h I__3060 (
            .O(N__17821),
            .I(N__17729));
    LocalMux I__3059 (
            .O(N__17818),
            .I(N__17726));
    InMux I__3058 (
            .O(N__17817),
            .I(N__17715));
    InMux I__3057 (
            .O(N__17814),
            .I(N__17715));
    InMux I__3056 (
            .O(N__17811),
            .I(N__17715));
    InMux I__3055 (
            .O(N__17810),
            .I(N__17715));
    InMux I__3054 (
            .O(N__17807),
            .I(N__17715));
    CascadeMux I__3053 (
            .O(N__17806),
            .I(N__17710));
    CascadeMux I__3052 (
            .O(N__17805),
            .I(N__17706));
    CascadeMux I__3051 (
            .O(N__17804),
            .I(N__17702));
    SRMux I__3050 (
            .O(N__17803),
            .I(N__17699));
    LocalMux I__3049 (
            .O(N__17800),
            .I(N__17692));
    Span4Mux_v I__3048 (
            .O(N__17793),
            .I(N__17692));
    LocalMux I__3047 (
            .O(N__17790),
            .I(N__17692));
    Span4Mux_s0_h I__3046 (
            .O(N__17787),
            .I(N__17689));
    Span4Mux_v I__3045 (
            .O(N__17782),
            .I(N__17680));
    Span4Mux_v I__3044 (
            .O(N__17775),
            .I(N__17680));
    LocalMux I__3043 (
            .O(N__17772),
            .I(N__17680));
    LocalMux I__3042 (
            .O(N__17769),
            .I(N__17680));
    SRMux I__3041 (
            .O(N__17768),
            .I(N__17677));
    SRMux I__3040 (
            .O(N__17767),
            .I(N__17674));
    SRMux I__3039 (
            .O(N__17766),
            .I(N__17671));
    SRMux I__3038 (
            .O(N__17765),
            .I(N__17668));
    Span4Mux_v I__3037 (
            .O(N__17756),
            .I(N__17665));
    LocalMux I__3036 (
            .O(N__17753),
            .I(N__17662));
    SRMux I__3035 (
            .O(N__17752),
            .I(N__17659));
    Span4Mux_v I__3034 (
            .O(N__17749),
            .I(N__17654));
    Span4Mux_v I__3033 (
            .O(N__17740),
            .I(N__17654));
    SRMux I__3032 (
            .O(N__17739),
            .I(N__17651));
    SRMux I__3031 (
            .O(N__17738),
            .I(N__17648));
    Span4Mux_h I__3030 (
            .O(N__17735),
            .I(N__17645));
    Span4Mux_h I__3029 (
            .O(N__17732),
            .I(N__17642));
    Span4Mux_v I__3028 (
            .O(N__17729),
            .I(N__17639));
    Span4Mux_h I__3027 (
            .O(N__17726),
            .I(N__17636));
    LocalMux I__3026 (
            .O(N__17715),
            .I(N__17633));
    InMux I__3025 (
            .O(N__17714),
            .I(N__17618));
    InMux I__3024 (
            .O(N__17713),
            .I(N__17618));
    InMux I__3023 (
            .O(N__17710),
            .I(N__17618));
    InMux I__3022 (
            .O(N__17709),
            .I(N__17618));
    InMux I__3021 (
            .O(N__17706),
            .I(N__17618));
    InMux I__3020 (
            .O(N__17705),
            .I(N__17618));
    InMux I__3019 (
            .O(N__17702),
            .I(N__17618));
    LocalMux I__3018 (
            .O(N__17699),
            .I(N__17615));
    Span4Mux_v I__3017 (
            .O(N__17692),
            .I(N__17612));
    Span4Mux_h I__3016 (
            .O(N__17689),
            .I(N__17605));
    Span4Mux_v I__3015 (
            .O(N__17680),
            .I(N__17605));
    LocalMux I__3014 (
            .O(N__17677),
            .I(N__17605));
    LocalMux I__3013 (
            .O(N__17674),
            .I(N__17595));
    LocalMux I__3012 (
            .O(N__17671),
            .I(N__17595));
    LocalMux I__3011 (
            .O(N__17668),
            .I(N__17595));
    Sp12to4 I__3010 (
            .O(N__17665),
            .I(N__17592));
    Span12Mux_s6_v I__3009 (
            .O(N__17662),
            .I(N__17581));
    LocalMux I__3008 (
            .O(N__17659),
            .I(N__17581));
    Sp12to4 I__3007 (
            .O(N__17654),
            .I(N__17581));
    LocalMux I__3006 (
            .O(N__17651),
            .I(N__17581));
    LocalMux I__3005 (
            .O(N__17648),
            .I(N__17581));
    Span4Mux_h I__3004 (
            .O(N__17645),
            .I(N__17578));
    Span4Mux_v I__3003 (
            .O(N__17642),
            .I(N__17571));
    Span4Mux_h I__3002 (
            .O(N__17639),
            .I(N__17571));
    Span4Mux_h I__3001 (
            .O(N__17636),
            .I(N__17571));
    Span4Mux_v I__3000 (
            .O(N__17633),
            .I(N__17566));
    LocalMux I__2999 (
            .O(N__17618),
            .I(N__17566));
    Span4Mux_v I__2998 (
            .O(N__17615),
            .I(N__17559));
    Span4Mux_h I__2997 (
            .O(N__17612),
            .I(N__17559));
    Span4Mux_h I__2996 (
            .O(N__17605),
            .I(N__17559));
    CascadeMux I__2995 (
            .O(N__17604),
            .I(N__17555));
    CascadeMux I__2994 (
            .O(N__17603),
            .I(N__17551));
    CascadeMux I__2993 (
            .O(N__17602),
            .I(N__17547));
    Span12Mux_v I__2992 (
            .O(N__17595),
            .I(N__17540));
    Span12Mux_s7_h I__2991 (
            .O(N__17592),
            .I(N__17540));
    Span12Mux_v I__2990 (
            .O(N__17581),
            .I(N__17540));
    Span4Mux_h I__2989 (
            .O(N__17578),
            .I(N__17537));
    Span4Mux_h I__2988 (
            .O(N__17571),
            .I(N__17534));
    Span4Mux_v I__2987 (
            .O(N__17566),
            .I(N__17531));
    Span4Mux_h I__2986 (
            .O(N__17559),
            .I(N__17528));
    InMux I__2985 (
            .O(N__17558),
            .I(N__17515));
    InMux I__2984 (
            .O(N__17555),
            .I(N__17515));
    InMux I__2983 (
            .O(N__17554),
            .I(N__17515));
    InMux I__2982 (
            .O(N__17551),
            .I(N__17515));
    InMux I__2981 (
            .O(N__17550),
            .I(N__17515));
    InMux I__2980 (
            .O(N__17547),
            .I(N__17515));
    Odrv12 I__2979 (
            .O(N__17540),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2978 (
            .O(N__17537),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2977 (
            .O(N__17534),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2976 (
            .O(N__17531),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2975 (
            .O(N__17528),
            .I(CONSTANT_ONE_NET));
    LocalMux I__2974 (
            .O(N__17515),
            .I(CONSTANT_ONE_NET));
    InMux I__2973 (
            .O(N__17502),
            .I(\this_ppu.un1_M_count_q_1_cry_5_s1 ));
    InMux I__2972 (
            .O(N__17499),
            .I(\this_ppu.un1_M_count_q_1_cry_6_s1 ));
    InMux I__2971 (
            .O(N__17496),
            .I(N__17493));
    LocalMux I__2970 (
            .O(N__17493),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_7 ));
    InMux I__2969 (
            .O(N__17490),
            .I(N__17487));
    LocalMux I__2968 (
            .O(N__17487),
            .I(\this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ));
    InMux I__2967 (
            .O(N__17484),
            .I(N__17481));
    LocalMux I__2966 (
            .O(N__17481),
            .I(\this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ));
    InMux I__2965 (
            .O(N__17478),
            .I(N__17475));
    LocalMux I__2964 (
            .O(N__17475),
            .I(N__17472));
    Odrv12 I__2963 (
            .O(N__17472),
            .I(\this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ));
    CascadeMux I__2962 (
            .O(N__17469),
            .I(N__17466));
    InMux I__2961 (
            .O(N__17466),
            .I(N__17463));
    LocalMux I__2960 (
            .O(N__17463),
            .I(M_this_data_count_q_cry_1_THRU_CO));
    InMux I__2959 (
            .O(N__17460),
            .I(N__17457));
    LocalMux I__2958 (
            .O(N__17457),
            .I(M_this_data_count_q_cry_8_THRU_CO));
    CascadeMux I__2957 (
            .O(N__17454),
            .I(N__17450));
    InMux I__2956 (
            .O(N__17453),
            .I(N__17446));
    InMux I__2955 (
            .O(N__17450),
            .I(N__17443));
    InMux I__2954 (
            .O(N__17449),
            .I(N__17440));
    LocalMux I__2953 (
            .O(N__17446),
            .I(M_this_data_count_qZ0Z_9));
    LocalMux I__2952 (
            .O(N__17443),
            .I(M_this_data_count_qZ0Z_9));
    LocalMux I__2951 (
            .O(N__17440),
            .I(M_this_data_count_qZ0Z_9));
    InMux I__2950 (
            .O(N__17433),
            .I(N__17430));
    LocalMux I__2949 (
            .O(N__17430),
            .I(N__17427));
    Span4Mux_v I__2948 (
            .O(N__17427),
            .I(N__17424));
    Span4Mux_v I__2947 (
            .O(N__17424),
            .I(N__17421));
    Span4Mux_h I__2946 (
            .O(N__17421),
            .I(N__17418));
    Span4Mux_h I__2945 (
            .O(N__17418),
            .I(N__17415));
    Odrv4 I__2944 (
            .O(N__17415),
            .I(M_this_map_ram_read_data_1));
    CascadeMux I__2943 (
            .O(N__17412),
            .I(N__17408));
    CascadeMux I__2942 (
            .O(N__17411),
            .I(N__17402));
    InMux I__2941 (
            .O(N__17408),
            .I(N__17396));
    CascadeMux I__2940 (
            .O(N__17407),
            .I(N__17393));
    CascadeMux I__2939 (
            .O(N__17406),
            .I(N__17388));
    CascadeMux I__2938 (
            .O(N__17405),
            .I(N__17385));
    InMux I__2937 (
            .O(N__17402),
            .I(N__17381));
    CascadeMux I__2936 (
            .O(N__17401),
            .I(N__17377));
    CascadeMux I__2935 (
            .O(N__17400),
            .I(N__17374));
    CascadeMux I__2934 (
            .O(N__17399),
            .I(N__17371));
    LocalMux I__2933 (
            .O(N__17396),
            .I(N__17368));
    InMux I__2932 (
            .O(N__17393),
            .I(N__17365));
    CascadeMux I__2931 (
            .O(N__17392),
            .I(N__17362));
    CascadeMux I__2930 (
            .O(N__17391),
            .I(N__17359));
    InMux I__2929 (
            .O(N__17388),
            .I(N__17355));
    InMux I__2928 (
            .O(N__17385),
            .I(N__17352));
    CascadeMux I__2927 (
            .O(N__17384),
            .I(N__17349));
    LocalMux I__2926 (
            .O(N__17381),
            .I(N__17344));
    CascadeMux I__2925 (
            .O(N__17380),
            .I(N__17341));
    InMux I__2924 (
            .O(N__17377),
            .I(N__17338));
    InMux I__2923 (
            .O(N__17374),
            .I(N__17335));
    InMux I__2922 (
            .O(N__17371),
            .I(N__17332));
    Span4Mux_s2_v I__2921 (
            .O(N__17368),
            .I(N__17327));
    LocalMux I__2920 (
            .O(N__17365),
            .I(N__17327));
    InMux I__2919 (
            .O(N__17362),
            .I(N__17324));
    InMux I__2918 (
            .O(N__17359),
            .I(N__17321));
    CascadeMux I__2917 (
            .O(N__17358),
            .I(N__17318));
    LocalMux I__2916 (
            .O(N__17355),
            .I(N__17313));
    LocalMux I__2915 (
            .O(N__17352),
            .I(N__17313));
    InMux I__2914 (
            .O(N__17349),
            .I(N__17310));
    CascadeMux I__2913 (
            .O(N__17348),
            .I(N__17307));
    CascadeMux I__2912 (
            .O(N__17347),
            .I(N__17304));
    Span4Mux_v I__2911 (
            .O(N__17344),
            .I(N__17301));
    InMux I__2910 (
            .O(N__17341),
            .I(N__17298));
    LocalMux I__2909 (
            .O(N__17338),
            .I(N__17295));
    LocalMux I__2908 (
            .O(N__17335),
            .I(N__17292));
    LocalMux I__2907 (
            .O(N__17332),
            .I(N__17289));
    Span4Mux_v I__2906 (
            .O(N__17327),
            .I(N__17284));
    LocalMux I__2905 (
            .O(N__17324),
            .I(N__17284));
    LocalMux I__2904 (
            .O(N__17321),
            .I(N__17281));
    InMux I__2903 (
            .O(N__17318),
            .I(N__17278));
    Span4Mux_v I__2902 (
            .O(N__17313),
            .I(N__17272));
    LocalMux I__2901 (
            .O(N__17310),
            .I(N__17272));
    InMux I__2900 (
            .O(N__17307),
            .I(N__17269));
    InMux I__2899 (
            .O(N__17304),
            .I(N__17266));
    Sp12to4 I__2898 (
            .O(N__17301),
            .I(N__17261));
    LocalMux I__2897 (
            .O(N__17298),
            .I(N__17261));
    Span4Mux_h I__2896 (
            .O(N__17295),
            .I(N__17258));
    Span4Mux_h I__2895 (
            .O(N__17292),
            .I(N__17255));
    Span4Mux_h I__2894 (
            .O(N__17289),
            .I(N__17252));
    Span4Mux_v I__2893 (
            .O(N__17284),
            .I(N__17245));
    Span4Mux_h I__2892 (
            .O(N__17281),
            .I(N__17245));
    LocalMux I__2891 (
            .O(N__17278),
            .I(N__17245));
    CascadeMux I__2890 (
            .O(N__17277),
            .I(N__17242));
    Span4Mux_v I__2889 (
            .O(N__17272),
            .I(N__17237));
    LocalMux I__2888 (
            .O(N__17269),
            .I(N__17237));
    LocalMux I__2887 (
            .O(N__17266),
            .I(N__17234));
    Span12Mux_h I__2886 (
            .O(N__17261),
            .I(N__17231));
    Sp12to4 I__2885 (
            .O(N__17258),
            .I(N__17224));
    Sp12to4 I__2884 (
            .O(N__17255),
            .I(N__17224));
    Sp12to4 I__2883 (
            .O(N__17252),
            .I(N__17224));
    Span4Mux_v I__2882 (
            .O(N__17245),
            .I(N__17221));
    InMux I__2881 (
            .O(N__17242),
            .I(N__17218));
    Span4Mux_h I__2880 (
            .O(N__17237),
            .I(N__17215));
    Span12Mux_h I__2879 (
            .O(N__17234),
            .I(N__17212));
    Span12Mux_v I__2878 (
            .O(N__17231),
            .I(N__17203));
    Span12Mux_v I__2877 (
            .O(N__17224),
            .I(N__17203));
    Sp12to4 I__2876 (
            .O(N__17221),
            .I(N__17203));
    LocalMux I__2875 (
            .O(N__17218),
            .I(N__17203));
    Span4Mux_h I__2874 (
            .O(N__17215),
            .I(N__17200));
    Odrv12 I__2873 (
            .O(N__17212),
            .I(M_this_ppu_sprites_addr_7));
    Odrv12 I__2872 (
            .O(N__17203),
            .I(M_this_ppu_sprites_addr_7));
    Odrv4 I__2871 (
            .O(N__17200),
            .I(M_this_ppu_sprites_addr_7));
    CascadeMux I__2870 (
            .O(N__17193),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_7_cascade_ ));
    InMux I__2869 (
            .O(N__17190),
            .I(N__17186));
    InMux I__2868 (
            .O(N__17189),
            .I(N__17183));
    LocalMux I__2867 (
            .O(N__17186),
            .I(\this_vga_signals.un4_lvisibility_1 ));
    LocalMux I__2866 (
            .O(N__17183),
            .I(\this_vga_signals.un4_lvisibility_1 ));
    CascadeMux I__2865 (
            .O(N__17178),
            .I(N__17173));
    InMux I__2864 (
            .O(N__17177),
            .I(N__17163));
    InMux I__2863 (
            .O(N__17176),
            .I(N__17160));
    InMux I__2862 (
            .O(N__17173),
            .I(N__17157));
    InMux I__2861 (
            .O(N__17172),
            .I(N__17154));
    InMux I__2860 (
            .O(N__17171),
            .I(N__17151));
    InMux I__2859 (
            .O(N__17170),
            .I(N__17146));
    InMux I__2858 (
            .O(N__17169),
            .I(N__17146));
    InMux I__2857 (
            .O(N__17168),
            .I(N__17143));
    InMux I__2856 (
            .O(N__17167),
            .I(N__17140));
    InMux I__2855 (
            .O(N__17166),
            .I(N__17137));
    LocalMux I__2854 (
            .O(N__17163),
            .I(N__17129));
    LocalMux I__2853 (
            .O(N__17160),
            .I(N__17129));
    LocalMux I__2852 (
            .O(N__17157),
            .I(N__17129));
    LocalMux I__2851 (
            .O(N__17154),
            .I(N__17126));
    LocalMux I__2850 (
            .O(N__17151),
            .I(N__17123));
    LocalMux I__2849 (
            .O(N__17146),
            .I(N__17111));
    LocalMux I__2848 (
            .O(N__17143),
            .I(N__17111));
    LocalMux I__2847 (
            .O(N__17140),
            .I(N__17111));
    LocalMux I__2846 (
            .O(N__17137),
            .I(N__17111));
    InMux I__2845 (
            .O(N__17136),
            .I(N__17108));
    Span4Mux_v I__2844 (
            .O(N__17129),
            .I(N__17105));
    Span4Mux_v I__2843 (
            .O(N__17126),
            .I(N__17100));
    Span4Mux_h I__2842 (
            .O(N__17123),
            .I(N__17100));
    InMux I__2841 (
            .O(N__17122),
            .I(N__17095));
    InMux I__2840 (
            .O(N__17121),
            .I(N__17095));
    InMux I__2839 (
            .O(N__17120),
            .I(N__17092));
    Span4Mux_v I__2838 (
            .O(N__17111),
            .I(N__17087));
    LocalMux I__2837 (
            .O(N__17108),
            .I(N__17087));
    Span4Mux_h I__2836 (
            .O(N__17105),
            .I(N__17084));
    Odrv4 I__2835 (
            .O(N__17100),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2834 (
            .O(N__17095),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2833 (
            .O(N__17092),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2832 (
            .O(N__17087),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2831 (
            .O(N__17084),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    InMux I__2830 (
            .O(N__17073),
            .I(N__17069));
    InMux I__2829 (
            .O(N__17072),
            .I(N__17063));
    LocalMux I__2828 (
            .O(N__17069),
            .I(N__17060));
    InMux I__2827 (
            .O(N__17068),
            .I(N__17057));
    InMux I__2826 (
            .O(N__17067),
            .I(N__17052));
    InMux I__2825 (
            .O(N__17066),
            .I(N__17052));
    LocalMux I__2824 (
            .O(N__17063),
            .I(N__17042));
    Span4Mux_v I__2823 (
            .O(N__17060),
            .I(N__17042));
    LocalMux I__2822 (
            .O(N__17057),
            .I(N__17039));
    LocalMux I__2821 (
            .O(N__17052),
            .I(N__17036));
    InMux I__2820 (
            .O(N__17051),
            .I(N__17031));
    InMux I__2819 (
            .O(N__17050),
            .I(N__17031));
    InMux I__2818 (
            .O(N__17049),
            .I(N__17028));
    InMux I__2817 (
            .O(N__17048),
            .I(N__17025));
    InMux I__2816 (
            .O(N__17047),
            .I(N__17022));
    Span4Mux_h I__2815 (
            .O(N__17042),
            .I(N__17011));
    Span4Mux_v I__2814 (
            .O(N__17039),
            .I(N__17011));
    Sp12to4 I__2813 (
            .O(N__17036),
            .I(N__17004));
    LocalMux I__2812 (
            .O(N__17031),
            .I(N__17004));
    LocalMux I__2811 (
            .O(N__17028),
            .I(N__17004));
    LocalMux I__2810 (
            .O(N__17025),
            .I(N__16999));
    LocalMux I__2809 (
            .O(N__17022),
            .I(N__16999));
    InMux I__2808 (
            .O(N__17021),
            .I(N__16994));
    InMux I__2807 (
            .O(N__17020),
            .I(N__16994));
    InMux I__2806 (
            .O(N__17019),
            .I(N__16991));
    InMux I__2805 (
            .O(N__17018),
            .I(N__16988));
    InMux I__2804 (
            .O(N__17017),
            .I(N__16983));
    InMux I__2803 (
            .O(N__17016),
            .I(N__16983));
    Odrv4 I__2802 (
            .O(N__17011),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv12 I__2801 (
            .O(N__17004),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv12 I__2800 (
            .O(N__16999),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2799 (
            .O(N__16994),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2798 (
            .O(N__16991),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2797 (
            .O(N__16988),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2796 (
            .O(N__16983),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    InMux I__2795 (
            .O(N__16968),
            .I(\this_ppu.un1_M_count_q_1_cry_0_s1 ));
    InMux I__2794 (
            .O(N__16965),
            .I(N__16961));
    InMux I__2793 (
            .O(N__16964),
            .I(N__16958));
    LocalMux I__2792 (
            .O(N__16961),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__2791 (
            .O(N__16958),
            .I(M_this_data_count_qZ0Z_6));
    InMux I__2790 (
            .O(N__16953),
            .I(N__16950));
    LocalMux I__2789 (
            .O(N__16950),
            .I(M_this_data_count_q_cry_3_THRU_CO));
    InMux I__2788 (
            .O(N__16947),
            .I(N__16942));
    InMux I__2787 (
            .O(N__16946),
            .I(N__16937));
    InMux I__2786 (
            .O(N__16945),
            .I(N__16937));
    LocalMux I__2785 (
            .O(N__16942),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__2784 (
            .O(N__16937),
            .I(M_this_data_count_qZ0Z_4));
    InMux I__2783 (
            .O(N__16932),
            .I(N__16929));
    LocalMux I__2782 (
            .O(N__16929),
            .I(N__16926));
    Odrv4 I__2781 (
            .O(N__16926),
            .I(M_this_data_count_q_cry_4_THRU_CO));
    CascadeMux I__2780 (
            .O(N__16923),
            .I(N__16920));
    InMux I__2779 (
            .O(N__16920),
            .I(N__16915));
    InMux I__2778 (
            .O(N__16919),
            .I(N__16910));
    InMux I__2777 (
            .O(N__16918),
            .I(N__16910));
    LocalMux I__2776 (
            .O(N__16915),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__2775 (
            .O(N__16910),
            .I(M_this_data_count_qZ0Z_5));
    InMux I__2774 (
            .O(N__16905),
            .I(N__16902));
    LocalMux I__2773 (
            .O(N__16902),
            .I(M_this_data_count_q_cry_6_THRU_CO));
    CascadeMux I__2772 (
            .O(N__16899),
            .I(N__16895));
    CascadeMux I__2771 (
            .O(N__16898),
            .I(N__16891));
    InMux I__2770 (
            .O(N__16895),
            .I(N__16888));
    InMux I__2769 (
            .O(N__16894),
            .I(N__16883));
    InMux I__2768 (
            .O(N__16891),
            .I(N__16883));
    LocalMux I__2767 (
            .O(N__16888),
            .I(M_this_data_count_qZ0Z_7));
    LocalMux I__2766 (
            .O(N__16883),
            .I(M_this_data_count_qZ0Z_7));
    InMux I__2765 (
            .O(N__16878),
            .I(N__16875));
    LocalMux I__2764 (
            .O(N__16875),
            .I(M_this_data_count_q_cry_2_THRU_CO));
    InMux I__2763 (
            .O(N__16872),
            .I(N__16869));
    LocalMux I__2762 (
            .O(N__16869),
            .I(M_this_data_count_q_cry_10_THRU_CO));
    InMux I__2761 (
            .O(N__16866),
            .I(N__16863));
    LocalMux I__2760 (
            .O(N__16863),
            .I(M_this_data_count_q_cry_11_THRU_CO));
    InMux I__2759 (
            .O(N__16860),
            .I(N__16855));
    InMux I__2758 (
            .O(N__16859),
            .I(N__16850));
    InMux I__2757 (
            .O(N__16858),
            .I(N__16850));
    LocalMux I__2756 (
            .O(N__16855),
            .I(M_this_data_count_qZ0Z_12));
    LocalMux I__2755 (
            .O(N__16850),
            .I(M_this_data_count_qZ0Z_12));
    CascadeMux I__2754 (
            .O(N__16845),
            .I(N__16841));
    InMux I__2753 (
            .O(N__16844),
            .I(N__16838));
    InMux I__2752 (
            .O(N__16841),
            .I(N__16835));
    LocalMux I__2751 (
            .O(N__16838),
            .I(N__16830));
    LocalMux I__2750 (
            .O(N__16835),
            .I(N__16830));
    Odrv4 I__2749 (
            .O(N__16830),
            .I(M_this_data_count_qZ0Z_13));
    InMux I__2748 (
            .O(N__16827),
            .I(N__16824));
    LocalMux I__2747 (
            .O(N__16824),
            .I(M_this_data_count_q_cry_7_THRU_CO));
    InMux I__2746 (
            .O(N__16821),
            .I(N__16816));
    InMux I__2745 (
            .O(N__16820),
            .I(N__16811));
    InMux I__2744 (
            .O(N__16819),
            .I(N__16811));
    LocalMux I__2743 (
            .O(N__16816),
            .I(M_this_data_count_qZ0Z_8));
    LocalMux I__2742 (
            .O(N__16811),
            .I(M_this_data_count_qZ0Z_8));
    InMux I__2741 (
            .O(N__16806),
            .I(N__16803));
    LocalMux I__2740 (
            .O(N__16803),
            .I(M_this_state_q_RNIOE1SZ0Z_11));
    InMux I__2739 (
            .O(N__16800),
            .I(N__16797));
    LocalMux I__2738 (
            .O(N__16797),
            .I(un20_i_a2_x_3));
    InMux I__2737 (
            .O(N__16794),
            .I(N__16791));
    LocalMux I__2736 (
            .O(N__16791),
            .I(M_this_state_q_RNIG01LZ0Z_12));
    CascadeMux I__2735 (
            .O(N__16788),
            .I(\this_vga_signals.N_419_i_i_0Z0Z_1_cascade_ ));
    InMux I__2734 (
            .O(N__16785),
            .I(N__16782));
    LocalMux I__2733 (
            .O(N__16782),
            .I(M_this_data_count_q_s_6));
    CascadeMux I__2732 (
            .O(N__16779),
            .I(N__16772));
    CascadeMux I__2731 (
            .O(N__16778),
            .I(N__16768));
    CascadeMux I__2730 (
            .O(N__16777),
            .I(N__16761));
    CascadeMux I__2729 (
            .O(N__16776),
            .I(N__16757));
    CascadeMux I__2728 (
            .O(N__16775),
            .I(N__16754));
    InMux I__2727 (
            .O(N__16772),
            .I(N__16744));
    InMux I__2726 (
            .O(N__16771),
            .I(N__16744));
    InMux I__2725 (
            .O(N__16768),
            .I(N__16744));
    InMux I__2724 (
            .O(N__16767),
            .I(N__16744));
    InMux I__2723 (
            .O(N__16766),
            .I(N__16737));
    InMux I__2722 (
            .O(N__16765),
            .I(N__16737));
    InMux I__2721 (
            .O(N__16764),
            .I(N__16731));
    InMux I__2720 (
            .O(N__16761),
            .I(N__16731));
    InMux I__2719 (
            .O(N__16760),
            .I(N__16728));
    InMux I__2718 (
            .O(N__16757),
            .I(N__16725));
    InMux I__2717 (
            .O(N__16754),
            .I(N__16722));
    InMux I__2716 (
            .O(N__16753),
            .I(N__16719));
    LocalMux I__2715 (
            .O(N__16744),
            .I(N__16716));
    InMux I__2714 (
            .O(N__16743),
            .I(N__16713));
    CascadeMux I__2713 (
            .O(N__16742),
            .I(N__16708));
    LocalMux I__2712 (
            .O(N__16737),
            .I(N__16704));
    CascadeMux I__2711 (
            .O(N__16736),
            .I(N__16700));
    LocalMux I__2710 (
            .O(N__16731),
            .I(N__16697));
    LocalMux I__2709 (
            .O(N__16728),
            .I(N__16692));
    LocalMux I__2708 (
            .O(N__16725),
            .I(N__16692));
    LocalMux I__2707 (
            .O(N__16722),
            .I(N__16687));
    LocalMux I__2706 (
            .O(N__16719),
            .I(N__16682));
    Span4Mux_v I__2705 (
            .O(N__16716),
            .I(N__16677));
    LocalMux I__2704 (
            .O(N__16713),
            .I(N__16677));
    InMux I__2703 (
            .O(N__16712),
            .I(N__16668));
    InMux I__2702 (
            .O(N__16711),
            .I(N__16668));
    InMux I__2701 (
            .O(N__16708),
            .I(N__16668));
    InMux I__2700 (
            .O(N__16707),
            .I(N__16668));
    Span4Mux_v I__2699 (
            .O(N__16704),
            .I(N__16665));
    InMux I__2698 (
            .O(N__16703),
            .I(N__16662));
    InMux I__2697 (
            .O(N__16700),
            .I(N__16659));
    Span4Mux_h I__2696 (
            .O(N__16697),
            .I(N__16656));
    Span4Mux_v I__2695 (
            .O(N__16692),
            .I(N__16653));
    InMux I__2694 (
            .O(N__16691),
            .I(N__16648));
    InMux I__2693 (
            .O(N__16690),
            .I(N__16648));
    Span4Mux_h I__2692 (
            .O(N__16687),
            .I(N__16645));
    InMux I__2691 (
            .O(N__16686),
            .I(N__16640));
    InMux I__2690 (
            .O(N__16685),
            .I(N__16640));
    Span4Mux_v I__2689 (
            .O(N__16682),
            .I(N__16635));
    Span4Mux_h I__2688 (
            .O(N__16677),
            .I(N__16635));
    LocalMux I__2687 (
            .O(N__16668),
            .I(N__16630));
    Span4Mux_h I__2686 (
            .O(N__16665),
            .I(N__16630));
    LocalMux I__2685 (
            .O(N__16662),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2684 (
            .O(N__16659),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2683 (
            .O(N__16656),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2682 (
            .O(N__16653),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2681 (
            .O(N__16648),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2680 (
            .O(N__16645),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2679 (
            .O(N__16640),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2678 (
            .O(N__16635),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2677 (
            .O(N__16630),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    InMux I__2676 (
            .O(N__16611),
            .I(N__16603));
    InMux I__2675 (
            .O(N__16610),
            .I(N__16603));
    InMux I__2674 (
            .O(N__16609),
            .I(N__16593));
    InMux I__2673 (
            .O(N__16608),
            .I(N__16590));
    LocalMux I__2672 (
            .O(N__16603),
            .I(N__16587));
    CascadeMux I__2671 (
            .O(N__16602),
            .I(N__16584));
    InMux I__2670 (
            .O(N__16601),
            .I(N__16578));
    InMux I__2669 (
            .O(N__16600),
            .I(N__16578));
    InMux I__2668 (
            .O(N__16599),
            .I(N__16571));
    InMux I__2667 (
            .O(N__16598),
            .I(N__16571));
    InMux I__2666 (
            .O(N__16597),
            .I(N__16571));
    InMux I__2665 (
            .O(N__16596),
            .I(N__16568));
    LocalMux I__2664 (
            .O(N__16593),
            .I(N__16565));
    LocalMux I__2663 (
            .O(N__16590),
            .I(N__16560));
    Span4Mux_h I__2662 (
            .O(N__16587),
            .I(N__16560));
    InMux I__2661 (
            .O(N__16584),
            .I(N__16557));
    InMux I__2660 (
            .O(N__16583),
            .I(N__16554));
    LocalMux I__2659 (
            .O(N__16578),
            .I(N__16551));
    LocalMux I__2658 (
            .O(N__16571),
            .I(N__16535));
    LocalMux I__2657 (
            .O(N__16568),
            .I(N__16535));
    Span4Mux_h I__2656 (
            .O(N__16565),
            .I(N__16535));
    Span4Mux_h I__2655 (
            .O(N__16560),
            .I(N__16535));
    LocalMux I__2654 (
            .O(N__16557),
            .I(N__16535));
    LocalMux I__2653 (
            .O(N__16554),
            .I(N__16535));
    Span4Mux_v I__2652 (
            .O(N__16551),
            .I(N__16531));
    InMux I__2651 (
            .O(N__16550),
            .I(N__16526));
    InMux I__2650 (
            .O(N__16549),
            .I(N__16526));
    InMux I__2649 (
            .O(N__16548),
            .I(N__16523));
    Span4Mux_v I__2648 (
            .O(N__16535),
            .I(N__16520));
    InMux I__2647 (
            .O(N__16534),
            .I(N__16517));
    Odrv4 I__2646 (
            .O(N__16531),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2645 (
            .O(N__16526),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2644 (
            .O(N__16523),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2643 (
            .O(N__16520),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2642 (
            .O(N__16517),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    CascadeMux I__2641 (
            .O(N__16506),
            .I(N__16503));
    InMux I__2640 (
            .O(N__16503),
            .I(N__16497));
    InMux I__2639 (
            .O(N__16502),
            .I(N__16497));
    LocalMux I__2638 (
            .O(N__16497),
            .I(\this_vga_signals.M_vcounter_d7lt8_0 ));
    CascadeMux I__2637 (
            .O(N__16494),
            .I(\this_vga_signals.M_vcounter_d7lto8_1_cascade_ ));
    InMux I__2636 (
            .O(N__16491),
            .I(N__16485));
    CascadeMux I__2635 (
            .O(N__16490),
            .I(N__16470));
    InMux I__2634 (
            .O(N__16489),
            .I(N__16466));
    InMux I__2633 (
            .O(N__16488),
            .I(N__16463));
    LocalMux I__2632 (
            .O(N__16485),
            .I(N__16460));
    CascadeMux I__2631 (
            .O(N__16484),
            .I(N__16452));
    InMux I__2630 (
            .O(N__16483),
            .I(N__16446));
    InMux I__2629 (
            .O(N__16482),
            .I(N__16446));
    CascadeMux I__2628 (
            .O(N__16481),
            .I(N__16443));
    CascadeMux I__2627 (
            .O(N__16480),
            .I(N__16440));
    InMux I__2626 (
            .O(N__16479),
            .I(N__16437));
    InMux I__2625 (
            .O(N__16478),
            .I(N__16434));
    InMux I__2624 (
            .O(N__16477),
            .I(N__16431));
    InMux I__2623 (
            .O(N__16476),
            .I(N__16428));
    InMux I__2622 (
            .O(N__16475),
            .I(N__16415));
    InMux I__2621 (
            .O(N__16474),
            .I(N__16415));
    InMux I__2620 (
            .O(N__16473),
            .I(N__16415));
    InMux I__2619 (
            .O(N__16470),
            .I(N__16415));
    InMux I__2618 (
            .O(N__16469),
            .I(N__16412));
    LocalMux I__2617 (
            .O(N__16466),
            .I(N__16405));
    LocalMux I__2616 (
            .O(N__16463),
            .I(N__16405));
    Span4Mux_h I__2615 (
            .O(N__16460),
            .I(N__16405));
    InMux I__2614 (
            .O(N__16459),
            .I(N__16400));
    InMux I__2613 (
            .O(N__16458),
            .I(N__16400));
    InMux I__2612 (
            .O(N__16457),
            .I(N__16395));
    InMux I__2611 (
            .O(N__16456),
            .I(N__16395));
    InMux I__2610 (
            .O(N__16455),
            .I(N__16389));
    InMux I__2609 (
            .O(N__16452),
            .I(N__16389));
    CascadeMux I__2608 (
            .O(N__16451),
            .I(N__16386));
    LocalMux I__2607 (
            .O(N__16446),
            .I(N__16382));
    InMux I__2606 (
            .O(N__16443),
            .I(N__16377));
    InMux I__2605 (
            .O(N__16440),
            .I(N__16377));
    LocalMux I__2604 (
            .O(N__16437),
            .I(N__16370));
    LocalMux I__2603 (
            .O(N__16434),
            .I(N__16370));
    LocalMux I__2602 (
            .O(N__16431),
            .I(N__16370));
    LocalMux I__2601 (
            .O(N__16428),
            .I(N__16367));
    InMux I__2600 (
            .O(N__16427),
            .I(N__16357));
    InMux I__2599 (
            .O(N__16426),
            .I(N__16357));
    InMux I__2598 (
            .O(N__16425),
            .I(N__16357));
    InMux I__2597 (
            .O(N__16424),
            .I(N__16357));
    LocalMux I__2596 (
            .O(N__16415),
            .I(N__16354));
    LocalMux I__2595 (
            .O(N__16412),
            .I(N__16347));
    Span4Mux_v I__2594 (
            .O(N__16405),
            .I(N__16347));
    LocalMux I__2593 (
            .O(N__16400),
            .I(N__16347));
    LocalMux I__2592 (
            .O(N__16395),
            .I(N__16344));
    InMux I__2591 (
            .O(N__16394),
            .I(N__16341));
    LocalMux I__2590 (
            .O(N__16389),
            .I(N__16338));
    InMux I__2589 (
            .O(N__16386),
            .I(N__16333));
    InMux I__2588 (
            .O(N__16385),
            .I(N__16333));
    Span4Mux_h I__2587 (
            .O(N__16382),
            .I(N__16324));
    LocalMux I__2586 (
            .O(N__16377),
            .I(N__16324));
    Span4Mux_v I__2585 (
            .O(N__16370),
            .I(N__16324));
    Span4Mux_h I__2584 (
            .O(N__16367),
            .I(N__16324));
    InMux I__2583 (
            .O(N__16366),
            .I(N__16321));
    LocalMux I__2582 (
            .O(N__16357),
            .I(N__16312));
    Span4Mux_h I__2581 (
            .O(N__16354),
            .I(N__16312));
    Span4Mux_h I__2580 (
            .O(N__16347),
            .I(N__16312));
    Span4Mux_v I__2579 (
            .O(N__16344),
            .I(N__16312));
    LocalMux I__2578 (
            .O(N__16341),
            .I(N__16307));
    Span4Mux_h I__2577 (
            .O(N__16338),
            .I(N__16307));
    LocalMux I__2576 (
            .O(N__16333),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2575 (
            .O(N__16324),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2574 (
            .O(N__16321),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2573 (
            .O(N__16312),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2572 (
            .O(N__16307),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    CascadeMux I__2571 (
            .O(N__16296),
            .I(\this_vga_signals.M_vcounter_d8_cascade_ ));
    IoInMux I__2570 (
            .O(N__16293),
            .I(N__16290));
    LocalMux I__2569 (
            .O(N__16290),
            .I(N__16287));
    Span12Mux_s7_h I__2568 (
            .O(N__16287),
            .I(N__16284));
    Odrv12 I__2567 (
            .O(N__16284),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ));
    InMux I__2566 (
            .O(N__16281),
            .I(N__16276));
    InMux I__2565 (
            .O(N__16280),
            .I(N__16271));
    InMux I__2564 (
            .O(N__16279),
            .I(N__16271));
    LocalMux I__2563 (
            .O(N__16276),
            .I(this_pixel_clk_M_counter_q_0));
    LocalMux I__2562 (
            .O(N__16271),
            .I(this_pixel_clk_M_counter_q_0));
    CascadeMux I__2561 (
            .O(N__16266),
            .I(N__16260));
    CascadeMux I__2560 (
            .O(N__16265),
            .I(N__16256));
    InMux I__2559 (
            .O(N__16264),
            .I(N__16252));
    InMux I__2558 (
            .O(N__16263),
            .I(N__16249));
    InMux I__2557 (
            .O(N__16260),
            .I(N__16240));
    InMux I__2556 (
            .O(N__16259),
            .I(N__16240));
    InMux I__2555 (
            .O(N__16256),
            .I(N__16240));
    InMux I__2554 (
            .O(N__16255),
            .I(N__16240));
    LocalMux I__2553 (
            .O(N__16252),
            .I(M_pcounter_q_ret_2_RNIH7PG8));
    LocalMux I__2552 (
            .O(N__16249),
            .I(M_pcounter_q_ret_2_RNIH7PG8));
    LocalMux I__2551 (
            .O(N__16240),
            .I(M_pcounter_q_ret_2_RNIH7PG8));
    InMux I__2550 (
            .O(N__16233),
            .I(N__16230));
    LocalMux I__2549 (
            .O(N__16230),
            .I(N__16226));
    CascadeMux I__2548 (
            .O(N__16229),
            .I(N__16223));
    Span4Mux_v I__2547 (
            .O(N__16226),
            .I(N__16220));
    InMux I__2546 (
            .O(N__16223),
            .I(N__16217));
    Odrv4 I__2545 (
            .O(N__16220),
            .I(\this_vga_ramdac.N_2865_reto ));
    LocalMux I__2544 (
            .O(N__16217),
            .I(\this_vga_ramdac.N_2865_reto ));
    CascadeMux I__2543 (
            .O(N__16212),
            .I(dma_ac0_5_0_cascade_));
    InMux I__2542 (
            .O(N__16209),
            .I(M_this_data_count_q_cry_8));
    CascadeMux I__2541 (
            .O(N__16206),
            .I(N__16203));
    InMux I__2540 (
            .O(N__16203),
            .I(N__16200));
    LocalMux I__2539 (
            .O(N__16200),
            .I(N__16197));
    Odrv4 I__2538 (
            .O(N__16197),
            .I(M_this_data_count_q_s_10));
    InMux I__2537 (
            .O(N__16194),
            .I(M_this_data_count_q_cry_9));
    InMux I__2536 (
            .O(N__16191),
            .I(M_this_data_count_q_cry_10));
    InMux I__2535 (
            .O(N__16188),
            .I(M_this_data_count_q_cry_11));
    InMux I__2534 (
            .O(N__16185),
            .I(M_this_data_count_q_cry_12));
    CascadeMux I__2533 (
            .O(N__16182),
            .I(N__16179));
    InMux I__2532 (
            .O(N__16179),
            .I(N__16176));
    LocalMux I__2531 (
            .O(N__16176),
            .I(N__16173));
    Odrv4 I__2530 (
            .O(N__16173),
            .I(M_this_data_count_q_s_13));
    InMux I__2529 (
            .O(N__16170),
            .I(N__16167));
    LocalMux I__2528 (
            .O(N__16167),
            .I(N__16164));
    Span12Mux_h I__2527 (
            .O(N__16164),
            .I(N__16161));
    Odrv12 I__2526 (
            .O(N__16161),
            .I(N_87_0));
    InMux I__2525 (
            .O(N__16158),
            .I(N__16155));
    LocalMux I__2524 (
            .O(N__16155),
            .I(N__16152));
    Odrv12 I__2523 (
            .O(N__16152),
            .I(N_81_0));
    InMux I__2522 (
            .O(N__16149),
            .I(M_this_data_count_q_cry_0));
    InMux I__2521 (
            .O(N__16146),
            .I(M_this_data_count_q_cry_1));
    InMux I__2520 (
            .O(N__16143),
            .I(M_this_data_count_q_cry_2));
    InMux I__2519 (
            .O(N__16140),
            .I(M_this_data_count_q_cry_3));
    InMux I__2518 (
            .O(N__16137),
            .I(M_this_data_count_q_cry_4));
    InMux I__2517 (
            .O(N__16134),
            .I(M_this_data_count_q_cry_5));
    InMux I__2516 (
            .O(N__16131),
            .I(M_this_data_count_q_cry_6));
    InMux I__2515 (
            .O(N__16128),
            .I(bfn_14_26_0_));
    InMux I__2514 (
            .O(N__16125),
            .I(N__16122));
    LocalMux I__2513 (
            .O(N__16122),
            .I(N__16119));
    Span4Mux_h I__2512 (
            .O(N__16119),
            .I(N__16116));
    Span4Mux_h I__2511 (
            .O(N__16116),
            .I(N__16113));
    Odrv4 I__2510 (
            .O(N__16113),
            .I(\this_vga_ramdac.i2_mux ));
    InMux I__2509 (
            .O(N__16110),
            .I(N__16106));
    InMux I__2508 (
            .O(N__16109),
            .I(N__16103));
    LocalMux I__2507 (
            .O(N__16106),
            .I(\this_vga_ramdac.N_2864_reto ));
    LocalMux I__2506 (
            .O(N__16103),
            .I(\this_vga_ramdac.N_2864_reto ));
    IoInMux I__2505 (
            .O(N__16098),
            .I(N__16091));
    IoInMux I__2504 (
            .O(N__16097),
            .I(N__16088));
    IoInMux I__2503 (
            .O(N__16096),
            .I(N__16085));
    IoInMux I__2502 (
            .O(N__16095),
            .I(N__16080));
    IoInMux I__2501 (
            .O(N__16094),
            .I(N__16077));
    LocalMux I__2500 (
            .O(N__16091),
            .I(N__16072));
    LocalMux I__2499 (
            .O(N__16088),
            .I(N__16072));
    LocalMux I__2498 (
            .O(N__16085),
            .I(N__16069));
    IoInMux I__2497 (
            .O(N__16084),
            .I(N__16066));
    IoInMux I__2496 (
            .O(N__16083),
            .I(N__16063));
    LocalMux I__2495 (
            .O(N__16080),
            .I(N__16058));
    LocalMux I__2494 (
            .O(N__16077),
            .I(N__16053));
    IoSpan4Mux I__2493 (
            .O(N__16072),
            .I(N__16050));
    IoSpan4Mux I__2492 (
            .O(N__16069),
            .I(N__16043));
    LocalMux I__2491 (
            .O(N__16066),
            .I(N__16043));
    LocalMux I__2490 (
            .O(N__16063),
            .I(N__16043));
    IoInMux I__2489 (
            .O(N__16062),
            .I(N__16040));
    IoInMux I__2488 (
            .O(N__16061),
            .I(N__16037));
    IoSpan4Mux I__2487 (
            .O(N__16058),
            .I(N__16034));
    IoInMux I__2486 (
            .O(N__16057),
            .I(N__16031));
    IoInMux I__2485 (
            .O(N__16056),
            .I(N__16028));
    IoSpan4Mux I__2484 (
            .O(N__16053),
            .I(N__16023));
    Span4Mux_s1_h I__2483 (
            .O(N__16050),
            .I(N__16019));
    IoSpan4Mux I__2482 (
            .O(N__16043),
            .I(N__16012));
    LocalMux I__2481 (
            .O(N__16040),
            .I(N__16012));
    LocalMux I__2480 (
            .O(N__16037),
            .I(N__16012));
    IoSpan4Mux I__2479 (
            .O(N__16034),
            .I(N__16007));
    LocalMux I__2478 (
            .O(N__16031),
            .I(N__16007));
    LocalMux I__2477 (
            .O(N__16028),
            .I(N__16004));
    IoInMux I__2476 (
            .O(N__16027),
            .I(N__16001));
    IoInMux I__2475 (
            .O(N__16026),
            .I(N__15996));
    Span4Mux_s3_h I__2474 (
            .O(N__16023),
            .I(N__15993));
    IoInMux I__2473 (
            .O(N__16022),
            .I(N__15990));
    Span4Mux_h I__2472 (
            .O(N__16019),
            .I(N__15984));
    IoSpan4Mux I__2471 (
            .O(N__16012),
            .I(N__15984));
    IoSpan4Mux I__2470 (
            .O(N__16007),
            .I(N__15977));
    IoSpan4Mux I__2469 (
            .O(N__16004),
            .I(N__15977));
    LocalMux I__2468 (
            .O(N__16001),
            .I(N__15977));
    IoInMux I__2467 (
            .O(N__16000),
            .I(N__15974));
    IoInMux I__2466 (
            .O(N__15999),
            .I(N__15971));
    LocalMux I__2465 (
            .O(N__15996),
            .I(N__15968));
    Span4Mux_h I__2464 (
            .O(N__15993),
            .I(N__15965));
    LocalMux I__2463 (
            .O(N__15990),
            .I(N__15962));
    IoInMux I__2462 (
            .O(N__15989),
            .I(N__15959));
    Span4Mux_s1_h I__2461 (
            .O(N__15984),
            .I(N__15956));
    IoSpan4Mux I__2460 (
            .O(N__15977),
            .I(N__15949));
    LocalMux I__2459 (
            .O(N__15974),
            .I(N__15949));
    LocalMux I__2458 (
            .O(N__15971),
            .I(N__15949));
    IoSpan4Mux I__2457 (
            .O(N__15968),
            .I(N__15946));
    Sp12to4 I__2456 (
            .O(N__15965),
            .I(N__15941));
    Span12Mux_s6_h I__2455 (
            .O(N__15962),
            .I(N__15941));
    LocalMux I__2454 (
            .O(N__15959),
            .I(N__15938));
    Sp12to4 I__2453 (
            .O(N__15956),
            .I(N__15935));
    IoSpan4Mux I__2452 (
            .O(N__15949),
            .I(N__15932));
    Span4Mux_s2_h I__2451 (
            .O(N__15946),
            .I(N__15929));
    Span12Mux_h I__2450 (
            .O(N__15941),
            .I(N__15926));
    Span12Mux_s2_v I__2449 (
            .O(N__15938),
            .I(N__15923));
    Span12Mux_s6_h I__2448 (
            .O(N__15935),
            .I(N__15920));
    Span4Mux_s2_v I__2447 (
            .O(N__15932),
            .I(N__15917));
    Span4Mux_h I__2446 (
            .O(N__15929),
            .I(N__15914));
    Span12Mux_v I__2445 (
            .O(N__15926),
            .I(N__15905));
    Span12Mux_h I__2444 (
            .O(N__15923),
            .I(N__15905));
    Span12Mux_h I__2443 (
            .O(N__15920),
            .I(N__15905));
    Sp12to4 I__2442 (
            .O(N__15917),
            .I(N__15905));
    Span4Mux_h I__2441 (
            .O(N__15914),
            .I(N__15902));
    Odrv12 I__2440 (
            .O(N__15905),
            .I(dma_0_i));
    Odrv4 I__2439 (
            .O(N__15902),
            .I(dma_0_i));
    InMux I__2438 (
            .O(N__15897),
            .I(N__15892));
    InMux I__2437 (
            .O(N__15896),
            .I(N__15887));
    InMux I__2436 (
            .O(N__15895),
            .I(N__15887));
    LocalMux I__2435 (
            .O(N__15892),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    LocalMux I__2434 (
            .O(N__15887),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    InMux I__2433 (
            .O(N__15882),
            .I(N__15879));
    LocalMux I__2432 (
            .O(N__15879),
            .I(\this_vga_signals.M_pcounter_q_3_0 ));
    CascadeMux I__2431 (
            .O(N__15876),
            .I(N__15871));
    CascadeMux I__2430 (
            .O(N__15875),
            .I(N__15868));
    InMux I__2429 (
            .O(N__15874),
            .I(N__15865));
    InMux I__2428 (
            .O(N__15871),
            .I(N__15860));
    InMux I__2427 (
            .O(N__15868),
            .I(N__15860));
    LocalMux I__2426 (
            .O(N__15865),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    LocalMux I__2425 (
            .O(N__15860),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    InMux I__2424 (
            .O(N__15855),
            .I(N__15852));
    LocalMux I__2423 (
            .O(N__15852),
            .I(\this_vga_signals.M_pcounter_q_3_1 ));
    CascadeMux I__2422 (
            .O(N__15849),
            .I(N__15846));
    InMux I__2421 (
            .O(N__15846),
            .I(N__15840));
    InMux I__2420 (
            .O(N__15845),
            .I(N__15840));
    LocalMux I__2419 (
            .O(N__15840),
            .I(\this_vga_signals.N_3_0 ));
    CascadeMux I__2418 (
            .O(N__15837),
            .I(\this_vga_signals.N_3_0_cascade_ ));
    InMux I__2417 (
            .O(N__15834),
            .I(N__15822));
    InMux I__2416 (
            .O(N__15833),
            .I(N__15822));
    InMux I__2415 (
            .O(N__15832),
            .I(N__15822));
    InMux I__2414 (
            .O(N__15831),
            .I(N__15822));
    LocalMux I__2413 (
            .O(N__15822),
            .I(\this_vga_signals.M_pcounter_q_i_3_1 ));
    InMux I__2412 (
            .O(N__15819),
            .I(N__15812));
    InMux I__2411 (
            .O(N__15818),
            .I(N__15812));
    InMux I__2410 (
            .O(N__15817),
            .I(N__15809));
    LocalMux I__2409 (
            .O(N__15812),
            .I(N__15806));
    LocalMux I__2408 (
            .O(N__15809),
            .I(N__15801));
    Span4Mux_h I__2407 (
            .O(N__15806),
            .I(N__15798));
    InMux I__2406 (
            .O(N__15805),
            .I(N__15795));
    InMux I__2405 (
            .O(N__15804),
            .I(N__15792));
    Span4Mux_v I__2404 (
            .O(N__15801),
            .I(N__15787));
    Span4Mux_h I__2403 (
            .O(N__15798),
            .I(N__15780));
    LocalMux I__2402 (
            .O(N__15795),
            .I(N__15780));
    LocalMux I__2401 (
            .O(N__15792),
            .I(N__15780));
    InMux I__2400 (
            .O(N__15791),
            .I(N__15777));
    InMux I__2399 (
            .O(N__15790),
            .I(N__15774));
    Odrv4 I__2398 (
            .O(N__15787),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    Odrv4 I__2397 (
            .O(N__15780),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    LocalMux I__2396 (
            .O(N__15777),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    LocalMux I__2395 (
            .O(N__15774),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ));
    InMux I__2394 (
            .O(N__15765),
            .I(N__15762));
    LocalMux I__2393 (
            .O(N__15762),
            .I(N__15758));
    InMux I__2392 (
            .O(N__15761),
            .I(N__15755));
    Odrv12 I__2391 (
            .O(N__15758),
            .I(\this_vga_ramdac.N_2867_reto ));
    LocalMux I__2390 (
            .O(N__15755),
            .I(\this_vga_ramdac.N_2867_reto ));
    IoInMux I__2389 (
            .O(N__15750),
            .I(N__15747));
    LocalMux I__2388 (
            .O(N__15747),
            .I(N__15744));
    Span4Mux_s3_h I__2387 (
            .O(N__15744),
            .I(N__15741));
    Span4Mux_h I__2386 (
            .O(N__15741),
            .I(N__15738));
    Sp12to4 I__2385 (
            .O(N__15738),
            .I(N__15735));
    Span12Mux_s11_v I__2384 (
            .O(N__15735),
            .I(N__15732));
    Odrv12 I__2383 (
            .O(N__15732),
            .I(rgb_c_5));
    InMux I__2382 (
            .O(N__15729),
            .I(N__15724));
    InMux I__2381 (
            .O(N__15728),
            .I(N__15719));
    InMux I__2380 (
            .O(N__15727),
            .I(N__15719));
    LocalMux I__2379 (
            .O(N__15724),
            .I(\this_vga_signals.N_2_0 ));
    LocalMux I__2378 (
            .O(N__15719),
            .I(\this_vga_signals.N_2_0 ));
    InMux I__2377 (
            .O(N__15714),
            .I(N__15710));
    InMux I__2376 (
            .O(N__15713),
            .I(N__15707));
    LocalMux I__2375 (
            .O(N__15710),
            .I(\this_vga_signals.M_pcounter_q_i_3_0 ));
    LocalMux I__2374 (
            .O(N__15707),
            .I(\this_vga_signals.M_pcounter_q_i_3_0 ));
    InMux I__2373 (
            .O(N__15702),
            .I(N__15696));
    InMux I__2372 (
            .O(N__15701),
            .I(N__15696));
    LocalMux I__2371 (
            .O(N__15696),
            .I(this_pixel_clk_M_counter_q_i_1));
    IoInMux I__2370 (
            .O(N__15693),
            .I(N__15690));
    LocalMux I__2369 (
            .O(N__15690),
            .I(N__15687));
    Span4Mux_s1_h I__2368 (
            .O(N__15687),
            .I(N__15684));
    Span4Mux_h I__2367 (
            .O(N__15684),
            .I(N__15681));
    Span4Mux_h I__2366 (
            .O(N__15681),
            .I(N__15678));
    Span4Mux_h I__2365 (
            .O(N__15678),
            .I(N__15675));
    Odrv4 I__2364 (
            .O(N__15675),
            .I(rgb_c_2));
    InMux I__2363 (
            .O(N__15672),
            .I(N__15669));
    LocalMux I__2362 (
            .O(N__15669),
            .I(N__15666));
    Odrv4 I__2361 (
            .O(N__15666),
            .I(\this_vga_ramdac.m6 ));
    InMux I__2360 (
            .O(N__15663),
            .I(N__15660));
    LocalMux I__2359 (
            .O(N__15660),
            .I(N__15657));
    Span4Mux_v I__2358 (
            .O(N__15657),
            .I(N__15654));
    Span4Mux_h I__2357 (
            .O(N__15654),
            .I(N__15650));
    CascadeMux I__2356 (
            .O(N__15653),
            .I(N__15647));
    Span4Mux_h I__2355 (
            .O(N__15650),
            .I(N__15644));
    InMux I__2354 (
            .O(N__15647),
            .I(N__15641));
    Odrv4 I__2353 (
            .O(N__15644),
            .I(\this_vga_ramdac.N_2863_reto ));
    LocalMux I__2352 (
            .O(N__15641),
            .I(\this_vga_ramdac.N_2863_reto ));
    InMux I__2351 (
            .O(N__15636),
            .I(N__15633));
    LocalMux I__2350 (
            .O(N__15633),
            .I(N__15630));
    Odrv4 I__2349 (
            .O(N__15630),
            .I(\this_vga_ramdac.i2_mux_0 ));
    InMux I__2348 (
            .O(N__15627),
            .I(N__15624));
    LocalMux I__2347 (
            .O(N__15624),
            .I(N__15621));
    Odrv4 I__2346 (
            .O(N__15621),
            .I(\this_vga_ramdac.m19 ));
    InMux I__2345 (
            .O(N__15618),
            .I(N__15615));
    LocalMux I__2344 (
            .O(N__15615),
            .I(N__15611));
    CascadeMux I__2343 (
            .O(N__15614),
            .I(N__15608));
    Span4Mux_h I__2342 (
            .O(N__15611),
            .I(N__15605));
    InMux I__2341 (
            .O(N__15608),
            .I(N__15602));
    Odrv4 I__2340 (
            .O(N__15605),
            .I(\this_vga_ramdac.N_2866_reto ));
    LocalMux I__2339 (
            .O(N__15602),
            .I(\this_vga_ramdac.N_2866_reto ));
    InMux I__2338 (
            .O(N__15597),
            .I(N__15594));
    LocalMux I__2337 (
            .O(N__15594),
            .I(\this_vga_signals.M_this_vga_signals_pixel_clk_0_0 ));
    InMux I__2336 (
            .O(N__15591),
            .I(N__15584));
    InMux I__2335 (
            .O(N__15590),
            .I(N__15581));
    InMux I__2334 (
            .O(N__15589),
            .I(N__15578));
    InMux I__2333 (
            .O(N__15588),
            .I(N__15573));
    InMux I__2332 (
            .O(N__15587),
            .I(N__15573));
    LocalMux I__2331 (
            .O(N__15584),
            .I(N__15570));
    LocalMux I__2330 (
            .O(N__15581),
            .I(N__15567));
    LocalMux I__2329 (
            .O(N__15578),
            .I(N__15562));
    LocalMux I__2328 (
            .O(N__15573),
            .I(N__15562));
    Span4Mux_h I__2327 (
            .O(N__15570),
            .I(N__15555));
    Span4Mux_h I__2326 (
            .O(N__15567),
            .I(N__15552));
    Span4Mux_h I__2325 (
            .O(N__15562),
            .I(N__15549));
    InMux I__2324 (
            .O(N__15561),
            .I(N__15546));
    InMux I__2323 (
            .O(N__15560),
            .I(N__15541));
    InMux I__2322 (
            .O(N__15559),
            .I(N__15541));
    InMux I__2321 (
            .O(N__15558),
            .I(N__15538));
    Odrv4 I__2320 (
            .O(N__15555),
            .I(M_this_vga_ramdac_en_0));
    Odrv4 I__2319 (
            .O(N__15552),
            .I(M_this_vga_ramdac_en_0));
    Odrv4 I__2318 (
            .O(N__15549),
            .I(M_this_vga_ramdac_en_0));
    LocalMux I__2317 (
            .O(N__15546),
            .I(M_this_vga_ramdac_en_0));
    LocalMux I__2316 (
            .O(N__15541),
            .I(M_this_vga_ramdac_en_0));
    LocalMux I__2315 (
            .O(N__15538),
            .I(M_this_vga_ramdac_en_0));
    CascadeMux I__2314 (
            .O(N__15525),
            .I(M_pcounter_q_ret_2_RNIH7PG8_cascade_));
    IoInMux I__2313 (
            .O(N__15522),
            .I(N__15519));
    LocalMux I__2312 (
            .O(N__15519),
            .I(N__15516));
    IoSpan4Mux I__2311 (
            .O(N__15516),
            .I(N__15513));
    Span4Mux_s2_h I__2310 (
            .O(N__15513),
            .I(N__15510));
    Span4Mux_h I__2309 (
            .O(N__15510),
            .I(N__15507));
    Span4Mux_h I__2308 (
            .O(N__15507),
            .I(N__15504));
    Odrv4 I__2307 (
            .O(N__15504),
            .I(rgb_c_3));
    InMux I__2306 (
            .O(N__15501),
            .I(N__15498));
    LocalMux I__2305 (
            .O(N__15498),
            .I(N__15495));
    Span4Mux_v I__2304 (
            .O(N__15495),
            .I(N__15492));
    Span4Mux_h I__2303 (
            .O(N__15492),
            .I(N__15489));
    Odrv4 I__2302 (
            .O(N__15489),
            .I(N_95_0));
    CascadeMux I__2301 (
            .O(N__15486),
            .I(N__15482));
    InMux I__2300 (
            .O(N__15485),
            .I(N__15478));
    InMux I__2299 (
            .O(N__15482),
            .I(N__15475));
    InMux I__2298 (
            .O(N__15481),
            .I(N__15472));
    LocalMux I__2297 (
            .O(N__15478),
            .I(N__15469));
    LocalMux I__2296 (
            .O(N__15475),
            .I(N__15464));
    LocalMux I__2295 (
            .O(N__15472),
            .I(N__15464));
    Span4Mux_v I__2294 (
            .O(N__15469),
            .I(N__15458));
    Span4Mux_v I__2293 (
            .O(N__15464),
            .I(N__15458));
    InMux I__2292 (
            .O(N__15463),
            .I(N__15452));
    Span4Mux_h I__2291 (
            .O(N__15458),
            .I(N__15449));
    InMux I__2290 (
            .O(N__15457),
            .I(N__15446));
    InMux I__2289 (
            .O(N__15456),
            .I(N__15443));
    InMux I__2288 (
            .O(N__15455),
            .I(N__15440));
    LocalMux I__2287 (
            .O(N__15452),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__2286 (
            .O(N__15449),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2285 (
            .O(N__15446),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2284 (
            .O(N__15443),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2283 (
            .O(N__15440),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    InMux I__2282 (
            .O(N__15429),
            .I(N__15426));
    LocalMux I__2281 (
            .O(N__15426),
            .I(N__15422));
    InMux I__2280 (
            .O(N__15425),
            .I(N__15418));
    Span4Mux_h I__2279 (
            .O(N__15422),
            .I(N__15415));
    InMux I__2278 (
            .O(N__15421),
            .I(N__15412));
    LocalMux I__2277 (
            .O(N__15418),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv4 I__2276 (
            .O(N__15415),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__2275 (
            .O(N__15412),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    InMux I__2274 (
            .O(N__15405),
            .I(N__15400));
    InMux I__2273 (
            .O(N__15404),
            .I(N__15397));
    CascadeMux I__2272 (
            .O(N__15403),
            .I(N__15388));
    LocalMux I__2271 (
            .O(N__15400),
            .I(N__15382));
    LocalMux I__2270 (
            .O(N__15397),
            .I(N__15382));
    InMux I__2269 (
            .O(N__15396),
            .I(N__15379));
    InMux I__2268 (
            .O(N__15395),
            .I(N__15374));
    InMux I__2267 (
            .O(N__15394),
            .I(N__15374));
    InMux I__2266 (
            .O(N__15393),
            .I(N__15371));
    InMux I__2265 (
            .O(N__15392),
            .I(N__15366));
    InMux I__2264 (
            .O(N__15391),
            .I(N__15366));
    InMux I__2263 (
            .O(N__15388),
            .I(N__15362));
    InMux I__2262 (
            .O(N__15387),
            .I(N__15357));
    Span4Mux_v I__2261 (
            .O(N__15382),
            .I(N__15352));
    LocalMux I__2260 (
            .O(N__15379),
            .I(N__15352));
    LocalMux I__2259 (
            .O(N__15374),
            .I(N__15347));
    LocalMux I__2258 (
            .O(N__15371),
            .I(N__15347));
    LocalMux I__2257 (
            .O(N__15366),
            .I(N__15344));
    CascadeMux I__2256 (
            .O(N__15365),
            .I(N__15341));
    LocalMux I__2255 (
            .O(N__15362),
            .I(N__15338));
    InMux I__2254 (
            .O(N__15361),
            .I(N__15335));
    InMux I__2253 (
            .O(N__15360),
            .I(N__15332));
    LocalMux I__2252 (
            .O(N__15357),
            .I(N__15325));
    Span4Mux_h I__2251 (
            .O(N__15352),
            .I(N__15325));
    Span4Mux_h I__2250 (
            .O(N__15347),
            .I(N__15325));
    Span12Mux_h I__2249 (
            .O(N__15344),
            .I(N__15322));
    InMux I__2248 (
            .O(N__15341),
            .I(N__15319));
    Odrv12 I__2247 (
            .O(N__15338),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__2246 (
            .O(N__15335),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__2245 (
            .O(N__15332),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2244 (
            .O(N__15325),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv12 I__2243 (
            .O(N__15322),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__2242 (
            .O(N__15319),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    CascadeMux I__2241 (
            .O(N__15306),
            .I(N__15303));
    InMux I__2240 (
            .O(N__15303),
            .I(N__15299));
    CascadeMux I__2239 (
            .O(N__15302),
            .I(N__15292));
    LocalMux I__2238 (
            .O(N__15299),
            .I(N__15288));
    InMux I__2237 (
            .O(N__15298),
            .I(N__15283));
    InMux I__2236 (
            .O(N__15297),
            .I(N__15283));
    InMux I__2235 (
            .O(N__15296),
            .I(N__15279));
    InMux I__2234 (
            .O(N__15295),
            .I(N__15276));
    InMux I__2233 (
            .O(N__15292),
            .I(N__15268));
    CascadeMux I__2232 (
            .O(N__15291),
            .I(N__15264));
    Span4Mux_v I__2231 (
            .O(N__15288),
            .I(N__15258));
    LocalMux I__2230 (
            .O(N__15283),
            .I(N__15258));
    InMux I__2229 (
            .O(N__15282),
            .I(N__15255));
    LocalMux I__2228 (
            .O(N__15279),
            .I(N__15250));
    LocalMux I__2227 (
            .O(N__15276),
            .I(N__15250));
    InMux I__2226 (
            .O(N__15275),
            .I(N__15247));
    InMux I__2225 (
            .O(N__15274),
            .I(N__15242));
    InMux I__2224 (
            .O(N__15273),
            .I(N__15242));
    CascadeMux I__2223 (
            .O(N__15272),
            .I(N__15237));
    CascadeMux I__2222 (
            .O(N__15271),
            .I(N__15231));
    LocalMux I__2221 (
            .O(N__15268),
            .I(N__15227));
    InMux I__2220 (
            .O(N__15267),
            .I(N__15222));
    InMux I__2219 (
            .O(N__15264),
            .I(N__15217));
    InMux I__2218 (
            .O(N__15263),
            .I(N__15217));
    Span4Mux_h I__2217 (
            .O(N__15258),
            .I(N__15214));
    LocalMux I__2216 (
            .O(N__15255),
            .I(N__15205));
    Span4Mux_v I__2215 (
            .O(N__15250),
            .I(N__15205));
    LocalMux I__2214 (
            .O(N__15247),
            .I(N__15205));
    LocalMux I__2213 (
            .O(N__15242),
            .I(N__15205));
    InMux I__2212 (
            .O(N__15241),
            .I(N__15198));
    InMux I__2211 (
            .O(N__15240),
            .I(N__15198));
    InMux I__2210 (
            .O(N__15237),
            .I(N__15198));
    InMux I__2209 (
            .O(N__15236),
            .I(N__15194));
    InMux I__2208 (
            .O(N__15235),
            .I(N__15185));
    InMux I__2207 (
            .O(N__15234),
            .I(N__15185));
    InMux I__2206 (
            .O(N__15231),
            .I(N__15185));
    InMux I__2205 (
            .O(N__15230),
            .I(N__15185));
    Span4Mux_v I__2204 (
            .O(N__15227),
            .I(N__15182));
    InMux I__2203 (
            .O(N__15226),
            .I(N__15177));
    InMux I__2202 (
            .O(N__15225),
            .I(N__15177));
    LocalMux I__2201 (
            .O(N__15222),
            .I(N__15166));
    LocalMux I__2200 (
            .O(N__15217),
            .I(N__15166));
    Span4Mux_h I__2199 (
            .O(N__15214),
            .I(N__15166));
    Span4Mux_h I__2198 (
            .O(N__15205),
            .I(N__15166));
    LocalMux I__2197 (
            .O(N__15198),
            .I(N__15166));
    InMux I__2196 (
            .O(N__15197),
            .I(N__15163));
    LocalMux I__2195 (
            .O(N__15194),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2194 (
            .O(N__15185),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2193 (
            .O(N__15182),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2192 (
            .O(N__15177),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2191 (
            .O(N__15166),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2190 (
            .O(N__15163),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    InMux I__2189 (
            .O(N__15150),
            .I(N__15147));
    LocalMux I__2188 (
            .O(N__15147),
            .I(N__15144));
    Span4Mux_h I__2187 (
            .O(N__15144),
            .I(N__15141));
    Span4Mux_v I__2186 (
            .O(N__15141),
            .I(N__15138));
    Span4Mux_v I__2185 (
            .O(N__15138),
            .I(N__15135));
    Odrv4 I__2184 (
            .O(N__15135),
            .I(M_this_map_ram_read_data_2));
    CascadeMux I__2183 (
            .O(N__15132),
            .I(N__15129));
    InMux I__2182 (
            .O(N__15129),
            .I(N__15122));
    CascadeMux I__2181 (
            .O(N__15128),
            .I(N__15119));
    CascadeMux I__2180 (
            .O(N__15127),
            .I(N__15114));
    CascadeMux I__2179 (
            .O(N__15126),
            .I(N__15111));
    CascadeMux I__2178 (
            .O(N__15125),
            .I(N__15108));
    LocalMux I__2177 (
            .O(N__15122),
            .I(N__15103));
    InMux I__2176 (
            .O(N__15119),
            .I(N__15100));
    CascadeMux I__2175 (
            .O(N__15118),
            .I(N__15097));
    CascadeMux I__2174 (
            .O(N__15117),
            .I(N__15094));
    InMux I__2173 (
            .O(N__15114),
            .I(N__15089));
    InMux I__2172 (
            .O(N__15111),
            .I(N__15085));
    InMux I__2171 (
            .O(N__15108),
            .I(N__15082));
    CascadeMux I__2170 (
            .O(N__15107),
            .I(N__15079));
    CascadeMux I__2169 (
            .O(N__15106),
            .I(N__15076));
    Span4Mux_h I__2168 (
            .O(N__15103),
            .I(N__15070));
    LocalMux I__2167 (
            .O(N__15100),
            .I(N__15070));
    InMux I__2166 (
            .O(N__15097),
            .I(N__15067));
    InMux I__2165 (
            .O(N__15094),
            .I(N__15064));
    CascadeMux I__2164 (
            .O(N__15093),
            .I(N__15061));
    CascadeMux I__2163 (
            .O(N__15092),
            .I(N__15058));
    LocalMux I__2162 (
            .O(N__15089),
            .I(N__15053));
    CascadeMux I__2161 (
            .O(N__15088),
            .I(N__15050));
    LocalMux I__2160 (
            .O(N__15085),
            .I(N__15045));
    LocalMux I__2159 (
            .O(N__15082),
            .I(N__15045));
    InMux I__2158 (
            .O(N__15079),
            .I(N__15042));
    InMux I__2157 (
            .O(N__15076),
            .I(N__15039));
    CascadeMux I__2156 (
            .O(N__15075),
            .I(N__15035));
    Span4Mux_v I__2155 (
            .O(N__15070),
            .I(N__15030));
    LocalMux I__2154 (
            .O(N__15067),
            .I(N__15030));
    LocalMux I__2153 (
            .O(N__15064),
            .I(N__15027));
    InMux I__2152 (
            .O(N__15061),
            .I(N__15024));
    InMux I__2151 (
            .O(N__15058),
            .I(N__15021));
    CascadeMux I__2150 (
            .O(N__15057),
            .I(N__15018));
    CascadeMux I__2149 (
            .O(N__15056),
            .I(N__15015));
    Span4Mux_v I__2148 (
            .O(N__15053),
            .I(N__15012));
    InMux I__2147 (
            .O(N__15050),
            .I(N__15009));
    Span4Mux_v I__2146 (
            .O(N__15045),
            .I(N__15002));
    LocalMux I__2145 (
            .O(N__15042),
            .I(N__15002));
    LocalMux I__2144 (
            .O(N__15039),
            .I(N__15002));
    CascadeMux I__2143 (
            .O(N__15038),
            .I(N__14999));
    InMux I__2142 (
            .O(N__15035),
            .I(N__14996));
    Span4Mux_h I__2141 (
            .O(N__15030),
            .I(N__14993));
    Span4Mux_v I__2140 (
            .O(N__15027),
            .I(N__14988));
    LocalMux I__2139 (
            .O(N__15024),
            .I(N__14988));
    LocalMux I__2138 (
            .O(N__15021),
            .I(N__14985));
    InMux I__2137 (
            .O(N__15018),
            .I(N__14982));
    InMux I__2136 (
            .O(N__15015),
            .I(N__14979));
    Sp12to4 I__2135 (
            .O(N__15012),
            .I(N__14974));
    LocalMux I__2134 (
            .O(N__15009),
            .I(N__14974));
    Span4Mux_v I__2133 (
            .O(N__15002),
            .I(N__14971));
    InMux I__2132 (
            .O(N__14999),
            .I(N__14968));
    LocalMux I__2131 (
            .O(N__14996),
            .I(N__14965));
    Span4Mux_v I__2130 (
            .O(N__14993),
            .I(N__14960));
    Span4Mux_h I__2129 (
            .O(N__14988),
            .I(N__14960));
    Span4Mux_h I__2128 (
            .O(N__14985),
            .I(N__14957));
    LocalMux I__2127 (
            .O(N__14982),
            .I(N__14954));
    LocalMux I__2126 (
            .O(N__14979),
            .I(N__14951));
    Span12Mux_h I__2125 (
            .O(N__14974),
            .I(N__14948));
    Sp12to4 I__2124 (
            .O(N__14971),
            .I(N__14943));
    LocalMux I__2123 (
            .O(N__14968),
            .I(N__14943));
    Span4Mux_h I__2122 (
            .O(N__14965),
            .I(N__14940));
    Span4Mux_h I__2121 (
            .O(N__14960),
            .I(N__14937));
    Span4Mux_v I__2120 (
            .O(N__14957),
            .I(N__14932));
    Span4Mux_h I__2119 (
            .O(N__14954),
            .I(N__14932));
    Span4Mux_h I__2118 (
            .O(N__14951),
            .I(N__14929));
    Span12Mux_v I__2117 (
            .O(N__14948),
            .I(N__14926));
    Span12Mux_h I__2116 (
            .O(N__14943),
            .I(N__14923));
    Span4Mux_v I__2115 (
            .O(N__14940),
            .I(N__14920));
    Span4Mux_h I__2114 (
            .O(N__14937),
            .I(N__14913));
    Span4Mux_h I__2113 (
            .O(N__14932),
            .I(N__14913));
    Span4Mux_h I__2112 (
            .O(N__14929),
            .I(N__14913));
    Odrv12 I__2111 (
            .O(N__14926),
            .I(M_this_ppu_sprites_addr_8));
    Odrv12 I__2110 (
            .O(N__14923),
            .I(M_this_ppu_sprites_addr_8));
    Odrv4 I__2109 (
            .O(N__14920),
            .I(M_this_ppu_sprites_addr_8));
    Odrv4 I__2108 (
            .O(N__14913),
            .I(M_this_ppu_sprites_addr_8));
    InMux I__2107 (
            .O(N__14904),
            .I(N__14901));
    LocalMux I__2106 (
            .O(N__14901),
            .I(\this_vga_ramdac.N_24_mux ));
    InMux I__2105 (
            .O(N__14898),
            .I(N__14895));
    LocalMux I__2104 (
            .O(N__14895),
            .I(N__14892));
    Span4Mux_h I__2103 (
            .O(N__14892),
            .I(N__14888));
    CascadeMux I__2102 (
            .O(N__14891),
            .I(N__14885));
    Span4Mux_h I__2101 (
            .O(N__14888),
            .I(N__14882));
    InMux I__2100 (
            .O(N__14885),
            .I(N__14879));
    Odrv4 I__2099 (
            .O(N__14882),
            .I(\this_vga_ramdac.N_2862_reto ));
    LocalMux I__2098 (
            .O(N__14879),
            .I(\this_vga_ramdac.N_2862_reto ));
    InMux I__2097 (
            .O(N__14874),
            .I(bfn_13_18_0_));
    InMux I__2096 (
            .O(N__14871),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    InMux I__2095 (
            .O(N__14868),
            .I(N__14863));
    InMux I__2094 (
            .O(N__14867),
            .I(N__14860));
    InMux I__2093 (
            .O(N__14866),
            .I(N__14857));
    LocalMux I__2092 (
            .O(N__14863),
            .I(N__14852));
    LocalMux I__2091 (
            .O(N__14860),
            .I(N__14852));
    LocalMux I__2090 (
            .O(N__14857),
            .I(N__14849));
    Span4Mux_v I__2089 (
            .O(N__14852),
            .I(N__14846));
    Span4Mux_h I__2088 (
            .O(N__14849),
            .I(N__14843));
    Odrv4 I__2087 (
            .O(N__14846),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    Odrv4 I__2086 (
            .O(N__14843),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    InMux I__2085 (
            .O(N__14838),
            .I(N__14834));
    InMux I__2084 (
            .O(N__14837),
            .I(N__14831));
    LocalMux I__2083 (
            .O(N__14834),
            .I(N__14826));
    LocalMux I__2082 (
            .O(N__14831),
            .I(N__14826));
    Span4Mux_v I__2081 (
            .O(N__14826),
            .I(N__14822));
    InMux I__2080 (
            .O(N__14825),
            .I(N__14819));
    Odrv4 I__2079 (
            .O(N__14822),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    LocalMux I__2078 (
            .O(N__14819),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    CascadeMux I__2077 (
            .O(N__14814),
            .I(N__14810));
    InMux I__2076 (
            .O(N__14813),
            .I(N__14807));
    InMux I__2075 (
            .O(N__14810),
            .I(N__14804));
    LocalMux I__2074 (
            .O(N__14807),
            .I(N__14799));
    LocalMux I__2073 (
            .O(N__14804),
            .I(N__14799));
    Odrv4 I__2072 (
            .O(N__14799),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    InMux I__2071 (
            .O(N__14796),
            .I(N__14792));
    InMux I__2070 (
            .O(N__14795),
            .I(N__14788));
    LocalMux I__2069 (
            .O(N__14792),
            .I(N__14785));
    InMux I__2068 (
            .O(N__14791),
            .I(N__14782));
    LocalMux I__2067 (
            .O(N__14788),
            .I(N__14779));
    Span4Mux_v I__2066 (
            .O(N__14785),
            .I(N__14774));
    LocalMux I__2065 (
            .O(N__14782),
            .I(N__14774));
    Odrv4 I__2064 (
            .O(N__14779),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    Odrv4 I__2063 (
            .O(N__14774),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    CEMux I__2062 (
            .O(N__14769),
            .I(N__14742));
    CEMux I__2061 (
            .O(N__14768),
            .I(N__14742));
    CEMux I__2060 (
            .O(N__14767),
            .I(N__14742));
    CEMux I__2059 (
            .O(N__14766),
            .I(N__14742));
    CEMux I__2058 (
            .O(N__14765),
            .I(N__14742));
    CEMux I__2057 (
            .O(N__14764),
            .I(N__14742));
    CEMux I__2056 (
            .O(N__14763),
            .I(N__14742));
    CEMux I__2055 (
            .O(N__14762),
            .I(N__14742));
    CEMux I__2054 (
            .O(N__14761),
            .I(N__14742));
    GlobalMux I__2053 (
            .O(N__14742),
            .I(N__14739));
    gio2CtrlBuf I__2052 (
            .O(N__14739),
            .I(\this_vga_signals.N_692_0_g ));
    InMux I__2051 (
            .O(N__14736),
            .I(N__14733));
    LocalMux I__2050 (
            .O(N__14733),
            .I(N__14720));
    SRMux I__2049 (
            .O(N__14732),
            .I(N__14697));
    SRMux I__2048 (
            .O(N__14731),
            .I(N__14697));
    SRMux I__2047 (
            .O(N__14730),
            .I(N__14697));
    SRMux I__2046 (
            .O(N__14729),
            .I(N__14697));
    SRMux I__2045 (
            .O(N__14728),
            .I(N__14697));
    SRMux I__2044 (
            .O(N__14727),
            .I(N__14697));
    SRMux I__2043 (
            .O(N__14726),
            .I(N__14697));
    SRMux I__2042 (
            .O(N__14725),
            .I(N__14697));
    SRMux I__2041 (
            .O(N__14724),
            .I(N__14697));
    SRMux I__2040 (
            .O(N__14723),
            .I(N__14697));
    Glb2LocalMux I__2039 (
            .O(N__14720),
            .I(N__14697));
    GlobalMux I__2038 (
            .O(N__14697),
            .I(N__14694));
    gio2CtrlBuf I__2037 (
            .O(N__14694),
            .I(\this_vga_signals.N_988_g ));
    InMux I__2036 (
            .O(N__14691),
            .I(N__14687));
    InMux I__2035 (
            .O(N__14690),
            .I(N__14684));
    LocalMux I__2034 (
            .O(N__14687),
            .I(N__14681));
    LocalMux I__2033 (
            .O(N__14684),
            .I(N__14675));
    Span4Mux_h I__2032 (
            .O(N__14681),
            .I(N__14672));
    InMux I__2031 (
            .O(N__14680),
            .I(N__14666));
    InMux I__2030 (
            .O(N__14679),
            .I(N__14666));
    InMux I__2029 (
            .O(N__14678),
            .I(N__14660));
    Span4Mux_h I__2028 (
            .O(N__14675),
            .I(N__14655));
    Span4Mux_v I__2027 (
            .O(N__14672),
            .I(N__14655));
    InMux I__2026 (
            .O(N__14671),
            .I(N__14652));
    LocalMux I__2025 (
            .O(N__14666),
            .I(N__14649));
    InMux I__2024 (
            .O(N__14665),
            .I(N__14642));
    InMux I__2023 (
            .O(N__14664),
            .I(N__14642));
    InMux I__2022 (
            .O(N__14663),
            .I(N__14642));
    LocalMux I__2021 (
            .O(N__14660),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__2020 (
            .O(N__14655),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2019 (
            .O(N__14652),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__2018 (
            .O(N__14649),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2017 (
            .O(N__14642),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    InMux I__2016 (
            .O(N__14631),
            .I(N__14628));
    LocalMux I__2015 (
            .O(N__14628),
            .I(N__14625));
    Odrv4 I__2014 (
            .O(N__14625),
            .I(\this_vga_signals.un4_hsynclt8_0 ));
    CascadeMux I__2013 (
            .O(N__14622),
            .I(N__14619));
    InMux I__2012 (
            .O(N__14619),
            .I(N__14616));
    LocalMux I__2011 (
            .O(N__14616),
            .I(N__14613));
    Span4Mux_h I__2010 (
            .O(N__14613),
            .I(N__14610));
    Odrv4 I__2009 (
            .O(N__14610),
            .I(\this_vga_signals.un2_hsynclt8_0 ));
    InMux I__2008 (
            .O(N__14607),
            .I(N__14603));
    CascadeMux I__2007 (
            .O(N__14606),
            .I(N__14598));
    LocalMux I__2006 (
            .O(N__14603),
            .I(N__14593));
    CascadeMux I__2005 (
            .O(N__14602),
            .I(N__14588));
    CascadeMux I__2004 (
            .O(N__14601),
            .I(N__14584));
    InMux I__2003 (
            .O(N__14598),
            .I(N__14581));
    InMux I__2002 (
            .O(N__14597),
            .I(N__14578));
    InMux I__2001 (
            .O(N__14596),
            .I(N__14575));
    Span4Mux_v I__2000 (
            .O(N__14593),
            .I(N__14572));
    InMux I__1999 (
            .O(N__14592),
            .I(N__14569));
    InMux I__1998 (
            .O(N__14591),
            .I(N__14566));
    InMux I__1997 (
            .O(N__14588),
            .I(N__14559));
    InMux I__1996 (
            .O(N__14587),
            .I(N__14559));
    InMux I__1995 (
            .O(N__14584),
            .I(N__14559));
    LocalMux I__1994 (
            .O(N__14581),
            .I(N__14552));
    LocalMux I__1993 (
            .O(N__14578),
            .I(N__14552));
    LocalMux I__1992 (
            .O(N__14575),
            .I(N__14552));
    Odrv4 I__1991 (
            .O(N__14572),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1990 (
            .O(N__14569),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1989 (
            .O(N__14566),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1988 (
            .O(N__14559),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__1987 (
            .O(N__14552),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    IoInMux I__1986 (
            .O(N__14541),
            .I(N__14538));
    LocalMux I__1985 (
            .O(N__14538),
            .I(N__14535));
    Span4Mux_s3_v I__1984 (
            .O(N__14535),
            .I(N__14532));
    Sp12to4 I__1983 (
            .O(N__14532),
            .I(N__14529));
    Span12Mux_h I__1982 (
            .O(N__14529),
            .I(N__14526));
    Odrv12 I__1981 (
            .O(N__14526),
            .I(this_vga_signals_hsync_1_i));
    InMux I__1980 (
            .O(N__14523),
            .I(N__14520));
    LocalMux I__1979 (
            .O(N__14520),
            .I(N__14517));
    Span4Mux_h I__1978 (
            .O(N__14517),
            .I(N__14514));
    Span4Mux_v I__1977 (
            .O(N__14514),
            .I(N__14511));
    Span4Mux_v I__1976 (
            .O(N__14511),
            .I(N__14508));
    Span4Mux_h I__1975 (
            .O(N__14508),
            .I(N__14505));
    Odrv4 I__1974 (
            .O(N__14505),
            .I(M_this_map_ram_read_data_0));
    CascadeMux I__1973 (
            .O(N__14502),
            .I(N__14497));
    CascadeMux I__1972 (
            .O(N__14501),
            .I(N__14491));
    CascadeMux I__1971 (
            .O(N__14500),
            .I(N__14484));
    InMux I__1970 (
            .O(N__14497),
            .I(N__14480));
    CascadeMux I__1969 (
            .O(N__14496),
            .I(N__14477));
    CascadeMux I__1968 (
            .O(N__14495),
            .I(N__14474));
    CascadeMux I__1967 (
            .O(N__14494),
            .I(N__14471));
    InMux I__1966 (
            .O(N__14491),
            .I(N__14466));
    CascadeMux I__1965 (
            .O(N__14490),
            .I(N__14461));
    CascadeMux I__1964 (
            .O(N__14489),
            .I(N__14457));
    CascadeMux I__1963 (
            .O(N__14488),
            .I(N__14454));
    CascadeMux I__1962 (
            .O(N__14487),
            .I(N__14451));
    InMux I__1961 (
            .O(N__14484),
            .I(N__14448));
    CascadeMux I__1960 (
            .O(N__14483),
            .I(N__14445));
    LocalMux I__1959 (
            .O(N__14480),
            .I(N__14442));
    InMux I__1958 (
            .O(N__14477),
            .I(N__14439));
    InMux I__1957 (
            .O(N__14474),
            .I(N__14436));
    InMux I__1956 (
            .O(N__14471),
            .I(N__14433));
    CascadeMux I__1955 (
            .O(N__14470),
            .I(N__14430));
    CascadeMux I__1954 (
            .O(N__14469),
            .I(N__14427));
    LocalMux I__1953 (
            .O(N__14466),
            .I(N__14424));
    CascadeMux I__1952 (
            .O(N__14465),
            .I(N__14421));
    CascadeMux I__1951 (
            .O(N__14464),
            .I(N__14418));
    InMux I__1950 (
            .O(N__14461),
            .I(N__14415));
    CascadeMux I__1949 (
            .O(N__14460),
            .I(N__14412));
    InMux I__1948 (
            .O(N__14457),
            .I(N__14409));
    InMux I__1947 (
            .O(N__14454),
            .I(N__14406));
    InMux I__1946 (
            .O(N__14451),
            .I(N__14403));
    LocalMux I__1945 (
            .O(N__14448),
            .I(N__14400));
    InMux I__1944 (
            .O(N__14445),
            .I(N__14397));
    Span4Mux_h I__1943 (
            .O(N__14442),
            .I(N__14394));
    LocalMux I__1942 (
            .O(N__14439),
            .I(N__14391));
    LocalMux I__1941 (
            .O(N__14436),
            .I(N__14386));
    LocalMux I__1940 (
            .O(N__14433),
            .I(N__14386));
    InMux I__1939 (
            .O(N__14430),
            .I(N__14383));
    InMux I__1938 (
            .O(N__14427),
            .I(N__14380));
    Span4Mux_v I__1937 (
            .O(N__14424),
            .I(N__14377));
    InMux I__1936 (
            .O(N__14421),
            .I(N__14374));
    InMux I__1935 (
            .O(N__14418),
            .I(N__14371));
    LocalMux I__1934 (
            .O(N__14415),
            .I(N__14368));
    InMux I__1933 (
            .O(N__14412),
            .I(N__14365));
    LocalMux I__1932 (
            .O(N__14409),
            .I(N__14362));
    LocalMux I__1931 (
            .O(N__14406),
            .I(N__14359));
    LocalMux I__1930 (
            .O(N__14403),
            .I(N__14356));
    Span4Mux_v I__1929 (
            .O(N__14400),
            .I(N__14351));
    LocalMux I__1928 (
            .O(N__14397),
            .I(N__14351));
    Span4Mux_v I__1927 (
            .O(N__14394),
            .I(N__14348));
    Span4Mux_v I__1926 (
            .O(N__14391),
            .I(N__14341));
    Span4Mux_v I__1925 (
            .O(N__14386),
            .I(N__14341));
    LocalMux I__1924 (
            .O(N__14383),
            .I(N__14341));
    LocalMux I__1923 (
            .O(N__14380),
            .I(N__14338));
    Span4Mux_h I__1922 (
            .O(N__14377),
            .I(N__14335));
    LocalMux I__1921 (
            .O(N__14374),
            .I(N__14328));
    LocalMux I__1920 (
            .O(N__14371),
            .I(N__14328));
    Sp12to4 I__1919 (
            .O(N__14368),
            .I(N__14328));
    LocalMux I__1918 (
            .O(N__14365),
            .I(N__14325));
    Span12Mux_h I__1917 (
            .O(N__14362),
            .I(N__14322));
    Span4Mux_v I__1916 (
            .O(N__14359),
            .I(N__14319));
    Span4Mux_v I__1915 (
            .O(N__14356),
            .I(N__14314));
    Span4Mux_v I__1914 (
            .O(N__14351),
            .I(N__14314));
    Sp12to4 I__1913 (
            .O(N__14348),
            .I(N__14309));
    Sp12to4 I__1912 (
            .O(N__14341),
            .I(N__14309));
    Sp12to4 I__1911 (
            .O(N__14338),
            .I(N__14302));
    Sp12to4 I__1910 (
            .O(N__14335),
            .I(N__14302));
    Span12Mux_s11_v I__1909 (
            .O(N__14328),
            .I(N__14302));
    Span12Mux_s9_h I__1908 (
            .O(N__14325),
            .I(N__14299));
    Span12Mux_v I__1907 (
            .O(N__14322),
            .I(N__14296));
    Span4Mux_h I__1906 (
            .O(N__14319),
            .I(N__14291));
    Span4Mux_h I__1905 (
            .O(N__14314),
            .I(N__14291));
    Span12Mux_h I__1904 (
            .O(N__14309),
            .I(N__14286));
    Span12Mux_h I__1903 (
            .O(N__14302),
            .I(N__14286));
    Odrv12 I__1902 (
            .O(N__14299),
            .I(M_this_ppu_sprites_addr_6));
    Odrv12 I__1901 (
            .O(N__14296),
            .I(M_this_ppu_sprites_addr_6));
    Odrv4 I__1900 (
            .O(N__14291),
            .I(M_this_ppu_sprites_addr_6));
    Odrv12 I__1899 (
            .O(N__14286),
            .I(M_this_ppu_sprites_addr_6));
    InMux I__1898 (
            .O(N__14277),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    InMux I__1897 (
            .O(N__14274),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__1896 (
            .O(N__14271),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__1895 (
            .O(N__14268),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__1894 (
            .O(N__14265),
            .I(N__14259));
    InMux I__1893 (
            .O(N__14264),
            .I(N__14259));
    LocalMux I__1892 (
            .O(N__14259),
            .I(N__14255));
    InMux I__1891 (
            .O(N__14258),
            .I(N__14252));
    Span4Mux_v I__1890 (
            .O(N__14255),
            .I(N__14247));
    LocalMux I__1889 (
            .O(N__14252),
            .I(N__14247));
    Odrv4 I__1888 (
            .O(N__14247),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    InMux I__1887 (
            .O(N__14244),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__1886 (
            .O(N__14241),
            .I(N__14237));
    InMux I__1885 (
            .O(N__14240),
            .I(N__14234));
    LocalMux I__1884 (
            .O(N__14237),
            .I(N__14230));
    LocalMux I__1883 (
            .O(N__14234),
            .I(N__14227));
    InMux I__1882 (
            .O(N__14233),
            .I(N__14224));
    Span4Mux_h I__1881 (
            .O(N__14230),
            .I(N__14221));
    Span4Mux_h I__1880 (
            .O(N__14227),
            .I(N__14218));
    LocalMux I__1879 (
            .O(N__14224),
            .I(N__14215));
    Odrv4 I__1878 (
            .O(N__14221),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    Odrv4 I__1877 (
            .O(N__14218),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    Odrv12 I__1876 (
            .O(N__14215),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    InMux I__1875 (
            .O(N__14208),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__1874 (
            .O(N__14205),
            .I(N__14202));
    LocalMux I__1873 (
            .O(N__14202),
            .I(N__14198));
    InMux I__1872 (
            .O(N__14201),
            .I(N__14195));
    Span4Mux_h I__1871 (
            .O(N__14198),
            .I(N__14192));
    LocalMux I__1870 (
            .O(N__14195),
            .I(N__14189));
    Odrv4 I__1869 (
            .O(N__14192),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    Odrv12 I__1868 (
            .O(N__14189),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    InMux I__1867 (
            .O(N__14184),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    CascadeMux I__1866 (
            .O(N__14181),
            .I(N__14178));
    InMux I__1865 (
            .O(N__14178),
            .I(N__14175));
    LocalMux I__1864 (
            .O(N__14175),
            .I(N__14168));
    InMux I__1863 (
            .O(N__14174),
            .I(N__14165));
    CascadeMux I__1862 (
            .O(N__14173),
            .I(N__14161));
    InMux I__1861 (
            .O(N__14172),
            .I(N__14155));
    InMux I__1860 (
            .O(N__14171),
            .I(N__14152));
    Span4Mux_h I__1859 (
            .O(N__14168),
            .I(N__14149));
    LocalMux I__1858 (
            .O(N__14165),
            .I(N__14146));
    InMux I__1857 (
            .O(N__14164),
            .I(N__14139));
    InMux I__1856 (
            .O(N__14161),
            .I(N__14139));
    InMux I__1855 (
            .O(N__14160),
            .I(N__14139));
    InMux I__1854 (
            .O(N__14159),
            .I(N__14134));
    InMux I__1853 (
            .O(N__14158),
            .I(N__14134));
    LocalMux I__1852 (
            .O(N__14155),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1851 (
            .O(N__14152),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__1850 (
            .O(N__14149),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__1849 (
            .O(N__14146),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1848 (
            .O(N__14139),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1847 (
            .O(N__14134),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__1846 (
            .O(N__14121),
            .I(N__14115));
    InMux I__1845 (
            .O(N__14120),
            .I(N__14115));
    LocalMux I__1844 (
            .O(N__14115),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ));
    CascadeMux I__1843 (
            .O(N__14112),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_ ));
    InMux I__1842 (
            .O(N__14109),
            .I(N__14106));
    LocalMux I__1841 (
            .O(N__14106),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0_0_0 ));
    CascadeMux I__1840 (
            .O(N__14103),
            .I(N__14097));
    CascadeMux I__1839 (
            .O(N__14102),
            .I(N__14094));
    CascadeMux I__1838 (
            .O(N__14101),
            .I(N__14090));
    InMux I__1837 (
            .O(N__14100),
            .I(N__14084));
    InMux I__1836 (
            .O(N__14097),
            .I(N__14079));
    InMux I__1835 (
            .O(N__14094),
            .I(N__14079));
    InMux I__1834 (
            .O(N__14093),
            .I(N__14074));
    InMux I__1833 (
            .O(N__14090),
            .I(N__14074));
    InMux I__1832 (
            .O(N__14089),
            .I(N__14070));
    InMux I__1831 (
            .O(N__14088),
            .I(N__14067));
    InMux I__1830 (
            .O(N__14087),
            .I(N__14064));
    LocalMux I__1829 (
            .O(N__14084),
            .I(N__14057));
    LocalMux I__1828 (
            .O(N__14079),
            .I(N__14057));
    LocalMux I__1827 (
            .O(N__14074),
            .I(N__14057));
    InMux I__1826 (
            .O(N__14073),
            .I(N__14054));
    LocalMux I__1825 (
            .O(N__14070),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1824 (
            .O(N__14067),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1823 (
            .O(N__14064),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1822 (
            .O(N__14057),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1821 (
            .O(N__14054),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__1820 (
            .O(N__14043),
            .I(N__14033));
    InMux I__1819 (
            .O(N__14042),
            .I(N__14033));
    InMux I__1818 (
            .O(N__14041),
            .I(N__14028));
    InMux I__1817 (
            .O(N__14040),
            .I(N__14028));
    InMux I__1816 (
            .O(N__14039),
            .I(N__14024));
    InMux I__1815 (
            .O(N__14038),
            .I(N__14021));
    LocalMux I__1814 (
            .O(N__14033),
            .I(N__14018));
    LocalMux I__1813 (
            .O(N__14028),
            .I(N__14015));
    InMux I__1812 (
            .O(N__14027),
            .I(N__14012));
    LocalMux I__1811 (
            .O(N__14024),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__1810 (
            .O(N__14021),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1809 (
            .O(N__14018),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1808 (
            .O(N__14015),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__1807 (
            .O(N__14012),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__1806 (
            .O(N__14001),
            .I(N__13995));
    InMux I__1805 (
            .O(N__14000),
            .I(N__13991));
    CascadeMux I__1804 (
            .O(N__13999),
            .I(N__13987));
    CascadeMux I__1803 (
            .O(N__13998),
            .I(N__13984));
    LocalMux I__1802 (
            .O(N__13995),
            .I(N__13981));
    CascadeMux I__1801 (
            .O(N__13994),
            .I(N__13977));
    LocalMux I__1800 (
            .O(N__13991),
            .I(N__13974));
    InMux I__1799 (
            .O(N__13990),
            .I(N__13971));
    InMux I__1798 (
            .O(N__13987),
            .I(N__13966));
    InMux I__1797 (
            .O(N__13984),
            .I(N__13966));
    Span4Mux_v I__1796 (
            .O(N__13981),
            .I(N__13963));
    InMux I__1795 (
            .O(N__13980),
            .I(N__13960));
    InMux I__1794 (
            .O(N__13977),
            .I(N__13957));
    Span4Mux_h I__1793 (
            .O(N__13974),
            .I(N__13954));
    LocalMux I__1792 (
            .O(N__13971),
            .I(N__13949));
    LocalMux I__1791 (
            .O(N__13966),
            .I(N__13949));
    Odrv4 I__1790 (
            .O(N__13963),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__1789 (
            .O(N__13960),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__1788 (
            .O(N__13957),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__1787 (
            .O(N__13954),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__1786 (
            .O(N__13949),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    InMux I__1785 (
            .O(N__13938),
            .I(N__13934));
    InMux I__1784 (
            .O(N__13937),
            .I(N__13921));
    LocalMux I__1783 (
            .O(N__13934),
            .I(N__13918));
    InMux I__1782 (
            .O(N__13933),
            .I(N__13913));
    InMux I__1781 (
            .O(N__13932),
            .I(N__13913));
    InMux I__1780 (
            .O(N__13931),
            .I(N__13908));
    InMux I__1779 (
            .O(N__13930),
            .I(N__13908));
    InMux I__1778 (
            .O(N__13929),
            .I(N__13895));
    InMux I__1777 (
            .O(N__13928),
            .I(N__13895));
    InMux I__1776 (
            .O(N__13927),
            .I(N__13895));
    InMux I__1775 (
            .O(N__13926),
            .I(N__13895));
    InMux I__1774 (
            .O(N__13925),
            .I(N__13895));
    InMux I__1773 (
            .O(N__13924),
            .I(N__13895));
    LocalMux I__1772 (
            .O(N__13921),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1771 (
            .O(N__13918),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1770 (
            .O(N__13913),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1769 (
            .O(N__13908),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1768 (
            .O(N__13895),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    CascadeMux I__1767 (
            .O(N__13884),
            .I(N__13874));
    CascadeMux I__1766 (
            .O(N__13883),
            .I(N__13871));
    InMux I__1765 (
            .O(N__13882),
            .I(N__13866));
    InMux I__1764 (
            .O(N__13881),
            .I(N__13861));
    InMux I__1763 (
            .O(N__13880),
            .I(N__13861));
    InMux I__1762 (
            .O(N__13879),
            .I(N__13858));
    InMux I__1761 (
            .O(N__13878),
            .I(N__13849));
    InMux I__1760 (
            .O(N__13877),
            .I(N__13849));
    InMux I__1759 (
            .O(N__13874),
            .I(N__13849));
    InMux I__1758 (
            .O(N__13871),
            .I(N__13849));
    InMux I__1757 (
            .O(N__13870),
            .I(N__13844));
    InMux I__1756 (
            .O(N__13869),
            .I(N__13844));
    LocalMux I__1755 (
            .O(N__13866),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1754 (
            .O(N__13861),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1753 (
            .O(N__13858),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1752 (
            .O(N__13849),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1751 (
            .O(N__13844),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    CascadeMux I__1750 (
            .O(N__13833),
            .I(\this_vga_signals.un4_hsynclt4_0_cascade_ ));
    InMux I__1749 (
            .O(N__13830),
            .I(N__13821));
    InMux I__1748 (
            .O(N__13829),
            .I(N__13816));
    InMux I__1747 (
            .O(N__13828),
            .I(N__13816));
    InMux I__1746 (
            .O(N__13827),
            .I(N__13811));
    InMux I__1745 (
            .O(N__13826),
            .I(N__13811));
    InMux I__1744 (
            .O(N__13825),
            .I(N__13802));
    InMux I__1743 (
            .O(N__13824),
            .I(N__13799));
    LocalMux I__1742 (
            .O(N__13821),
            .I(N__13796));
    LocalMux I__1741 (
            .O(N__13816),
            .I(N__13793));
    LocalMux I__1740 (
            .O(N__13811),
            .I(N__13790));
    InMux I__1739 (
            .O(N__13810),
            .I(N__13783));
    InMux I__1738 (
            .O(N__13809),
            .I(N__13783));
    InMux I__1737 (
            .O(N__13808),
            .I(N__13783));
    InMux I__1736 (
            .O(N__13807),
            .I(N__13776));
    InMux I__1735 (
            .O(N__13806),
            .I(N__13776));
    InMux I__1734 (
            .O(N__13805),
            .I(N__13776));
    LocalMux I__1733 (
            .O(N__13802),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1732 (
            .O(N__13799),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1731 (
            .O(N__13796),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1730 (
            .O(N__13793),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1729 (
            .O(N__13790),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1728 (
            .O(N__13783),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1727 (
            .O(N__13776),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__1726 (
            .O(N__13761),
            .I(N__13758));
    LocalMux I__1725 (
            .O(N__13758),
            .I(N__13755));
    Odrv12 I__1724 (
            .O(N__13755),
            .I(N_91_0));
    InMux I__1723 (
            .O(N__13752),
            .I(N__13749));
    LocalMux I__1722 (
            .O(N__13749),
            .I(N__13746));
    Span4Mux_h I__1721 (
            .O(N__13746),
            .I(N__13743));
    Odrv4 I__1720 (
            .O(N__13743),
            .I(N_93_0));
    InMux I__1719 (
            .O(N__13740),
            .I(N__13737));
    LocalMux I__1718 (
            .O(N__13737),
            .I(N__13734));
    Sp12to4 I__1717 (
            .O(N__13734),
            .I(N__13731));
    Span12Mux_v I__1716 (
            .O(N__13731),
            .I(N__13728));
    Odrv12 I__1715 (
            .O(N__13728),
            .I(M_this_map_ram_read_data_3));
    CascadeMux I__1714 (
            .O(N__13725),
            .I(N__13721));
    CascadeMux I__1713 (
            .O(N__13724),
            .I(N__13718));
    InMux I__1712 (
            .O(N__13721),
            .I(N__13712));
    InMux I__1711 (
            .O(N__13718),
            .I(N__13708));
    CascadeMux I__1710 (
            .O(N__13717),
            .I(N__13705));
    CascadeMux I__1709 (
            .O(N__13716),
            .I(N__13701));
    CascadeMux I__1708 (
            .O(N__13715),
            .I(N__13697));
    LocalMux I__1707 (
            .O(N__13712),
            .I(N__13692));
    CascadeMux I__1706 (
            .O(N__13711),
            .I(N__13689));
    LocalMux I__1705 (
            .O(N__13708),
            .I(N__13685));
    InMux I__1704 (
            .O(N__13705),
            .I(N__13682));
    CascadeMux I__1703 (
            .O(N__13704),
            .I(N__13679));
    InMux I__1702 (
            .O(N__13701),
            .I(N__13675));
    CascadeMux I__1701 (
            .O(N__13700),
            .I(N__13672));
    InMux I__1700 (
            .O(N__13697),
            .I(N__13667));
    CascadeMux I__1699 (
            .O(N__13696),
            .I(N__13664));
    CascadeMux I__1698 (
            .O(N__13695),
            .I(N__13661));
    Span4Mux_v I__1697 (
            .O(N__13692),
            .I(N__13658));
    InMux I__1696 (
            .O(N__13689),
            .I(N__13655));
    CascadeMux I__1695 (
            .O(N__13688),
            .I(N__13652));
    Span4Mux_v I__1694 (
            .O(N__13685),
            .I(N__13647));
    LocalMux I__1693 (
            .O(N__13682),
            .I(N__13647));
    InMux I__1692 (
            .O(N__13679),
            .I(N__13644));
    CascadeMux I__1691 (
            .O(N__13678),
            .I(N__13641));
    LocalMux I__1690 (
            .O(N__13675),
            .I(N__13638));
    InMux I__1689 (
            .O(N__13672),
            .I(N__13635));
    CascadeMux I__1688 (
            .O(N__13671),
            .I(N__13632));
    CascadeMux I__1687 (
            .O(N__13670),
            .I(N__13628));
    LocalMux I__1686 (
            .O(N__13667),
            .I(N__13625));
    InMux I__1685 (
            .O(N__13664),
            .I(N__13622));
    InMux I__1684 (
            .O(N__13661),
            .I(N__13619));
    Span4Mux_v I__1683 (
            .O(N__13658),
            .I(N__13616));
    LocalMux I__1682 (
            .O(N__13655),
            .I(N__13613));
    InMux I__1681 (
            .O(N__13652),
            .I(N__13610));
    Span4Mux_h I__1680 (
            .O(N__13647),
            .I(N__13605));
    LocalMux I__1679 (
            .O(N__13644),
            .I(N__13605));
    InMux I__1678 (
            .O(N__13641),
            .I(N__13602));
    Span4Mux_h I__1677 (
            .O(N__13638),
            .I(N__13596));
    LocalMux I__1676 (
            .O(N__13635),
            .I(N__13596));
    InMux I__1675 (
            .O(N__13632),
            .I(N__13593));
    CascadeMux I__1674 (
            .O(N__13631),
            .I(N__13590));
    InMux I__1673 (
            .O(N__13628),
            .I(N__13587));
    Span4Mux_h I__1672 (
            .O(N__13625),
            .I(N__13584));
    LocalMux I__1671 (
            .O(N__13622),
            .I(N__13581));
    LocalMux I__1670 (
            .O(N__13619),
            .I(N__13578));
    Span4Mux_v I__1669 (
            .O(N__13616),
            .I(N__13571));
    Span4Mux_v I__1668 (
            .O(N__13613),
            .I(N__13571));
    LocalMux I__1667 (
            .O(N__13610),
            .I(N__13571));
    Span4Mux_v I__1666 (
            .O(N__13605),
            .I(N__13566));
    LocalMux I__1665 (
            .O(N__13602),
            .I(N__13566));
    CascadeMux I__1664 (
            .O(N__13601),
            .I(N__13563));
    Span4Mux_v I__1663 (
            .O(N__13596),
            .I(N__13558));
    LocalMux I__1662 (
            .O(N__13593),
            .I(N__13558));
    InMux I__1661 (
            .O(N__13590),
            .I(N__13555));
    LocalMux I__1660 (
            .O(N__13587),
            .I(N__13552));
    Span4Mux_v I__1659 (
            .O(N__13584),
            .I(N__13547));
    Span4Mux_h I__1658 (
            .O(N__13581),
            .I(N__13547));
    Span4Mux_h I__1657 (
            .O(N__13578),
            .I(N__13544));
    Span4Mux_v I__1656 (
            .O(N__13571),
            .I(N__13539));
    Span4Mux_v I__1655 (
            .O(N__13566),
            .I(N__13539));
    InMux I__1654 (
            .O(N__13563),
            .I(N__13536));
    Span4Mux_v I__1653 (
            .O(N__13558),
            .I(N__13531));
    LocalMux I__1652 (
            .O(N__13555),
            .I(N__13531));
    Span12Mux_s9_h I__1651 (
            .O(N__13552),
            .I(N__13526));
    Sp12to4 I__1650 (
            .O(N__13547),
            .I(N__13526));
    Span4Mux_v I__1649 (
            .O(N__13544),
            .I(N__13521));
    Span4Mux_h I__1648 (
            .O(N__13539),
            .I(N__13521));
    LocalMux I__1647 (
            .O(N__13536),
            .I(N__13518));
    Span4Mux_h I__1646 (
            .O(N__13531),
            .I(N__13515));
    Span12Mux_v I__1645 (
            .O(N__13526),
            .I(N__13508));
    Sp12to4 I__1644 (
            .O(N__13521),
            .I(N__13508));
    Span12Mux_s9_h I__1643 (
            .O(N__13518),
            .I(N__13508));
    Span4Mux_h I__1642 (
            .O(N__13515),
            .I(N__13505));
    Odrv12 I__1641 (
            .O(N__13508),
            .I(M_this_ppu_sprites_addr_9));
    Odrv4 I__1640 (
            .O(N__13505),
            .I(M_this_ppu_sprites_addr_9));
    CascadeMux I__1639 (
            .O(N__13500),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ));
    CascadeMux I__1638 (
            .O(N__13497),
            .I(N__13494));
    InMux I__1637 (
            .O(N__13494),
            .I(N__13485));
    InMux I__1636 (
            .O(N__13493),
            .I(N__13485));
    InMux I__1635 (
            .O(N__13492),
            .I(N__13485));
    LocalMux I__1634 (
            .O(N__13485),
            .I(\this_vga_signals.mult1_un68_sum_axb2_1 ));
    CascadeMux I__1633 (
            .O(N__13482),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1_cascade_ ));
    CascadeMux I__1632 (
            .O(N__13479),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_ ));
    InMux I__1631 (
            .O(N__13476),
            .I(N__13473));
    LocalMux I__1630 (
            .O(N__13473),
            .I(N__13470));
    Span4Mux_h I__1629 (
            .O(N__13470),
            .I(N__13467));
    Span4Mux_v I__1628 (
            .O(N__13467),
            .I(N__13460));
    InMux I__1627 (
            .O(N__13466),
            .I(N__13455));
    InMux I__1626 (
            .O(N__13465),
            .I(N__13455));
    InMux I__1625 (
            .O(N__13464),
            .I(N__13450));
    InMux I__1624 (
            .O(N__13463),
            .I(N__13450));
    Odrv4 I__1623 (
            .O(N__13460),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1622 (
            .O(N__13455),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1621 (
            .O(N__13450),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    CascadeMux I__1620 (
            .O(N__13443),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_ ));
    InMux I__1619 (
            .O(N__13440),
            .I(N__13437));
    LocalMux I__1618 (
            .O(N__13437),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_0 ));
    InMux I__1617 (
            .O(N__13434),
            .I(N__13431));
    LocalMux I__1616 (
            .O(N__13431),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    CascadeMux I__1615 (
            .O(N__13428),
            .I(N__13425));
    InMux I__1614 (
            .O(N__13425),
            .I(N__13422));
    LocalMux I__1613 (
            .O(N__13422),
            .I(N__13419));
    Span12Mux_s11_h I__1612 (
            .O(N__13419),
            .I(N__13416));
    Odrv12 I__1611 (
            .O(N__13416),
            .I(M_this_vga_signals_address_5));
    InMux I__1610 (
            .O(N__13413),
            .I(N__13407));
    InMux I__1609 (
            .O(N__13412),
            .I(N__13407));
    LocalMux I__1608 (
            .O(N__13407),
            .I(\this_vga_signals.SUM_3 ));
    CascadeMux I__1607 (
            .O(N__13404),
            .I(\this_vga_signals.SUM_3_cascade_ ));
    InMux I__1606 (
            .O(N__13401),
            .I(N__13398));
    LocalMux I__1605 (
            .O(N__13398),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0 ));
    InMux I__1604 (
            .O(N__13395),
            .I(N__13392));
    LocalMux I__1603 (
            .O(N__13392),
            .I(\this_vga_signals.N_6_1 ));
    InMux I__1602 (
            .O(N__13389),
            .I(N__13378));
    InMux I__1601 (
            .O(N__13388),
            .I(N__13378));
    InMux I__1600 (
            .O(N__13387),
            .I(N__13370));
    InMux I__1599 (
            .O(N__13386),
            .I(N__13370));
    InMux I__1598 (
            .O(N__13385),
            .I(N__13370));
    InMux I__1597 (
            .O(N__13384),
            .I(N__13358));
    InMux I__1596 (
            .O(N__13383),
            .I(N__13355));
    LocalMux I__1595 (
            .O(N__13378),
            .I(N__13352));
    InMux I__1594 (
            .O(N__13377),
            .I(N__13349));
    LocalMux I__1593 (
            .O(N__13370),
            .I(N__13346));
    InMux I__1592 (
            .O(N__13369),
            .I(N__13339));
    InMux I__1591 (
            .O(N__13368),
            .I(N__13339));
    InMux I__1590 (
            .O(N__13367),
            .I(N__13339));
    InMux I__1589 (
            .O(N__13366),
            .I(N__13332));
    InMux I__1588 (
            .O(N__13365),
            .I(N__13332));
    InMux I__1587 (
            .O(N__13364),
            .I(N__13332));
    InMux I__1586 (
            .O(N__13363),
            .I(N__13325));
    InMux I__1585 (
            .O(N__13362),
            .I(N__13325));
    InMux I__1584 (
            .O(N__13361),
            .I(N__13325));
    LocalMux I__1583 (
            .O(N__13358),
            .I(\this_vga_signals.mult1_un68_sum_axb1_571 ));
    LocalMux I__1582 (
            .O(N__13355),
            .I(\this_vga_signals.mult1_un68_sum_axb1_571 ));
    Odrv4 I__1581 (
            .O(N__13352),
            .I(\this_vga_signals.mult1_un68_sum_axb1_571 ));
    LocalMux I__1580 (
            .O(N__13349),
            .I(\this_vga_signals.mult1_un68_sum_axb1_571 ));
    Odrv4 I__1579 (
            .O(N__13346),
            .I(\this_vga_signals.mult1_un68_sum_axb1_571 ));
    LocalMux I__1578 (
            .O(N__13339),
            .I(\this_vga_signals.mult1_un68_sum_axb1_571 ));
    LocalMux I__1577 (
            .O(N__13332),
            .I(\this_vga_signals.mult1_un68_sum_axb1_571 ));
    LocalMux I__1576 (
            .O(N__13325),
            .I(\this_vga_signals.mult1_un68_sum_axb1_571 ));
    CascadeMux I__1575 (
            .O(N__13308),
            .I(N__13303));
    InMux I__1574 (
            .O(N__13307),
            .I(N__13300));
    InMux I__1573 (
            .O(N__13306),
            .I(N__13290));
    InMux I__1572 (
            .O(N__13303),
            .I(N__13287));
    LocalMux I__1571 (
            .O(N__13300),
            .I(N__13284));
    InMux I__1570 (
            .O(N__13299),
            .I(N__13277));
    InMux I__1569 (
            .O(N__13298),
            .I(N__13277));
    InMux I__1568 (
            .O(N__13297),
            .I(N__13277));
    CascadeMux I__1567 (
            .O(N__13296),
            .I(N__13271));
    CascadeMux I__1566 (
            .O(N__13295),
            .I(N__13265));
    InMux I__1565 (
            .O(N__13294),
            .I(N__13261));
    InMux I__1564 (
            .O(N__13293),
            .I(N__13258));
    LocalMux I__1563 (
            .O(N__13290),
            .I(N__13251));
    LocalMux I__1562 (
            .O(N__13287),
            .I(N__13251));
    Span4Mux_h I__1561 (
            .O(N__13284),
            .I(N__13251));
    LocalMux I__1560 (
            .O(N__13277),
            .I(N__13248));
    InMux I__1559 (
            .O(N__13276),
            .I(N__13245));
    InMux I__1558 (
            .O(N__13275),
            .I(N__13236));
    InMux I__1557 (
            .O(N__13274),
            .I(N__13236));
    InMux I__1556 (
            .O(N__13271),
            .I(N__13236));
    InMux I__1555 (
            .O(N__13270),
            .I(N__13236));
    InMux I__1554 (
            .O(N__13269),
            .I(N__13227));
    InMux I__1553 (
            .O(N__13268),
            .I(N__13227));
    InMux I__1552 (
            .O(N__13265),
            .I(N__13227));
    InMux I__1551 (
            .O(N__13264),
            .I(N__13227));
    LocalMux I__1550 (
            .O(N__13261),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1549 (
            .O(N__13258),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    Odrv4 I__1548 (
            .O(N__13251),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    Odrv4 I__1547 (
            .O(N__13248),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1546 (
            .O(N__13245),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1545 (
            .O(N__13236),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1544 (
            .O(N__13227),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    InMux I__1543 (
            .O(N__13212),
            .I(N__13208));
    InMux I__1542 (
            .O(N__13211),
            .I(N__13205));
    LocalMux I__1541 (
            .O(N__13208),
            .I(N__13202));
    LocalMux I__1540 (
            .O(N__13205),
            .I(\this_vga_signals.N_4_0_0_1 ));
    Odrv4 I__1539 (
            .O(N__13202),
            .I(\this_vga_signals.N_4_0_0_1 ));
    CascadeMux I__1538 (
            .O(N__13197),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_cascade_ ));
    CascadeMux I__1537 (
            .O(N__13194),
            .I(N__13191));
    InMux I__1536 (
            .O(N__13191),
            .I(N__13188));
    LocalMux I__1535 (
            .O(N__13188),
            .I(N__13185));
    Span4Mux_h I__1534 (
            .O(N__13185),
            .I(N__13182));
    Odrv4 I__1533 (
            .O(N__13182),
            .I(M_this_vga_signals_address_3));
    InMux I__1532 (
            .O(N__13179),
            .I(N__13176));
    LocalMux I__1531 (
            .O(N__13176),
            .I(\this_vga_signals.if_m2_0 ));
    InMux I__1530 (
            .O(N__13173),
            .I(N__13167));
    InMux I__1529 (
            .O(N__13172),
            .I(N__13167));
    LocalMux I__1528 (
            .O(N__13167),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    InMux I__1527 (
            .O(N__13164),
            .I(N__13161));
    LocalMux I__1526 (
            .O(N__13161),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1 ));
    CascadeMux I__1525 (
            .O(N__13158),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ));
    InMux I__1524 (
            .O(N__13155),
            .I(N__13152));
    LocalMux I__1523 (
            .O(N__13152),
            .I(\this_vga_signals.mult1_un82_sum_c3_0 ));
    InMux I__1522 (
            .O(N__13149),
            .I(N__13144));
    InMux I__1521 (
            .O(N__13148),
            .I(N__13139));
    InMux I__1520 (
            .O(N__13147),
            .I(N__13139));
    LocalMux I__1519 (
            .O(N__13144),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0 ));
    LocalMux I__1518 (
            .O(N__13139),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0 ));
    CascadeMux I__1517 (
            .O(N__13134),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_cascade_ ));
    InMux I__1516 (
            .O(N__13131),
            .I(N__13128));
    LocalMux I__1515 (
            .O(N__13128),
            .I(N__13125));
    Span4Mux_h I__1514 (
            .O(N__13125),
            .I(N__13122));
    Span4Mux_h I__1513 (
            .O(N__13122),
            .I(N__13117));
    InMux I__1512 (
            .O(N__13121),
            .I(N__13114));
    InMux I__1511 (
            .O(N__13120),
            .I(N__13111));
    Odrv4 I__1510 (
            .O(N__13117),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__1509 (
            .O(N__13114),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__1508 (
            .O(N__13111),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    CascadeMux I__1507 (
            .O(N__13104),
            .I(N__13101));
    InMux I__1506 (
            .O(N__13101),
            .I(N__13098));
    LocalMux I__1505 (
            .O(N__13098),
            .I(N__13095));
    Span4Mux_h I__1504 (
            .O(N__13095),
            .I(N__13092));
    Odrv4 I__1503 (
            .O(N__13092),
            .I(M_this_vga_signals_address_1));
    InMux I__1502 (
            .O(N__13089),
            .I(N__13082));
    InMux I__1501 (
            .O(N__13088),
            .I(N__13082));
    InMux I__1500 (
            .O(N__13087),
            .I(N__13079));
    LocalMux I__1499 (
            .O(N__13082),
            .I(N__13076));
    LocalMux I__1498 (
            .O(N__13079),
            .I(\this_vga_signals.mult1_un75_sum_axb1 ));
    Odrv4 I__1497 (
            .O(N__13076),
            .I(\this_vga_signals.mult1_un75_sum_axb1 ));
    InMux I__1496 (
            .O(N__13071),
            .I(N__13067));
    InMux I__1495 (
            .O(N__13070),
            .I(N__13064));
    LocalMux I__1494 (
            .O(N__13067),
            .I(\this_vga_signals.mult1_un68_sum_ac0_2 ));
    LocalMux I__1493 (
            .O(N__13064),
            .I(\this_vga_signals.mult1_un68_sum_ac0_2 ));
    CascadeMux I__1492 (
            .O(N__13059),
            .I(\this_vga_signals.g2_0_0_cascade_ ));
    InMux I__1491 (
            .O(N__13056),
            .I(N__13053));
    LocalMux I__1490 (
            .O(N__13053),
            .I(\this_vga_signals.g0_0_0_a3_0 ));
    InMux I__1489 (
            .O(N__13050),
            .I(N__13047));
    LocalMux I__1488 (
            .O(N__13047),
            .I(N__13044));
    Span4Mux_h I__1487 (
            .O(N__13044),
            .I(N__13040));
    InMux I__1486 (
            .O(N__13043),
            .I(N__13037));
    Odrv4 I__1485 (
            .O(N__13040),
            .I(\this_vga_signals.vaddress_c3_0 ));
    LocalMux I__1484 (
            .O(N__13037),
            .I(\this_vga_signals.vaddress_c3_0 ));
    CascadeMux I__1483 (
            .O(N__13032),
            .I(N__13029));
    InMux I__1482 (
            .O(N__13029),
            .I(N__13026));
    LocalMux I__1481 (
            .O(N__13026),
            .I(N__13022));
    InMux I__1480 (
            .O(N__13025),
            .I(N__13019));
    Span4Mux_h I__1479 (
            .O(N__13022),
            .I(N__13014));
    LocalMux I__1478 (
            .O(N__13019),
            .I(N__13014));
    Odrv4 I__1477 (
            .O(N__13014),
            .I(\this_vga_signals.SUM_2_i_1_1_3 ));
    InMux I__1476 (
            .O(N__13011),
            .I(N__13008));
    LocalMux I__1475 (
            .O(N__13008),
            .I(N__13005));
    Span4Mux_h I__1474 (
            .O(N__13005),
            .I(N__13001));
    InMux I__1473 (
            .O(N__13004),
            .I(N__12998));
    Odrv4 I__1472 (
            .O(N__13001),
            .I(\this_vga_signals.SUM_2_i_1_2_3 ));
    LocalMux I__1471 (
            .O(N__12998),
            .I(\this_vga_signals.SUM_2_i_1_2_3 ));
    CascadeMux I__1470 (
            .O(N__12993),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i_0_cascade_ ));
    InMux I__1469 (
            .O(N__12990),
            .I(N__12987));
    LocalMux I__1468 (
            .O(N__12987),
            .I(\this_vga_signals.g0_i_x4_0 ));
    CascadeMux I__1467 (
            .O(N__12984),
            .I(\this_vga_signals.g0_i_x4_4_1_cascade_ ));
    InMux I__1466 (
            .O(N__12981),
            .I(N__12978));
    LocalMux I__1465 (
            .O(N__12978),
            .I(N__12975));
    Span4Mux_h I__1464 (
            .O(N__12975),
            .I(N__12972));
    Odrv4 I__1463 (
            .O(N__12972),
            .I(\this_vga_signals.g0_i_x4_4 ));
    InMux I__1462 (
            .O(N__12969),
            .I(N__12958));
    InMux I__1461 (
            .O(N__12968),
            .I(N__12958));
    InMux I__1460 (
            .O(N__12967),
            .I(N__12955));
    InMux I__1459 (
            .O(N__12966),
            .I(N__12950));
    InMux I__1458 (
            .O(N__12965),
            .I(N__12950));
    CascadeMux I__1457 (
            .O(N__12964),
            .I(N__12946));
    CascadeMux I__1456 (
            .O(N__12963),
            .I(N__12940));
    LocalMux I__1455 (
            .O(N__12958),
            .I(N__12932));
    LocalMux I__1454 (
            .O(N__12955),
            .I(N__12932));
    LocalMux I__1453 (
            .O(N__12950),
            .I(N__12929));
    InMux I__1452 (
            .O(N__12949),
            .I(N__12926));
    InMux I__1451 (
            .O(N__12946),
            .I(N__12921));
    InMux I__1450 (
            .O(N__12945),
            .I(N__12921));
    InMux I__1449 (
            .O(N__12944),
            .I(N__12918));
    InMux I__1448 (
            .O(N__12943),
            .I(N__12911));
    InMux I__1447 (
            .O(N__12940),
            .I(N__12911));
    InMux I__1446 (
            .O(N__12939),
            .I(N__12911));
    InMux I__1445 (
            .O(N__12938),
            .I(N__12908));
    InMux I__1444 (
            .O(N__12937),
            .I(N__12905));
    Span4Mux_v I__1443 (
            .O(N__12932),
            .I(N__12902));
    Span4Mux_h I__1442 (
            .O(N__12929),
            .I(N__12891));
    LocalMux I__1441 (
            .O(N__12926),
            .I(N__12891));
    LocalMux I__1440 (
            .O(N__12921),
            .I(N__12891));
    LocalMux I__1439 (
            .O(N__12918),
            .I(N__12891));
    LocalMux I__1438 (
            .O(N__12911),
            .I(N__12891));
    LocalMux I__1437 (
            .O(N__12908),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__1436 (
            .O(N__12905),
            .I(\this_vga_signals.vaddress_6 ));
    Odrv4 I__1435 (
            .O(N__12902),
            .I(\this_vga_signals.vaddress_6 ));
    Odrv4 I__1434 (
            .O(N__12891),
            .I(\this_vga_signals.vaddress_6 ));
    InMux I__1433 (
            .O(N__12882),
            .I(N__12876));
    InMux I__1432 (
            .O(N__12881),
            .I(N__12872));
    InMux I__1431 (
            .O(N__12880),
            .I(N__12869));
    InMux I__1430 (
            .O(N__12879),
            .I(N__12866));
    LocalMux I__1429 (
            .O(N__12876),
            .I(N__12863));
    InMux I__1428 (
            .O(N__12875),
            .I(N__12859));
    LocalMux I__1427 (
            .O(N__12872),
            .I(N__12856));
    LocalMux I__1426 (
            .O(N__12869),
            .I(N__12846));
    LocalMux I__1425 (
            .O(N__12866),
            .I(N__12841));
    Span4Mux_h I__1424 (
            .O(N__12863),
            .I(N__12841));
    InMux I__1423 (
            .O(N__12862),
            .I(N__12838));
    LocalMux I__1422 (
            .O(N__12859),
            .I(N__12833));
    Span4Mux_h I__1421 (
            .O(N__12856),
            .I(N__12833));
    InMux I__1420 (
            .O(N__12855),
            .I(N__12826));
    InMux I__1419 (
            .O(N__12854),
            .I(N__12826));
    InMux I__1418 (
            .O(N__12853),
            .I(N__12826));
    InMux I__1417 (
            .O(N__12852),
            .I(N__12823));
    InMux I__1416 (
            .O(N__12851),
            .I(N__12816));
    InMux I__1415 (
            .O(N__12850),
            .I(N__12816));
    InMux I__1414 (
            .O(N__12849),
            .I(N__12816));
    Odrv4 I__1413 (
            .O(N__12846),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__1412 (
            .O(N__12841),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1411 (
            .O(N__12838),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__1410 (
            .O(N__12833),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1409 (
            .O(N__12826),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1408 (
            .O(N__12823),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1407 (
            .O(N__12816),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    InMux I__1406 (
            .O(N__12801),
            .I(N__12798));
    LocalMux I__1405 (
            .O(N__12798),
            .I(\this_vga_signals.g2_0 ));
    InMux I__1404 (
            .O(N__12795),
            .I(N__12792));
    LocalMux I__1403 (
            .O(N__12792),
            .I(N__12789));
    Span4Mux_v I__1402 (
            .O(N__12789),
            .I(N__12786));
    Odrv4 I__1401 (
            .O(N__12786),
            .I(\this_vga_signals.g0_2_0_a2 ));
    InMux I__1400 (
            .O(N__12783),
            .I(N__12777));
    InMux I__1399 (
            .O(N__12782),
            .I(N__12777));
    LocalMux I__1398 (
            .O(N__12777),
            .I(N__12773));
    CascadeMux I__1397 (
            .O(N__12776),
            .I(N__12769));
    Span4Mux_v I__1396 (
            .O(N__12773),
            .I(N__12764));
    InMux I__1395 (
            .O(N__12772),
            .I(N__12759));
    InMux I__1394 (
            .O(N__12769),
            .I(N__12759));
    InMux I__1393 (
            .O(N__12768),
            .I(N__12754));
    InMux I__1392 (
            .O(N__12767),
            .I(N__12754));
    Odrv4 I__1391 (
            .O(N__12764),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_ns ));
    LocalMux I__1390 (
            .O(N__12759),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_ns ));
    LocalMux I__1389 (
            .O(N__12754),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_ns ));
    InMux I__1388 (
            .O(N__12747),
            .I(N__12744));
    LocalMux I__1387 (
            .O(N__12744),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3 ));
    CascadeMux I__1386 (
            .O(N__12741),
            .I(\this_vga_signals.g0_13_x0_cascade_ ));
    InMux I__1385 (
            .O(N__12738),
            .I(N__12735));
    LocalMux I__1384 (
            .O(N__12735),
            .I(\this_vga_signals.mult1_un68_sum_axb1_1 ));
    InMux I__1383 (
            .O(N__12732),
            .I(N__12729));
    LocalMux I__1382 (
            .O(N__12729),
            .I(\this_vga_signals.mult1_un47_sum_c3_1 ));
    InMux I__1381 (
            .O(N__12726),
            .I(N__12721));
    CascadeMux I__1380 (
            .O(N__12725),
            .I(N__12718));
    InMux I__1379 (
            .O(N__12724),
            .I(N__12714));
    LocalMux I__1378 (
            .O(N__12721),
            .I(N__12708));
    InMux I__1377 (
            .O(N__12718),
            .I(N__12703));
    InMux I__1376 (
            .O(N__12717),
            .I(N__12703));
    LocalMux I__1375 (
            .O(N__12714),
            .I(N__12700));
    InMux I__1374 (
            .O(N__12713),
            .I(N__12697));
    InMux I__1373 (
            .O(N__12712),
            .I(N__12694));
    InMux I__1372 (
            .O(N__12711),
            .I(N__12691));
    Odrv4 I__1371 (
            .O(N__12708),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__1370 (
            .O(N__12703),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    Odrv4 I__1369 (
            .O(N__12700),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__1368 (
            .O(N__12697),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__1367 (
            .O(N__12694),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__1366 (
            .O(N__12691),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    InMux I__1365 (
            .O(N__12678),
            .I(N__12675));
    LocalMux I__1364 (
            .O(N__12675),
            .I(N__12671));
    InMux I__1363 (
            .O(N__12674),
            .I(N__12668));
    Odrv4 I__1362 (
            .O(N__12671),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_2 ));
    LocalMux I__1361 (
            .O(N__12668),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_2 ));
    CascadeMux I__1360 (
            .O(N__12663),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_2_cascade_ ));
    InMux I__1359 (
            .O(N__12660),
            .I(N__12657));
    LocalMux I__1358 (
            .O(N__12657),
            .I(\this_vga_signals.g0_13_x1 ));
    InMux I__1357 (
            .O(N__12654),
            .I(N__12648));
    InMux I__1356 (
            .O(N__12653),
            .I(N__12642));
    InMux I__1355 (
            .O(N__12652),
            .I(N__12637));
    InMux I__1354 (
            .O(N__12651),
            .I(N__12637));
    LocalMux I__1353 (
            .O(N__12648),
            .I(N__12634));
    InMux I__1352 (
            .O(N__12647),
            .I(N__12631));
    InMux I__1351 (
            .O(N__12646),
            .I(N__12626));
    InMux I__1350 (
            .O(N__12645),
            .I(N__12626));
    LocalMux I__1349 (
            .O(N__12642),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1348 (
            .O(N__12637),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    Odrv4 I__1347 (
            .O(N__12634),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1346 (
            .O(N__12631),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1345 (
            .O(N__12626),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    InMux I__1344 (
            .O(N__12615),
            .I(N__12612));
    LocalMux I__1343 (
            .O(N__12612),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_x0 ));
    CascadeMux I__1342 (
            .O(N__12609),
            .I(\this_vga_signals.mult1_un61_sum_c3_cascade_ ));
    InMux I__1341 (
            .O(N__12606),
            .I(N__12598));
    InMux I__1340 (
            .O(N__12605),
            .I(N__12598));
    CascadeMux I__1339 (
            .O(N__12604),
            .I(N__12594));
    CascadeMux I__1338 (
            .O(N__12603),
            .I(N__12590));
    LocalMux I__1337 (
            .O(N__12598),
            .I(N__12586));
    InMux I__1336 (
            .O(N__12597),
            .I(N__12583));
    InMux I__1335 (
            .O(N__12594),
            .I(N__12572));
    InMux I__1334 (
            .O(N__12593),
            .I(N__12572));
    InMux I__1333 (
            .O(N__12590),
            .I(N__12572));
    InMux I__1332 (
            .O(N__12589),
            .I(N__12572));
    Span4Mux_h I__1331 (
            .O(N__12586),
            .I(N__12569));
    LocalMux I__1330 (
            .O(N__12583),
            .I(N__12566));
    InMux I__1329 (
            .O(N__12582),
            .I(N__12563));
    InMux I__1328 (
            .O(N__12581),
            .I(N__12560));
    LocalMux I__1327 (
            .O(N__12572),
            .I(N__12557));
    Odrv4 I__1326 (
            .O(N__12569),
            .I(\this_vga_signals.vaddress_5 ));
    Odrv4 I__1325 (
            .O(N__12566),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__1324 (
            .O(N__12563),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__1323 (
            .O(N__12560),
            .I(\this_vga_signals.vaddress_5 ));
    Odrv4 I__1322 (
            .O(N__12557),
            .I(\this_vga_signals.vaddress_5 ));
    InMux I__1321 (
            .O(N__12546),
            .I(N__12543));
    LocalMux I__1320 (
            .O(N__12543),
            .I(N__12534));
    InMux I__1319 (
            .O(N__12542),
            .I(N__12529));
    InMux I__1318 (
            .O(N__12541),
            .I(N__12529));
    InMux I__1317 (
            .O(N__12540),
            .I(N__12524));
    InMux I__1316 (
            .O(N__12539),
            .I(N__12524));
    InMux I__1315 (
            .O(N__12538),
            .I(N__12519));
    InMux I__1314 (
            .O(N__12537),
            .I(N__12519));
    Odrv4 I__1313 (
            .O(N__12534),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__1312 (
            .O(N__12529),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__1311 (
            .O(N__12524),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__1310 (
            .O(N__12519),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    CascadeMux I__1309 (
            .O(N__12510),
            .I(N__12507));
    InMux I__1308 (
            .O(N__12507),
            .I(N__12504));
    LocalMux I__1307 (
            .O(N__12504),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_x1 ));
    InMux I__1306 (
            .O(N__12501),
            .I(N__12498));
    LocalMux I__1305 (
            .O(N__12498),
            .I(\this_vga_signals.g1_2_1_0 ));
    InMux I__1304 (
            .O(N__12495),
            .I(N__12492));
    LocalMux I__1303 (
            .O(N__12492),
            .I(N__12489));
    Odrv12 I__1302 (
            .O(N__12489),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_0_0 ));
    CascadeMux I__1301 (
            .O(N__12486),
            .I(\this_vga_signals.M_vcounter_q_RNITVMCUZ0Z_3_cascade_ ));
    InMux I__1300 (
            .O(N__12483),
            .I(N__12480));
    LocalMux I__1299 (
            .O(N__12480),
            .I(\this_vga_signals.M_vcounter_q_RNIANU4QZ0Z_3 ));
    InMux I__1298 (
            .O(N__12477),
            .I(N__12474));
    LocalMux I__1297 (
            .O(N__12474),
            .I(N__12471));
    Odrv4 I__1296 (
            .O(N__12471),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0 ));
    CascadeMux I__1295 (
            .O(N__12468),
            .I(\this_vga_signals.g1_0_1_cascade_ ));
    InMux I__1294 (
            .O(N__12465),
            .I(N__12462));
    LocalMux I__1293 (
            .O(N__12462),
            .I(\this_vga_signals.g0_i_x4_0_0 ));
    InMux I__1292 (
            .O(N__12459),
            .I(N__12456));
    LocalMux I__1291 (
            .O(N__12456),
            .I(N__12453));
    Odrv4 I__1290 (
            .O(N__12453),
            .I(\this_vga_signals.g1 ));
    CascadeMux I__1289 (
            .O(N__12450),
            .I(N__12447));
    InMux I__1288 (
            .O(N__12447),
            .I(N__12444));
    LocalMux I__1287 (
            .O(N__12444),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_0_1 ));
    InMux I__1286 (
            .O(N__12441),
            .I(N__12438));
    LocalMux I__1285 (
            .O(N__12438),
            .I(N__12435));
    Span4Mux_v I__1284 (
            .O(N__12435),
            .I(N__12432));
    Odrv4 I__1283 (
            .O(N__12432),
            .I(\this_vga_signals.g0_1_0_0 ));
    CascadeMux I__1282 (
            .O(N__12429),
            .I(\this_vga_signals.g1_2_1_cascade_ ));
    InMux I__1281 (
            .O(N__12426),
            .I(N__12423));
    LocalMux I__1280 (
            .O(N__12423),
            .I(\this_vga_signals.g0_0_0_0_0 ));
    InMux I__1279 (
            .O(N__12420),
            .I(N__12417));
    LocalMux I__1278 (
            .O(N__12417),
            .I(\this_vga_signals.g0_2_0_a2_1 ));
    CascadeMux I__1277 (
            .O(N__12414),
            .I(\this_vga_signals.g0_2_0_a2_1_cascade_ ));
    InMux I__1276 (
            .O(N__12411),
            .I(N__12408));
    LocalMux I__1275 (
            .O(N__12408),
            .I(\this_vga_signals.g0_3_x1 ));
    InMux I__1274 (
            .O(N__12405),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__1273 (
            .O(N__12402),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__1272 (
            .O(N__12399),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__1271 (
            .O(N__12396),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__1270 (
            .O(N__12393),
            .I(bfn_11_24_0_));
    CEMux I__1269 (
            .O(N__12390),
            .I(N__12387));
    LocalMux I__1268 (
            .O(N__12387),
            .I(N__12384));
    Span4Mux_h I__1267 (
            .O(N__12384),
            .I(N__12381));
    Odrv4 I__1266 (
            .O(N__12381),
            .I(\this_vga_signals.N_692_1 ));
    SRMux I__1265 (
            .O(N__12378),
            .I(N__12375));
    LocalMux I__1264 (
            .O(N__12375),
            .I(N__12370));
    SRMux I__1263 (
            .O(N__12374),
            .I(N__12367));
    SRMux I__1262 (
            .O(N__12373),
            .I(N__12364));
    Span4Mux_v I__1261 (
            .O(N__12370),
            .I(N__12358));
    LocalMux I__1260 (
            .O(N__12367),
            .I(N__12358));
    LocalMux I__1259 (
            .O(N__12364),
            .I(N__12355));
    InMux I__1258 (
            .O(N__12363),
            .I(N__12352));
    Span4Mux_h I__1257 (
            .O(N__12358),
            .I(N__12349));
    Span4Mux_h I__1256 (
            .O(N__12355),
            .I(N__12344));
    LocalMux I__1255 (
            .O(N__12352),
            .I(N__12344));
    Odrv4 I__1254 (
            .O(N__12349),
            .I(\this_vga_signals.M_vcounter_q_379_0 ));
    Odrv4 I__1253 (
            .O(N__12344),
            .I(\this_vga_signals.M_vcounter_q_379_0 ));
    CascadeMux I__1252 (
            .O(N__12339),
            .I(\this_vga_signals.g0_3_x0_cascade_ ));
    InMux I__1251 (
            .O(N__12336),
            .I(N__12333));
    LocalMux I__1250 (
            .O(N__12333),
            .I(N__12330));
    Odrv4 I__1249 (
            .O(N__12330),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_0 ));
    InMux I__1248 (
            .O(N__12327),
            .I(N__12324));
    LocalMux I__1247 (
            .O(N__12324),
            .I(\this_vga_signals.M_hcounter_d7lto7_1 ));
    InMux I__1246 (
            .O(N__12321),
            .I(N__12318));
    LocalMux I__1245 (
            .O(N__12318),
            .I(\this_vga_signals.un2_hsynclto3_0 ));
    CascadeMux I__1244 (
            .O(N__12315),
            .I(\this_vga_signals.un2_hsynclto3_0_cascade_ ));
    CascadeMux I__1243 (
            .O(N__12312),
            .I(\this_vga_signals.un2_hsynclto6_0_cascade_ ));
    IoInMux I__1242 (
            .O(N__12309),
            .I(N__12306));
    LocalMux I__1241 (
            .O(N__12306),
            .I(N__12303));
    Span4Mux_s3_h I__1240 (
            .O(N__12303),
            .I(N__12300));
    Span4Mux_h I__1239 (
            .O(N__12300),
            .I(N__12297));
    Span4Mux_v I__1238 (
            .O(N__12297),
            .I(N__12294));
    Span4Mux_v I__1237 (
            .O(N__12294),
            .I(N__12291));
    Odrv4 I__1236 (
            .O(N__12291),
            .I(rgb_c_4));
    CascadeMux I__1235 (
            .O(N__12288),
            .I(N__12284));
    InMux I__1234 (
            .O(N__12287),
            .I(N__12277));
    InMux I__1233 (
            .O(N__12284),
            .I(N__12272));
    InMux I__1232 (
            .O(N__12283),
            .I(N__12272));
    InMux I__1231 (
            .O(N__12282),
            .I(N__12269));
    InMux I__1230 (
            .O(N__12281),
            .I(N__12264));
    InMux I__1229 (
            .O(N__12280),
            .I(N__12264));
    LocalMux I__1228 (
            .O(N__12277),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1227 (
            .O(N__12272),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1226 (
            .O(N__12269),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1225 (
            .O(N__12264),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    InMux I__1224 (
            .O(N__12255),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__1223 (
            .O(N__12252),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__1222 (
            .O(N__12249),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    CascadeMux I__1221 (
            .O(N__12246),
            .I(\this_vga_signals.g3_0_0_0_cascade_ ));
    InMux I__1220 (
            .O(N__12243),
            .I(N__12240));
    LocalMux I__1219 (
            .O(N__12240),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_0_0 ));
    CascadeMux I__1218 (
            .O(N__12237),
            .I(\this_vga_signals.M_hcounter_d7lt7_0_cascade_ ));
    CascadeMux I__1217 (
            .O(N__12234),
            .I(\this_vga_signals.if_m2_0_cascade_ ));
    CascadeMux I__1216 (
            .O(N__12231),
            .I(\this_vga_signals.mult1_un89_sum_c3_0_1_cascade_ ));
    CascadeMux I__1215 (
            .O(N__12228),
            .I(\this_vga_signals.haddress_1_0_cascade_ ));
    CascadeMux I__1214 (
            .O(N__12225),
            .I(N__12222));
    InMux I__1213 (
            .O(N__12222),
            .I(N__12219));
    LocalMux I__1212 (
            .O(N__12219),
            .I(N__12216));
    Span4Mux_h I__1211 (
            .O(N__12216),
            .I(N__12213));
    Span4Mux_v I__1210 (
            .O(N__12213),
            .I(N__12210));
    Odrv4 I__1209 (
            .O(N__12210),
            .I(M_this_vga_signals_address_0));
    InMux I__1208 (
            .O(N__12207),
            .I(N__12200));
    InMux I__1207 (
            .O(N__12206),
            .I(N__12197));
    InMux I__1206 (
            .O(N__12205),
            .I(N__12192));
    InMux I__1205 (
            .O(N__12204),
            .I(N__12192));
    InMux I__1204 (
            .O(N__12203),
            .I(N__12189));
    LocalMux I__1203 (
            .O(N__12200),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__1202 (
            .O(N__12197),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__1201 (
            .O(N__12192),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__1200 (
            .O(N__12189),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    InMux I__1199 (
            .O(N__12180),
            .I(N__12169));
    InMux I__1198 (
            .O(N__12179),
            .I(N__12169));
    InMux I__1197 (
            .O(N__12178),
            .I(N__12169));
    InMux I__1196 (
            .O(N__12177),
            .I(N__12160));
    InMux I__1195 (
            .O(N__12176),
            .I(N__12160));
    LocalMux I__1194 (
            .O(N__12169),
            .I(N__12157));
    InMux I__1193 (
            .O(N__12168),
            .I(N__12147));
    InMux I__1192 (
            .O(N__12167),
            .I(N__12147));
    InMux I__1191 (
            .O(N__12166),
            .I(N__12147));
    InMux I__1190 (
            .O(N__12165),
            .I(N__12147));
    LocalMux I__1189 (
            .O(N__12160),
            .I(N__12142));
    Span4Mux_h I__1188 (
            .O(N__12157),
            .I(N__12142));
    InMux I__1187 (
            .O(N__12156),
            .I(N__12139));
    LocalMux I__1186 (
            .O(N__12147),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__1185 (
            .O(N__12142),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__1184 (
            .O(N__12139),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    CascadeMux I__1183 (
            .O(N__12132),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_cascade_ ));
    CascadeMux I__1182 (
            .O(N__12129),
            .I(N__12126));
    InMux I__1181 (
            .O(N__12126),
            .I(N__12123));
    LocalMux I__1180 (
            .O(N__12123),
            .I(N__12120));
    Span4Mux_h I__1179 (
            .O(N__12120),
            .I(N__12117));
    Odrv4 I__1178 (
            .O(N__12117),
            .I(\this_vga_signals.if_m8_0_a3_1_1_6 ));
    InMux I__1177 (
            .O(N__12114),
            .I(N__12111));
    LocalMux I__1176 (
            .O(N__12111),
            .I(N__12108));
    Odrv4 I__1175 (
            .O(N__12108),
            .I(\this_vga_signals.N_5_i_0 ));
    CascadeMux I__1174 (
            .O(N__12105),
            .I(\this_vga_signals.g1_2_1_0_0_cascade_ ));
    CascadeMux I__1173 (
            .O(N__12102),
            .I(\this_vga_signals.g1_0_4_1_cascade_ ));
    InMux I__1172 (
            .O(N__12099),
            .I(N__12096));
    LocalMux I__1171 (
            .O(N__12096),
            .I(\this_vga_signals.mult1_un47_sum_c3_2_0 ));
    CascadeMux I__1170 (
            .O(N__12093),
            .I(N__12090));
    InMux I__1169 (
            .O(N__12090),
            .I(N__12087));
    LocalMux I__1168 (
            .O(N__12087),
            .I(N__12084));
    Odrv4 I__1167 (
            .O(N__12084),
            .I(\this_vga_signals.g1_0_4 ));
    CascadeMux I__1166 (
            .O(N__12081),
            .I(N__12078));
    InMux I__1165 (
            .O(N__12078),
            .I(N__12075));
    LocalMux I__1164 (
            .O(N__12075),
            .I(N__12072));
    Span4Mux_v I__1163 (
            .O(N__12072),
            .I(N__12069));
    Odrv4 I__1162 (
            .O(N__12069),
            .I(\this_vga_signals.if_m8_0_a3_1_1_4 ));
    InMux I__1161 (
            .O(N__12066),
            .I(N__12063));
    LocalMux I__1160 (
            .O(N__12063),
            .I(\this_vga_signals.g1_0 ));
    InMux I__1159 (
            .O(N__12060),
            .I(N__12057));
    LocalMux I__1158 (
            .O(N__12057),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0 ));
    CascadeMux I__1157 (
            .O(N__12054),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0_cascade_ ));
    InMux I__1156 (
            .O(N__12051),
            .I(N__12048));
    LocalMux I__1155 (
            .O(N__12048),
            .I(\this_vga_signals.g0_1_0_0_0 ));
    CascadeMux I__1154 (
            .O(N__12045),
            .I(\this_vga_signals.g2_1_0_1_cascade_ ));
    InMux I__1153 (
            .O(N__12042),
            .I(N__12034));
    InMux I__1152 (
            .O(N__12041),
            .I(N__12034));
    InMux I__1151 (
            .O(N__12040),
            .I(N__12029));
    InMux I__1150 (
            .O(N__12039),
            .I(N__12029));
    LocalMux I__1149 (
            .O(N__12034),
            .I(N__12024));
    LocalMux I__1148 (
            .O(N__12029),
            .I(N__12024));
    Odrv4 I__1147 (
            .O(N__12024),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    CascadeMux I__1146 (
            .O(N__12021),
            .I(N__12016));
    InMux I__1145 (
            .O(N__12020),
            .I(N__12012));
    InMux I__1144 (
            .O(N__12019),
            .I(N__12009));
    InMux I__1143 (
            .O(N__12016),
            .I(N__12004));
    InMux I__1142 (
            .O(N__12015),
            .I(N__12004));
    LocalMux I__1141 (
            .O(N__12012),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__1140 (
            .O(N__12009),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__1139 (
            .O(N__12004),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    CascadeMux I__1138 (
            .O(N__11997),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ));
    InMux I__1137 (
            .O(N__11994),
            .I(N__11987));
    InMux I__1136 (
            .O(N__11993),
            .I(N__11987));
    CascadeMux I__1135 (
            .O(N__11992),
            .I(N__11984));
    LocalMux I__1134 (
            .O(N__11987),
            .I(N__11979));
    InMux I__1133 (
            .O(N__11984),
            .I(N__11976));
    InMux I__1132 (
            .O(N__11983),
            .I(N__11971));
    InMux I__1131 (
            .O(N__11982),
            .I(N__11971));
    Odrv4 I__1130 (
            .O(N__11979),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__1129 (
            .O(N__11976),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__1128 (
            .O(N__11971),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    InMux I__1127 (
            .O(N__11964),
            .I(N__11961));
    LocalMux I__1126 (
            .O(N__11961),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_0 ));
    InMux I__1125 (
            .O(N__11958),
            .I(N__11947));
    InMux I__1124 (
            .O(N__11957),
            .I(N__11947));
    InMux I__1123 (
            .O(N__11956),
            .I(N__11944));
    InMux I__1122 (
            .O(N__11955),
            .I(N__11939));
    InMux I__1121 (
            .O(N__11954),
            .I(N__11939));
    InMux I__1120 (
            .O(N__11953),
            .I(N__11934));
    InMux I__1119 (
            .O(N__11952),
            .I(N__11934));
    LocalMux I__1118 (
            .O(N__11947),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1117 (
            .O(N__11944),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1116 (
            .O(N__11939),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1115 (
            .O(N__11934),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    CascadeMux I__1114 (
            .O(N__11925),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ));
    InMux I__1113 (
            .O(N__11922),
            .I(N__11919));
    LocalMux I__1112 (
            .O(N__11919),
            .I(N__11914));
    InMux I__1111 (
            .O(N__11918),
            .I(N__11911));
    InMux I__1110 (
            .O(N__11917),
            .I(N__11908));
    Odrv4 I__1109 (
            .O(N__11914),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__1108 (
            .O(N__11911),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__1107 (
            .O(N__11908),
            .I(\this_vga_signals.vaddress_c2 ));
    CascadeMux I__1106 (
            .O(N__11901),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ));
    InMux I__1105 (
            .O(N__11898),
            .I(N__11895));
    LocalMux I__1104 (
            .O(N__11895),
            .I(N__11892));
    Span4Mux_h I__1103 (
            .O(N__11892),
            .I(N__11889));
    Odrv4 I__1102 (
            .O(N__11889),
            .I(\this_vga_signals.g1_0_0_0 ));
    InMux I__1101 (
            .O(N__11886),
            .I(N__11883));
    LocalMux I__1100 (
            .O(N__11883),
            .I(N__11880));
    Odrv4 I__1099 (
            .O(N__11880),
            .I(\this_vga_signals.vaddress_2_5 ));
    CascadeMux I__1098 (
            .O(N__11877),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_x0_cascade_ ));
    InMux I__1097 (
            .O(N__11874),
            .I(N__11867));
    InMux I__1096 (
            .O(N__11873),
            .I(N__11859));
    InMux I__1095 (
            .O(N__11872),
            .I(N__11859));
    InMux I__1094 (
            .O(N__11871),
            .I(N__11859));
    InMux I__1093 (
            .O(N__11870),
            .I(N__11856));
    LocalMux I__1092 (
            .O(N__11867),
            .I(N__11853));
    InMux I__1091 (
            .O(N__11866),
            .I(N__11850));
    LocalMux I__1090 (
            .O(N__11859),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__1089 (
            .O(N__11856),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__1088 (
            .O(N__11853),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__1087 (
            .O(N__11850),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    InMux I__1086 (
            .O(N__11841),
            .I(N__11837));
    InMux I__1085 (
            .O(N__11840),
            .I(N__11834));
    LocalMux I__1084 (
            .O(N__11837),
            .I(N__11831));
    LocalMux I__1083 (
            .O(N__11834),
            .I(N__11828));
    Odrv4 I__1082 (
            .O(N__11831),
            .I(\this_vga_signals.if_m8_0_a3_1_1_1 ));
    Odrv4 I__1081 (
            .O(N__11828),
            .I(\this_vga_signals.if_m8_0_a3_1_1_1 ));
    CascadeMux I__1080 (
            .O(N__11823),
            .I(\this_vga_signals.if_N_5_cascade_ ));
    InMux I__1079 (
            .O(N__11820),
            .I(N__11817));
    LocalMux I__1078 (
            .O(N__11817),
            .I(N__11814));
    Odrv4 I__1077 (
            .O(N__11814),
            .I(\this_vga_signals.if_m8_0_a3_1_1_0 ));
    CascadeMux I__1076 (
            .O(N__11811),
            .I(\this_vga_signals.N_5_i_0_cascade_ ));
    InMux I__1075 (
            .O(N__11808),
            .I(N__11805));
    LocalMux I__1074 (
            .O(N__11805),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    InMux I__1073 (
            .O(N__11802),
            .I(N__11797));
    InMux I__1072 (
            .O(N__11801),
            .I(N__11792));
    InMux I__1071 (
            .O(N__11800),
            .I(N__11792));
    LocalMux I__1070 (
            .O(N__11797),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__1069 (
            .O(N__11792),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    InMux I__1068 (
            .O(N__11787),
            .I(N__11782));
    InMux I__1067 (
            .O(N__11786),
            .I(N__11777));
    InMux I__1066 (
            .O(N__11785),
            .I(N__11777));
    LocalMux I__1065 (
            .O(N__11782),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__1064 (
            .O(N__11777),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    InMux I__1063 (
            .O(N__11772),
            .I(N__11769));
    LocalMux I__1062 (
            .O(N__11769),
            .I(N__11766));
    Span4Mux_h I__1061 (
            .O(N__11766),
            .I(N__11763));
    Odrv4 I__1060 (
            .O(N__11763),
            .I(\this_vga_signals.SUM_3_1_tz ));
    IoInMux I__1059 (
            .O(N__11760),
            .I(N__11757));
    LocalMux I__1058 (
            .O(N__11757),
            .I(N__11754));
    IoSpan4Mux I__1057 (
            .O(N__11754),
            .I(N__11751));
    IoSpan4Mux I__1056 (
            .O(N__11751),
            .I(N__11748));
    Span4Mux_s1_v I__1055 (
            .O(N__11748),
            .I(N__11745));
    Span4Mux_v I__1054 (
            .O(N__11745),
            .I(N__11742));
    Odrv4 I__1053 (
            .O(N__11742),
            .I(this_vga_signals_hvisibility_i));
    SRMux I__1052 (
            .O(N__11739),
            .I(N__11736));
    LocalMux I__1051 (
            .O(N__11736),
            .I(N__11732));
    SRMux I__1050 (
            .O(N__11735),
            .I(N__11729));
    Span4Mux_h I__1049 (
            .O(N__11732),
            .I(N__11726));
    LocalMux I__1048 (
            .O(N__11729),
            .I(N__11723));
    Odrv4 I__1047 (
            .O(N__11726),
            .I(M_stage_q_RNIC68K4_9));
    Odrv12 I__1046 (
            .O(N__11723),
            .I(M_stage_q_RNIC68K4_9));
    CascadeMux I__1045 (
            .O(N__11718),
            .I(N__11715));
    InMux I__1044 (
            .O(N__11715),
            .I(N__11712));
    LocalMux I__1043 (
            .O(N__11712),
            .I(N__11708));
    InMux I__1042 (
            .O(N__11711),
            .I(N__11705));
    Span4Mux_h I__1041 (
            .O(N__11708),
            .I(N__11702));
    LocalMux I__1040 (
            .O(N__11705),
            .I(\this_vga_signals.vaddress_3_5 ));
    Odrv4 I__1039 (
            .O(N__11702),
            .I(\this_vga_signals.vaddress_3_5 ));
    CascadeMux I__1038 (
            .O(N__11697),
            .I(\this_vga_signals.if_m8_0_a3_1_1_5_cascade_ ));
    InMux I__1037 (
            .O(N__11694),
            .I(N__11691));
    LocalMux I__1036 (
            .O(N__11691),
            .I(N__11688));
    Span4Mux_v I__1035 (
            .O(N__11688),
            .I(N__11685));
    Odrv4 I__1034 (
            .O(N__11685),
            .I(\this_vga_signals.g0_6_0_0 ));
    CascadeMux I__1033 (
            .O(N__11682),
            .I(\this_vga_signals.un6_vvisibilitylt8_cascade_ ));
    CascadeMux I__1032 (
            .O(N__11679),
            .I(N__11676));
    InMux I__1031 (
            .O(N__11676),
            .I(N__11673));
    LocalMux I__1030 (
            .O(N__11673),
            .I(\this_vga_signals.vvisibility_1 ));
    InMux I__1029 (
            .O(N__11670),
            .I(N__11667));
    LocalMux I__1028 (
            .O(N__11667),
            .I(\this_vga_signals.vaddress_0_5 ));
    CascadeMux I__1027 (
            .O(N__11664),
            .I(\this_vga_signals.if_m8_0_a3_1_1_3_cascade_ ));
    CascadeMux I__1026 (
            .O(N__11661),
            .I(\this_vga_signals.g0_6_0_cascade_ ));
    InMux I__1025 (
            .O(N__11658),
            .I(N__11655));
    LocalMux I__1024 (
            .O(N__11655),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d ));
    InMux I__1023 (
            .O(N__11652),
            .I(N__11649));
    LocalMux I__1022 (
            .O(N__11649),
            .I(N__11646));
    Odrv4 I__1021 (
            .O(N__11646),
            .I(\this_vga_signals.i6_mux_0 ));
    CascadeMux I__1020 (
            .O(N__11643),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_0_cascade_ ));
    InMux I__1019 (
            .O(N__11640),
            .I(N__11637));
    LocalMux I__1018 (
            .O(N__11637),
            .I(\this_vga_signals.g0_i_x4_0_a2_1 ));
    InMux I__1017 (
            .O(N__11634),
            .I(N__11631));
    LocalMux I__1016 (
            .O(N__11631),
            .I(N__11628));
    Span4Mux_v I__1015 (
            .O(N__11628),
            .I(N__11625));
    Odrv4 I__1014 (
            .O(N__11625),
            .I(\this_vga_signals.if_m8_0_a3_1_1_2 ));
    CascadeMux I__1013 (
            .O(N__11622),
            .I(\this_vga_signals.vaddress_1_0_5_cascade_ ));
    CascadeMux I__1012 (
            .O(N__11619),
            .I(\this_vga_signals.SUM_2_i_1_1_3_cascade_ ));
    CascadeMux I__1011 (
            .O(N__11616),
            .I(N__11613));
    InMux I__1010 (
            .O(N__11613),
            .I(N__11610));
    LocalMux I__1009 (
            .O(N__11610),
            .I(\this_vga_signals.SUM_2_i_1_1_1_3 ));
    InMux I__1008 (
            .O(N__11607),
            .I(N__11604));
    LocalMux I__1007 (
            .O(N__11604),
            .I(N__11601));
    Odrv4 I__1006 (
            .O(N__11601),
            .I(\this_vga_signals.N_1_3_1 ));
    CascadeMux I__1005 (
            .O(N__11598),
            .I(\this_vga_signals.N_1_3_1_cascade_ ));
    InMux I__1004 (
            .O(N__11595),
            .I(N__11592));
    LocalMux I__1003 (
            .O(N__11592),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    CascadeMux I__1002 (
            .O(N__11589),
            .I(N__11586));
    CascadeBuf I__1001 (
            .O(N__11586),
            .I(N__11583));
    CascadeMux I__1000 (
            .O(N__11583),
            .I(N__11580));
    InMux I__999 (
            .O(N__11580),
            .I(N__11577));
    LocalMux I__998 (
            .O(N__11577),
            .I(N__11573));
    InMux I__997 (
            .O(N__11576),
            .I(N__11570));
    Span4Mux_v I__996 (
            .O(N__11573),
            .I(N__11567));
    LocalMux I__995 (
            .O(N__11570),
            .I(M_this_map_address_qZ0Z_6));
    Odrv4 I__994 (
            .O(N__11567),
            .I(M_this_map_address_qZ0Z_6));
    InMux I__993 (
            .O(N__11562),
            .I(un1_M_this_map_address_q_cry_5));
    CascadeMux I__992 (
            .O(N__11559),
            .I(N__11556));
    CascadeBuf I__991 (
            .O(N__11556),
            .I(N__11553));
    CascadeMux I__990 (
            .O(N__11553),
            .I(N__11550));
    InMux I__989 (
            .O(N__11550),
            .I(N__11547));
    LocalMux I__988 (
            .O(N__11547),
            .I(N__11543));
    InMux I__987 (
            .O(N__11546),
            .I(N__11540));
    Span4Mux_v I__986 (
            .O(N__11543),
            .I(N__11537));
    LocalMux I__985 (
            .O(N__11540),
            .I(M_this_map_address_qZ0Z_7));
    Odrv4 I__984 (
            .O(N__11537),
            .I(M_this_map_address_qZ0Z_7));
    InMux I__983 (
            .O(N__11532),
            .I(un1_M_this_map_address_q_cry_6));
    CascadeMux I__982 (
            .O(N__11529),
            .I(N__11526));
    CascadeBuf I__981 (
            .O(N__11526),
            .I(N__11523));
    CascadeMux I__980 (
            .O(N__11523),
            .I(N__11520));
    InMux I__979 (
            .O(N__11520),
            .I(N__11517));
    LocalMux I__978 (
            .O(N__11517),
            .I(N__11513));
    InMux I__977 (
            .O(N__11516),
            .I(N__11510));
    Span4Mux_v I__976 (
            .O(N__11513),
            .I(N__11507));
    LocalMux I__975 (
            .O(N__11510),
            .I(M_this_map_address_qZ0Z_8));
    Odrv4 I__974 (
            .O(N__11507),
            .I(M_this_map_address_qZ0Z_8));
    InMux I__973 (
            .O(N__11502),
            .I(bfn_9_24_0_));
    InMux I__972 (
            .O(N__11499),
            .I(un1_M_this_map_address_q_cry_8));
    CascadeMux I__971 (
            .O(N__11496),
            .I(N__11493));
    CascadeBuf I__970 (
            .O(N__11493),
            .I(N__11490));
    CascadeMux I__969 (
            .O(N__11490),
            .I(N__11487));
    InMux I__968 (
            .O(N__11487),
            .I(N__11484));
    LocalMux I__967 (
            .O(N__11484),
            .I(N__11480));
    InMux I__966 (
            .O(N__11483),
            .I(N__11477));
    Span4Mux_v I__965 (
            .O(N__11480),
            .I(N__11474));
    LocalMux I__964 (
            .O(N__11477),
            .I(M_this_map_address_qZ0Z_9));
    Odrv4 I__963 (
            .O(N__11474),
            .I(M_this_map_address_qZ0Z_9));
    InMux I__962 (
            .O(N__11469),
            .I(N__11466));
    LocalMux I__961 (
            .O(N__11466),
            .I(N_89_0));
    InMux I__960 (
            .O(N__11463),
            .I(N__11460));
    LocalMux I__959 (
            .O(N__11460),
            .I(N_83_0));
    InMux I__958 (
            .O(N__11457),
            .I(N__11454));
    LocalMux I__957 (
            .O(N__11454),
            .I(N__11451));
    Odrv4 I__956 (
            .O(N__11451),
            .I(N_85_0));
    CascadeMux I__955 (
            .O(N__11448),
            .I(\this_vga_signals.vaddress_3_0_5_cascade_ ));
    InMux I__954 (
            .O(N__11445),
            .I(N__11442));
    LocalMux I__953 (
            .O(N__11442),
            .I(N__11439));
    Span4Mux_h I__952 (
            .O(N__11439),
            .I(N__11436));
    Odrv4 I__951 (
            .O(N__11436),
            .I(\this_vga_signals.g0_6_0_0_0 ));
    InMux I__950 (
            .O(N__11433),
            .I(N__11430));
    LocalMux I__949 (
            .O(N__11430),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    InMux I__948 (
            .O(N__11427),
            .I(N__11424));
    LocalMux I__947 (
            .O(N__11424),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    InMux I__946 (
            .O(N__11421),
            .I(N__11418));
    LocalMux I__945 (
            .O(N__11418),
            .I(\this_vga_signals.g0_0_0 ));
    CascadeMux I__944 (
            .O(N__11415),
            .I(N__11412));
    CascadeBuf I__943 (
            .O(N__11412),
            .I(N__11409));
    CascadeMux I__942 (
            .O(N__11409),
            .I(N__11406));
    InMux I__941 (
            .O(N__11406),
            .I(N__11403));
    LocalMux I__940 (
            .O(N__11403),
            .I(N__11399));
    InMux I__939 (
            .O(N__11402),
            .I(N__11396));
    Sp12to4 I__938 (
            .O(N__11399),
            .I(N__11393));
    LocalMux I__937 (
            .O(N__11396),
            .I(M_this_map_address_qZ0Z_0));
    Odrv12 I__936 (
            .O(N__11393),
            .I(M_this_map_address_qZ0Z_0));
    CascadeMux I__935 (
            .O(N__11388),
            .I(N__11385));
    CascadeBuf I__934 (
            .O(N__11385),
            .I(N__11382));
    CascadeMux I__933 (
            .O(N__11382),
            .I(N__11379));
    InMux I__932 (
            .O(N__11379),
            .I(N__11376));
    LocalMux I__931 (
            .O(N__11376),
            .I(N__11372));
    InMux I__930 (
            .O(N__11375),
            .I(N__11369));
    Span4Mux_v I__929 (
            .O(N__11372),
            .I(N__11366));
    LocalMux I__928 (
            .O(N__11369),
            .I(M_this_map_address_qZ0Z_1));
    Odrv4 I__927 (
            .O(N__11366),
            .I(M_this_map_address_qZ0Z_1));
    InMux I__926 (
            .O(N__11361),
            .I(un1_M_this_map_address_q_cry_0));
    CascadeMux I__925 (
            .O(N__11358),
            .I(N__11355));
    CascadeBuf I__924 (
            .O(N__11355),
            .I(N__11352));
    CascadeMux I__923 (
            .O(N__11352),
            .I(N__11349));
    InMux I__922 (
            .O(N__11349),
            .I(N__11346));
    LocalMux I__921 (
            .O(N__11346),
            .I(N__11342));
    InMux I__920 (
            .O(N__11345),
            .I(N__11339));
    Span4Mux_v I__919 (
            .O(N__11342),
            .I(N__11336));
    LocalMux I__918 (
            .O(N__11339),
            .I(M_this_map_address_qZ0Z_2));
    Odrv4 I__917 (
            .O(N__11336),
            .I(M_this_map_address_qZ0Z_2));
    InMux I__916 (
            .O(N__11331),
            .I(un1_M_this_map_address_q_cry_1));
    CascadeMux I__915 (
            .O(N__11328),
            .I(N__11325));
    CascadeBuf I__914 (
            .O(N__11325),
            .I(N__11322));
    CascadeMux I__913 (
            .O(N__11322),
            .I(N__11319));
    InMux I__912 (
            .O(N__11319),
            .I(N__11316));
    LocalMux I__911 (
            .O(N__11316),
            .I(N__11312));
    InMux I__910 (
            .O(N__11315),
            .I(N__11309));
    Span4Mux_v I__909 (
            .O(N__11312),
            .I(N__11306));
    LocalMux I__908 (
            .O(N__11309),
            .I(M_this_map_address_qZ0Z_3));
    Odrv4 I__907 (
            .O(N__11306),
            .I(M_this_map_address_qZ0Z_3));
    InMux I__906 (
            .O(N__11301),
            .I(un1_M_this_map_address_q_cry_2));
    CascadeMux I__905 (
            .O(N__11298),
            .I(N__11295));
    CascadeBuf I__904 (
            .O(N__11295),
            .I(N__11292));
    CascadeMux I__903 (
            .O(N__11292),
            .I(N__11289));
    InMux I__902 (
            .O(N__11289),
            .I(N__11286));
    LocalMux I__901 (
            .O(N__11286),
            .I(N__11282));
    InMux I__900 (
            .O(N__11285),
            .I(N__11279));
    Span4Mux_v I__899 (
            .O(N__11282),
            .I(N__11276));
    LocalMux I__898 (
            .O(N__11279),
            .I(M_this_map_address_qZ0Z_4));
    Odrv4 I__897 (
            .O(N__11276),
            .I(M_this_map_address_qZ0Z_4));
    InMux I__896 (
            .O(N__11271),
            .I(un1_M_this_map_address_q_cry_3));
    CascadeMux I__895 (
            .O(N__11268),
            .I(N__11265));
    CascadeBuf I__894 (
            .O(N__11265),
            .I(N__11262));
    CascadeMux I__893 (
            .O(N__11262),
            .I(N__11259));
    InMux I__892 (
            .O(N__11259),
            .I(N__11256));
    LocalMux I__891 (
            .O(N__11256),
            .I(N__11252));
    InMux I__890 (
            .O(N__11255),
            .I(N__11249));
    Span4Mux_v I__889 (
            .O(N__11252),
            .I(N__11246));
    LocalMux I__888 (
            .O(N__11249),
            .I(M_this_map_address_qZ0Z_5));
    Odrv4 I__887 (
            .O(N__11246),
            .I(M_this_map_address_qZ0Z_5));
    InMux I__886 (
            .O(N__11241),
            .I(un1_M_this_map_address_q_cry_4));
    CascadeMux I__885 (
            .O(N__11238),
            .I(\this_vga_signals.vsync_1_3_cascade_ ));
    IoInMux I__884 (
            .O(N__11235),
            .I(N__11232));
    LocalMux I__883 (
            .O(N__11232),
            .I(N__11229));
    IoSpan4Mux I__882 (
            .O(N__11229),
            .I(N__11226));
    Sp12to4 I__881 (
            .O(N__11226),
            .I(N__11223));
    Span12Mux_v I__880 (
            .O(N__11223),
            .I(N__11220));
    Odrv12 I__879 (
            .O(N__11220),
            .I(this_vga_signals_vsync_1_i));
    CascadeMux I__878 (
            .O(N__11217),
            .I(\this_vga_signals.g0_2_0_cascade_ ));
    CascadeMux I__877 (
            .O(N__11214),
            .I(\this_vga_signals.N_43_1_cascade_ ));
    InMux I__876 (
            .O(N__11211),
            .I(N__11208));
    LocalMux I__875 (
            .O(N__11208),
            .I(\this_vga_signals.un2_vsynclt8 ));
    InMux I__874 (
            .O(N__11205),
            .I(N__11202));
    LocalMux I__873 (
            .O(N__11202),
            .I(\this_vga_signals.vsync_1_2 ));
    InMux I__872 (
            .O(N__11199),
            .I(N__11196));
    LocalMux I__871 (
            .O(N__11196),
            .I(\this_vga_signals.g1_1 ));
    InMux I__870 (
            .O(N__11193),
            .I(N__11190));
    LocalMux I__869 (
            .O(N__11190),
            .I(N__11187));
    Span12Mux_h I__868 (
            .O(N__11187),
            .I(N__11184));
    Odrv12 I__867 (
            .O(N__11184),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    CascadeMux I__866 (
            .O(N__11181),
            .I(\this_vga_signals.g0_0_0_0_cascade_ ));
    CascadeMux I__865 (
            .O(N__11178),
            .I(\this_vga_signals.g1_1_1_cascade_ ));
    InMux I__864 (
            .O(N__11175),
            .I(N__11172));
    LocalMux I__863 (
            .O(N__11172),
            .I(N__11169));
    Odrv4 I__862 (
            .O(N__11169),
            .I(\this_vga_signals.g1_1_0 ));
    InMux I__861 (
            .O(N__11166),
            .I(N__11163));
    LocalMux I__860 (
            .O(N__11163),
            .I(\this_vga_signals.N_4_0_0 ));
    CascadeMux I__859 (
            .O(N__11160),
            .I(\this_vga_signals.mult1_un47_sum_c3_0_cascade_ ));
    InMux I__858 (
            .O(N__11157),
            .I(N__11154));
    LocalMux I__857 (
            .O(N__11154),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_1 ));
    CascadeMux I__856 (
            .O(N__11151),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_d_1_cascade_ ));
    CascadeMux I__855 (
            .O(N__11148),
            .I(\this_vga_signals.g2_1_cascade_ ));
    InMux I__854 (
            .O(N__11145),
            .I(N__11142));
    LocalMux I__853 (
            .O(N__11142),
            .I(\this_vga_signals.g2 ));
    IoInMux I__852 (
            .O(N__11139),
            .I(N__11136));
    LocalMux I__851 (
            .O(N__11136),
            .I(N__11133));
    Span12Mux_s8_h I__850 (
            .O(N__11133),
            .I(N__11130));
    Span12Mux_v I__849 (
            .O(N__11130),
            .I(N__11127));
    Odrv12 I__848 (
            .O(N__11127),
            .I(rgb_c_0));
    IoInMux I__847 (
            .O(N__11124),
            .I(N__11121));
    LocalMux I__846 (
            .O(N__11121),
            .I(N__11118));
    Odrv12 I__845 (
            .O(N__11118),
            .I(rgb_c_1));
    CascadeMux I__844 (
            .O(N__11115),
            .I(N__11112));
    InMux I__843 (
            .O(N__11112),
            .I(N__11109));
    LocalMux I__842 (
            .O(N__11109),
            .I(M_this_vga_signals_address_2));
    CascadeMux I__841 (
            .O(N__11106),
            .I(N__11103));
    InMux I__840 (
            .O(N__11103),
            .I(N__11100));
    LocalMux I__839 (
            .O(N__11100),
            .I(N__11097));
    Odrv4 I__838 (
            .O(N__11097),
            .I(M_this_vga_signals_address_6));
    CascadeMux I__837 (
            .O(N__11094),
            .I(N__11091));
    InMux I__836 (
            .O(N__11091),
            .I(N__11088));
    LocalMux I__835 (
            .O(N__11088),
            .I(M_this_vga_signals_address_4));
    CascadeMux I__834 (
            .O(N__11085),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_ ));
    CascadeMux I__833 (
            .O(N__11082),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_0_cascade_ ));
    CascadeMux I__832 (
            .O(N__11079),
            .I(N__11076));
    InMux I__831 (
            .O(N__11076),
            .I(N__11073));
    LocalMux I__830 (
            .O(N__11073),
            .I(M_this_vga_signals_address_7));
    IoInMux I__829 (
            .O(N__11070),
            .I(N__11067));
    LocalMux I__828 (
            .O(N__11067),
            .I(\this_vga_signals.N_692_0 ));
    InMux I__827 (
            .O(N__11064),
            .I(N__11061));
    LocalMux I__826 (
            .O(N__11061),
            .I(port_clk_c));
    IoInMux I__825 (
            .O(N__11058),
            .I(N__11055));
    LocalMux I__824 (
            .O(N__11055),
            .I(port_data_rw_0_i));
    IoInMux I__823 (
            .O(N__11052),
            .I(N__11049));
    LocalMux I__822 (
            .O(N__11049),
            .I(N__11046));
    Span4Mux_s2_h I__821 (
            .O(N__11046),
            .I(N__11043));
    Span4Mux_v I__820 (
            .O(N__11043),
            .I(N__11040));
    Odrv4 I__819 (
            .O(N__11040),
            .I(port_nmib_0_i));
    IoInMux I__818 (
            .O(N__11037),
            .I(N__11034));
    LocalMux I__817 (
            .O(N__11034),
            .I(N__11031));
    Span12Mux_s2_v I__816 (
            .O(N__11031),
            .I(N__11028));
    Odrv12 I__815 (
            .O(N__11028),
            .I(this_vga_signals_vvisibility_i));
    defparam IN_MUX_bfv_24_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_22_0_));
    defparam IN_MUX_bfv_24_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_23_0_ (
            .carryinitin(un1_M_this_external_address_q_cry_7),
            .carryinitout(bfn_24_23_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_11_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_24_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_11_24_0_));
    defparam IN_MUX_bfv_23_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_19_0_));
    defparam IN_MUX_bfv_23_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_20_0_ (
            .carryinitin(\this_ppu.un1_M_vaddress_q_cry_7 ),
            .carryinitout(bfn_23_20_0_));
    defparam IN_MUX_bfv_22_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_19_0_));
    defparam IN_MUX_bfv_22_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_20_0_ (
            .carryinitin(\this_ppu.un1_M_haddress_q_cry_7 ),
            .carryinitout(bfn_22_20_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(M_this_data_count_q_cry_7),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_23_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_16_0_));
    defparam IN_MUX_bfv_21_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_16_0_));
    defparam IN_MUX_bfv_22_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_17_0_));
    defparam IN_MUX_bfv_22_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_18_0_ (
            .carryinitin(\this_ppu.un1_M_vaddress_q_3_cry_7 ),
            .carryinitout(bfn_22_18_0_));
    defparam IN_MUX_bfv_21_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_18_0_));
    defparam IN_MUX_bfv_21_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_19_0_ (
            .carryinitin(\this_ppu.un1_M_haddress_q_2_cry_7 ),
            .carryinitout(bfn_21_19_0_));
    defparam IN_MUX_bfv_19_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_22_0_));
    defparam IN_MUX_bfv_19_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_23_0_ (
            .carryinitin(un1_M_this_sprites_address_q_cry_7),
            .carryinitout(bfn_19_23_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(un1_M_this_map_address_q_cry_7),
            .carryinitout(bfn_9_24_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNIR1G77_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__11070),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_692_0_g ));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNI67JU6_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__16293),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_988_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_9  (
            .USERSIGNALTOGLOBALBUFFER(N__22858),
            .GLOBALBUFFEROUTPUT(M_this_reset_cond_out_g_0));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_1_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_1_17_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__19056),
            .in2(_gnd_net_),
            .in3(N__14736),
            .lcout(\this_vga_signals.N_692_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_1_21_2 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_1_21_2 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_1_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_1_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11064),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34592),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.port_data_rw_0_i_LC_1_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.port_data_rw_0_i_LC_1_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.port_data_rw_0_i_LC_1_21_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \this_vga_signals.port_data_rw_0_i_LC_1_21_5  (
            .in0(N__21710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22923),
            .lcout(port_data_rw_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKCDU5_9_LC_3_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKCDU5_9_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKCDU5_9_LC_3_16_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIKCDU5_9_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(N__22931),
            .in2(_gnd_net_),
            .in3(N__22989),
            .lcout(port_nmib_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_0_9_LC_5_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_0_9_LC_5_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_0_9_LC_5_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_0_9_LC_5_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22978),
            .lcout(this_vga_signals_vvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_6_18_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_6_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_6_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_6_18_5  (
            .in0(_gnd_net_),
            .in1(N__15818),
            .in2(_gnd_net_),
            .in3(N__14898),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_6_18_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_6_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_6_18_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_6_18_7  (
            .in0(N__15663),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15819),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGJMLD1_9_LC_7_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGJMLD1_9_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGJMLD1_9_LC_7_18_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIGJMLD1_9_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(N__15590),
            .in2(_gnd_net_),
            .in3(N__13131),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_7_18_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_7_18_6 .LUT_INIT=16'b0001010100111101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_7_18_6  (
            .in0(N__18858),
            .in1(N__18813),
            .in2(N__18759),
            .in3(N__18702),
            .lcout(\this_vga_ramdac.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNILR5N4_8_LC_9_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNILR5N4_8_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNILR5N4_8_LC_9_17_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNILR5N4_8_LC_9_17_1  (
            .in0(N__11772),
            .in1(N__15587),
            .in2(_gnd_net_),
            .in3(N__14691),
            .lcout(M_this_vga_signals_address_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI9V9QB_9_LC_9_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI9V9QB_9_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI9V9QB_9_LC_9_17_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI9V9QB_9_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__15588),
            .in2(_gnd_net_),
            .in3(N__13476),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_LC_9_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_LC_9_17_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_LC_9_17_5  (
            .in0(N__12795),
            .in1(N__12477),
            .in2(N__15403),
            .in3(N__12336),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_9_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_9_17_6 .LUT_INIT=16'b0101110011000101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_m2_LC_9_17_6  (
            .in0(N__15485),
            .in1(N__12459),
            .in2(N__11085),
            .in3(N__12981),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIOIKI4Q_1_LC_9_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIOIKI4Q_1_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIOIKI4Q_1_LC_9_17_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIOIKI4Q_1_LC_9_17_7  (
            .in0(N__15589),
            .in1(N__11175),
            .in2(N__11082),
            .in3(N__11898),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_9_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_9_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14205),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34541),
            .ce(N__14762),
            .sr(N__14732));
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_9_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_9_19_0 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_0_LC_9_19_0  (
            .in0(N__11445),
            .in1(N__11157),
            .in2(_gnd_net_),
            .in3(N__13387),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_9_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_9_19_1 .LUT_INIT=16'b1101100010001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_2_LC_9_19_1  (
            .in0(N__11166),
            .in1(N__11145),
            .in2(N__11181),
            .in3(N__13299),
            .lcout(),
            .ltout(\this_vga_signals.g1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIO70OS4_1_LC_9_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIO70OS4_1_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIO70OS4_1_LC_9_19_2 .LUT_INIT=16'b0100110111010100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIO70OS4_1_LC_9_19_2  (
            .in0(N__15481),
            .in1(N__15392),
            .in2(N__11178),
            .in3(N__11640),
            .lcout(\this_vga_signals.g1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_0_a2_LC_9_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_a2_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_a2_LC_9_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_0_a2_LC_9_19_3  (
            .in0(N__13386),
            .in1(N__16483),
            .in2(N__15306),
            .in3(N__13297),
            .lcout(\this_vga_signals.N_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_9_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_9_19_4 .LUT_INIT=16'b1001000111011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_19_LC_9_19_4  (
            .in0(N__12967),
            .in1(N__12206),
            .in2(N__11718),
            .in3(N__12881),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_9_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_9_19_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_12_LC_9_19_5  (
            .in0(N__16703),
            .in1(N__16482),
            .in2(N__11160),
            .in3(N__12724),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_3_d_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_3_d_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_9_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_9_19_6 .LUT_INIT=16'b0000101011110101;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_1_LC_9_19_6  (
            .in0(N__11694),
            .in1(_gnd_net_),
            .in2(N__11151),
            .in3(N__13385),
            .lcout(),
            .ltout(\this_vga_signals.g2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_LC_9_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_LC_9_19_7 .LUT_INIT=16'b1101010001001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_LC_9_19_7  (
            .in0(N__15391),
            .in1(N__15295),
            .in2(N__11148),
            .in3(N__13298),
            .lcout(\this_vga_signals.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_9_LC_9_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_9_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_9_LC_9_20_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_9_LC_9_20_0  (
            .in0(N__17172),
            .in1(N__20108),
            .in2(N__16779),
            .in3(N__16475),
            .lcout(),
            .ltout(\this_vga_signals.vsync_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_9_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_9_20_1 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_9_20_1  (
            .in0(N__11211),
            .in1(N__11205),
            .in2(N__11238),
            .in3(N__16601),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_LC_9_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_LC_9_20_2 .LUT_INIT=16'b1110101000010101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_LC_9_20_2  (
            .in0(N__16600),
            .in1(N__16473),
            .in2(N__16778),
            .in3(N__17066),
            .lcout(),
            .ltout(\this_vga_signals.g0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_9_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_9_20_3 .LUT_INIT=16'b0010110111110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_LC_9_20_3  (
            .in0(N__11607),
            .in1(N__11421),
            .in2(N__11217),
            .in3(N__13025),
            .lcout(),
            .ltout(\this_vga_signals.N_43_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_9_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_9_20_4 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_LC_9_20_4  (
            .in0(N__16771),
            .in1(N__11199),
            .in2(N__11214),
            .in3(N__12969),
            .lcout(\this_vga_signals.i6_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_9_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_9_20_5 .LUT_INIT=16'b0000000101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_9_20_5  (
            .in0(N__16474),
            .in1(N__15394),
            .in2(N__15486),
            .in3(N__15296),
            .lcout(\this_vga_signals.un2_vsynclt8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNICSHP_2_LC_9_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNICSHP_2_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNICSHP_2_LC_9_20_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNICSHP_2_LC_9_20_6  (
            .in0(N__15395),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17067),
            .lcout(\this_vga_signals.vsync_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_LC_9_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_LC_9_20_7 .LUT_INIT=16'b0001101110001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_LC_9_20_7  (
            .in0(N__12968),
            .in1(N__16767),
            .in2(N__16490),
            .in3(N__12882),
            .lcout(\this_vga_signals.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_9_21_1 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_9_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11427),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34566),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_9_21_4 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_9_21_4 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_9_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11193),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34566),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_9_21_6 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_9_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11433),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34566),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIP5821_9_LC_9_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIP5821_9_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIP5821_9_LC_9_21_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIP5821_9_LC_9_21_7  (
            .in0(N__20103),
            .in1(N__17167),
            .in2(_gnd_net_),
            .in3(N__16609),
            .lcout(\this_vga_signals.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_0_LC_9_23_0.C_ON=1'b1;
    defparam M_this_map_address_q_0_LC_9_23_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_0_LC_9_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_0_LC_9_23_0 (
            .in0(_gnd_net_),
            .in1(N__11402),
            .in2(N__18260),
            .in3(N__18255),
            .lcout(M_this_map_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(un1_M_this_map_address_q_cry_0),
            .clk(N__34575),
            .ce(),
            .sr(N__11739));
    defparam M_this_map_address_q_1_LC_9_23_1.C_ON=1'b1;
    defparam M_this_map_address_q_1_LC_9_23_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_1_LC_9_23_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_1_LC_9_23_1 (
            .in0(_gnd_net_),
            .in1(N__11375),
            .in2(_gnd_net_),
            .in3(N__11361),
            .lcout(M_this_map_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_0),
            .carryout(un1_M_this_map_address_q_cry_1),
            .clk(N__34575),
            .ce(),
            .sr(N__11739));
    defparam M_this_map_address_q_2_LC_9_23_2.C_ON=1'b1;
    defparam M_this_map_address_q_2_LC_9_23_2.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_2_LC_9_23_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_2_LC_9_23_2 (
            .in0(_gnd_net_),
            .in1(N__11345),
            .in2(_gnd_net_),
            .in3(N__11331),
            .lcout(M_this_map_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_1),
            .carryout(un1_M_this_map_address_q_cry_2),
            .clk(N__34575),
            .ce(),
            .sr(N__11739));
    defparam M_this_map_address_q_3_LC_9_23_3.C_ON=1'b1;
    defparam M_this_map_address_q_3_LC_9_23_3.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_3_LC_9_23_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_3_LC_9_23_3 (
            .in0(_gnd_net_),
            .in1(N__11315),
            .in2(_gnd_net_),
            .in3(N__11301),
            .lcout(M_this_map_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_2),
            .carryout(un1_M_this_map_address_q_cry_3),
            .clk(N__34575),
            .ce(),
            .sr(N__11739));
    defparam M_this_map_address_q_4_LC_9_23_4.C_ON=1'b1;
    defparam M_this_map_address_q_4_LC_9_23_4.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_4_LC_9_23_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_4_LC_9_23_4 (
            .in0(_gnd_net_),
            .in1(N__11285),
            .in2(_gnd_net_),
            .in3(N__11271),
            .lcout(M_this_map_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_3),
            .carryout(un1_M_this_map_address_q_cry_4),
            .clk(N__34575),
            .ce(),
            .sr(N__11739));
    defparam M_this_map_address_q_5_LC_9_23_5.C_ON=1'b1;
    defparam M_this_map_address_q_5_LC_9_23_5.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_5_LC_9_23_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_5_LC_9_23_5 (
            .in0(_gnd_net_),
            .in1(N__11255),
            .in2(_gnd_net_),
            .in3(N__11241),
            .lcout(M_this_map_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_4),
            .carryout(un1_M_this_map_address_q_cry_5),
            .clk(N__34575),
            .ce(),
            .sr(N__11739));
    defparam M_this_map_address_q_6_LC_9_23_6.C_ON=1'b1;
    defparam M_this_map_address_q_6_LC_9_23_6.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_6_LC_9_23_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_6_LC_9_23_6 (
            .in0(_gnd_net_),
            .in1(N__11576),
            .in2(_gnd_net_),
            .in3(N__11562),
            .lcout(M_this_map_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_5),
            .carryout(un1_M_this_map_address_q_cry_6),
            .clk(N__34575),
            .ce(),
            .sr(N__11739));
    defparam M_this_map_address_q_7_LC_9_23_7.C_ON=1'b1;
    defparam M_this_map_address_q_7_LC_9_23_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_7_LC_9_23_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_7_LC_9_23_7 (
            .in0(_gnd_net_),
            .in1(N__11546),
            .in2(_gnd_net_),
            .in3(N__11532),
            .lcout(M_this_map_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_6),
            .carryout(un1_M_this_map_address_q_cry_7),
            .clk(N__34575),
            .ce(),
            .sr(N__11739));
    defparam M_this_map_address_q_8_LC_9_24_0.C_ON=1'b1;
    defparam M_this_map_address_q_8_LC_9_24_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_8_LC_9_24_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_map_address_q_8_LC_9_24_0 (
            .in0(_gnd_net_),
            .in1(N__11516),
            .in2(_gnd_net_),
            .in3(N__11502),
            .lcout(M_this_map_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(un1_M_this_map_address_q_cry_8),
            .clk(N__34580),
            .ce(),
            .sr(N__11735));
    defparam M_this_map_address_q_9_LC_9_24_1.C_ON=1'b0;
    defparam M_this_map_address_q_9_LC_9_24_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_9_LC_9_24_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 M_this_map_address_q_9_LC_9_24_1 (
            .in0(_gnd_net_),
            .in1(N__11483),
            .in2(_gnd_net_),
            .in3(N__11499),
            .lcout(M_this_map_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34580),
            .ce(),
            .sr(N__11735));
    defparam \this_vga_signals.M_this_map_ram_write_data_i_3_LC_9_25_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_3_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_3_LC_9_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_i_3_LC_9_25_5  (
            .in0(N__32833),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18256),
            .lcout(N_89_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_i_6_LC_9_26_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_6_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_6_LC_9_26_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_i_6_LC_9_26_0  (
            .in0(N__18249),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32408),
            .lcout(N_83_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_i_5_LC_9_26_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_5_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_5_LC_9_26_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_i_5_LC_9_26_5  (
            .in0(_gnd_net_),
            .in1(N__34766),
            .in2(_gnd_net_),
            .in3(N__18248),
            .lcout(N_85_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_1_5_LC_10_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_1_5_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_1_5_LC_10_16_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_1_5_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__16753),
            .in2(_gnd_net_),
            .in3(N__16491),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_3_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_10_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_10_16_2 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_11_LC_10_16_2  (
            .in0(N__12875),
            .in1(N__11634),
            .in2(N__11448),
            .in3(N__12938),
            .lcout(\this_vga_signals.g0_6_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_10_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_10_16_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_10_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14241),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34506),
            .ce(N__14764),
            .sr(N__14729));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_10_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_10_16_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_10_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14838),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34506),
            .ce(N__14764),
            .sr(N__14729));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_10_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_10_16_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_10_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14868),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34506),
            .ce(N__14764),
            .sr(N__14729));
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_10_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_10_16_7 .LUT_INIT=16'b0111100110011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_LC_10_16_7  (
            .in0(N__17120),
            .in1(N__16534),
            .in2(N__20090),
            .in3(N__17019),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_10_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_10_17_0 .LUT_INIT=16'b0111100110011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_LC_10_17_0  (
            .in0(N__17136),
            .in1(N__16548),
            .in2(N__20078),
            .in3(N__17017),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_10_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_10_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14201),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34514),
            .ce(N__14761),
            .sr(N__14726));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_10_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_10_17_2 .LUT_INIT=16'b0111100110011111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_10_17_2  (
            .in0(N__12019),
            .in1(N__11954),
            .in2(N__11992),
            .in3(N__17016),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14837),
            .lcout(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34514),
            .ce(N__14761),
            .sr(N__14726));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_10_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_10_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14233),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34514),
            .ce(N__14761),
            .sr(N__14726));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_10_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_10_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14867),
            .lcout(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34514),
            .ce(N__14761),
            .sr(N__14726));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_0_LC_10_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_0_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_0_LC_10_17_6 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_0_LC_10_17_6  (
            .in0(N__11866),
            .in1(N__12156),
            .in2(_gnd_net_),
            .in3(N__11955),
            .lcout(\this_vga_signals.vaddress_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_10_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_10_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_10_17_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_10_17_7  (
            .in0(N__14791),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34514),
            .ce(N__14761),
            .sr(N__14726));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNI79KC_LC_10_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNI79KC_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_RNI79KC_LC_10_18_0 .LUT_INIT=16'b0000111111110001;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_RNI79KC_LC_10_18_0  (
            .in0(N__11958),
            .in1(N__11917),
            .in2(N__11616),
            .in3(N__11994),
            .lcout(\this_vga_signals.SUM_2_i_1_1_3 ),
            .ltout(\this_vga_signals.SUM_2_i_1_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_10_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_10_18_1 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_10_18_1  (
            .in0(N__17018),
            .in1(N__13043),
            .in2(N__11619),
            .in3(N__13004),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_10_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_10_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__11785),
            .in2(_gnd_net_),
            .in3(N__11800),
            .lcout(\this_vga_signals.vaddress_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1_9_LC_10_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1_9_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1_9_LC_10_18_3 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1_9_LC_10_18_3  (
            .in0(N__11595),
            .in1(N__12042),
            .in2(_gnd_net_),
            .in3(N__14813),
            .lcout(\this_vga_signals.SUM_2_i_1_1_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_4_LC_10_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_4_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_4_LC_10_18_4 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_4_LC_10_18_4  (
            .in0(N__12041),
            .in1(N__11786),
            .in2(_gnd_net_),
            .in3(N__11801),
            .lcout(\this_vga_signals.N_1_3_1 ),
            .ltout(\this_vga_signals.N_1_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_RNICPER_LC_10_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_RNICPER_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_RNICPER_LC_10_18_5 .LUT_INIT=16'b1111111101001111;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_RNICPER_LC_10_18_5  (
            .in0(N__11993),
            .in1(N__12020),
            .in2(N__11598),
            .in3(N__11957),
            .lcout(\this_vga_signals.SUM_2_i_1_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_10_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_10_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_9_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14866),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34525),
            .ce(N__14765),
            .sr(N__14730));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14796),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34525),
            .ce(N__14765),
            .sr(N__14730));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_10_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_10_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__16686),
            .in2(_gnd_net_),
            .in3(N__16476),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_1_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_10_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_10_19_1 .LUT_INIT=16'b1111011000000110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_25_LC_10_19_1  (
            .in0(N__12854),
            .in1(N__12945),
            .in2(N__11622),
            .in3(N__11841),
            .lcout(\this_vga_signals.g0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_10_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_10_19_2 .LUT_INIT=16'b1000001111001011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_24_LC_10_19_2  (
            .in0(N__12606),
            .in1(N__12207),
            .in2(N__12964),
            .in3(N__12855),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_10_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_10_19_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_10_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14264),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34534),
            .ce(N__14766),
            .sr(N__14731));
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_10_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_10_19_4 .LUT_INIT=16'b0111100010000111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_LC_10_19_4  (
            .in0(N__12176),
            .in1(N__16685),
            .in2(N__16602),
            .in3(N__12853),
            .lcout(\this_vga_signals.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_10_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_10_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14265),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34534),
            .ce(N__14766),
            .sr(N__14731));
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_10_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_10_19_6 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_LC_10_19_6  (
            .in0(N__16488),
            .in1(N__12717),
            .in2(N__16736),
            .in3(N__12651),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_3_d_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_d_LC_10_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_d_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_d_LC_10_19_7 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_d_LC_10_19_7  (
            .in0(N__12652),
            .in1(N__12605),
            .in2(N__12725),
            .in3(N__12177),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_3_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__16691),
            .in2(_gnd_net_),
            .in3(N__16459),
            .lcout(\this_vga_signals.vaddress_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_9_LC_10_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_9_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_9_LC_10_20_1 .LUT_INIT=16'b0001001100000011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIKT7S2_9_LC_10_20_1  (
            .in0(N__17169),
            .in1(N__20104),
            .in2(N__11679),
            .in3(N__11922),
            .lcout(this_vga_signals_vvisibility),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_10_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_10_20_2 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_10_20_2  (
            .in0(N__16598),
            .in1(N__16690),
            .in2(_gnd_net_),
            .in3(N__16458),
            .lcout(),
            .ltout(\this_vga_signals.un6_vvisibilitylt8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI81G42_8_LC_10_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI81G42_8_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI81G42_8_LC_10_20_3 .LUT_INIT=16'b0000100000011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI81G42_8_LC_10_20_3  (
            .in0(N__17051),
            .in1(N__17168),
            .in2(N__11682),
            .in3(N__16599),
            .lcout(\this_vga_signals.vvisibility_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_10_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_10_20_4 .LUT_INIT=16'b0111100110011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_LC_10_20_4  (
            .in0(N__16597),
            .in1(N__17170),
            .in2(N__20114),
            .in3(N__17050),
            .lcout(),
            .ltout(\this_vga_signals.if_m8_0_a3_1_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_0_LC_10_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_0_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_0_LC_10_20_5 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_0_LC_10_20_5  (
            .in0(N__12879),
            .in1(N__11670),
            .in2(N__11664),
            .in3(N__12949),
            .lcout(),
            .ltout(\this_vga_signals.g0_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_10_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_10_20_6 .LUT_INIT=16'b0111011100010111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_LC_10_20_6  (
            .in0(N__16469),
            .in1(N__15282),
            .in2(N__11661),
            .in3(N__11658),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_a2_1_LC_10_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_a2_1_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_a2_1_LC_10_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_0_a2_1_LC_10_20_7  (
            .in0(N__11652),
            .in1(N__13383),
            .in2(N__11643),
            .in3(N__13307),
            .lcout(\this_vga_signals.g0_i_x4_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_10_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_10_21_1 .LUT_INIT=16'b0111100110011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_23_LC_10_21_1  (
            .in0(N__17166),
            .in1(N__16596),
            .in2(N__20115),
            .in3(N__17049),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_10_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_10_21_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__19025),
            .in2(_gnd_net_),
            .in3(N__19102),
            .lcout(\this_vga_signals.M_vcounter_q_379_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIS6TO_9_LC_10_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIS6TO_9_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIS6TO_9_LC_10_21_3 .LUT_INIT=16'b1111000000000101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIS6TO_9_LC_10_21_3  (
            .in0(N__13938),
            .in1(_gnd_net_),
            .in2(N__14606),
            .in3(N__14174),
            .lcout(\this_vga_signals.SUM_3_1_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_10_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_10_22_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_10_22_6 .LUT_INIT=16'b0011111111000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(N__19064),
            .in2(N__12288),
            .in3(N__13980),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34555),
            .ce(),
            .sr(N__12374));
    defparam \this_vga_signals.M_hcounter_q_0_LC_10_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_10_22_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_10_22_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_10_22_7  (
            .in0(N__19065),
            .in1(N__12283),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34555),
            .ce(),
            .sr(N__12374));
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_10_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_10_23_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(N__12363),
            .in2(_gnd_net_),
            .in3(N__19055),
            .lcout(\this_vga_signals.N_692_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_24_4 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_24_4  (
            .in0(N__14172),
            .in1(N__14592),
            .in2(_gnd_net_),
            .in3(N__14678),
            .lcout(this_vga_signals_hvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_RNIC68K4_9_LC_10_24_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_RNIC68K4_9_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \this_reset_cond.M_stage_q_RNIC68K4_9_LC_10_24_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_reset_cond.M_stage_q_RNIC68K4_9_LC_10_24_7  (
            .in0(_gnd_net_),
            .in1(N__18282),
            .in2(_gnd_net_),
            .in3(N__34113),
            .lcout(M_stage_q_RNIC68K4_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_0_LC_11_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_0_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_0_LC_11_17_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_0_LC_11_17_0  (
            .in0(N__12168),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11873),
            .lcout(\this_vga_signals.vaddress_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_11_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_11_17_1 .LUT_INIT=16'b0111100110011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_20_LC_11_17_1  (
            .in0(N__17122),
            .in1(N__16549),
            .in2(N__20092),
            .in3(N__17020),
            .lcout(),
            .ltout(\this_vga_signals.if_m8_0_a3_1_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_11_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_11_17_2 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_18_LC_11_17_2  (
            .in0(N__11711),
            .in1(N__12937),
            .in2(N__11697),
            .in3(N__12862),
            .lcout(\this_vga_signals.g0_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_11_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_11_17_3 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_11_17_3  (
            .in0(N__11871),
            .in1(N__12166),
            .in2(_gnd_net_),
            .in3(N__11956),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_11_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14258),
            .lcout(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34507),
            .ce(N__14763),
            .sr(N__14725));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_11_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_11_17_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__11870),
            .in2(_gnd_net_),
            .in3(N__12165),
            .lcout(\this_vga_signals.vaddress_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_1_LC_11_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_1_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_1_LC_11_17_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_1_LC_11_17_6  (
            .in0(N__12167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11872),
            .lcout(\this_vga_signals.vaddress_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_11_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_11_17_7 .LUT_INIT=16'b0111100110011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_21_LC_11_17_7  (
            .in0(N__17121),
            .in1(N__16550),
            .in2(N__20091),
            .in3(N__17021),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_11_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_11_18_0 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_11_18_0  (
            .in0(N__11982),
            .in1(N__11952),
            .in2(N__12021),
            .in3(N__12039),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_11_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_11_18_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_9_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__16583),
            .in2(_gnd_net_),
            .in3(N__12852),
            .lcout(\this_vga_signals.N_5_i_0 ),
            .ltout(\this_vga_signals.N_5_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJ8O74_0_5_LC_11_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJ8O74_0_5_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJ8O74_0_5_LC_11_18_2 .LUT_INIT=16'b1110001010001011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIJ8O74_0_5_LC_11_18_2  (
            .in0(N__11820),
            .in1(N__16743),
            .in2(N__11811),
            .in3(N__16489),
            .lcout(\this_vga_signals.g1_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14240),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34515),
            .ce(N__14767),
            .sr(N__14727));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_18_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_11_18_4  (
            .in0(N__11808),
            .in1(N__11802),
            .in2(N__14814),
            .in3(N__11787),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_11_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_11_18_5 .LUT_INIT=16'b0000110100011011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_11_18_5  (
            .in0(N__12040),
            .in1(N__12015),
            .in2(N__11997),
            .in3(N__11983),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_11_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_11_18_6 .LUT_INIT=16'b1011000011010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_11_18_6  (
            .in0(N__11964),
            .in1(N__11953),
            .in2(N__11925),
            .in3(N__11918),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_11_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_11_18_7 .LUT_INIT=16'b1000111001010101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_11_18_7  (
            .in0(N__12944),
            .in1(N__12581),
            .in2(N__11901),
            .in3(N__12203),
            .lcout(\this_vga_signals.mult1_un47_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIC2H0Q9_1_LC_11_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIC2H0Q9_1_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIC2H0Q9_1_LC_11_19_0 .LUT_INIT=16'b0111110110000010;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIC2H0Q9_1_LC_11_19_0  (
            .in0(N__12426),
            .in1(N__12243),
            .in2(N__12093),
            .in3(N__13056),
            .lcout(\this_vga_signals.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_11_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_11_19_1 .LUT_INIT=16'b1000010110101101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_15_LC_11_19_1  (
            .in0(N__12205),
            .in1(N__11886),
            .in2(N__12963),
            .in3(N__12851),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x0_LC_11_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x0_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x0_LC_11_19_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x0_LC_11_19_2  (
            .in0(N__12646),
            .in1(N__12180),
            .in2(N__12604),
            .in3(N__12541),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_ns_LC_11_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_ns_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_ns_LC_11_19_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_ns_LC_11_19_3  (
            .in0(N__12542),
            .in1(_gnd_net_),
            .in2(N__11877),
            .in3(N__12712),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_11_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_11_19_4 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_11_19_4  (
            .in0(N__11874),
            .in1(N__12178),
            .in2(_gnd_net_),
            .in3(N__11840),
            .lcout(),
            .ltout(\this_vga_signals.if_N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_11_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_11_19_5 .LUT_INIT=16'b0000110100001110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_LC_11_19_5  (
            .in0(N__12939),
            .in1(N__12589),
            .in2(N__11823),
            .in3(N__12849),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_19_6 .LUT_INIT=16'b0100001010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_19_6  (
            .in0(N__12850),
            .in1(N__12943),
            .in2(N__12603),
            .in3(N__12204),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i ),
            .ltout(\this_vga_signals.mult1_un54_sum_axb2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_571_LC_11_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_571_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_571_LC_11_19_7 .LUT_INIT=16'b0001111001111000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_571_LC_11_19_7  (
            .in0(N__12179),
            .in1(N__12593),
            .in2(N__12132),
            .in3(N__12645),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_571 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJ8O74_5_LC_11_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJ8O74_5_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJ8O74_5_LC_11_20_0 .LUT_INIT=16'b1110100001110001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIJ8O74_5_LC_11_20_0  (
            .in0(N__16711),
            .in1(N__16426),
            .in2(N__12129),
            .in3(N__12114),
            .lcout(),
            .ltout(\this_vga_signals.g1_2_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIOV1AF_3_LC_11_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIOV1AF_3_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIOV1AF_3_LC_11_20_1 .LUT_INIT=16'b0100010011010100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIOV1AF_3_LC_11_20_1  (
            .in0(N__16427),
            .in1(N__15275),
            .in2(N__12105),
            .in3(N__12060),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI5FISK_2_LC_11_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI5FISK_2_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI5FISK_2_LC_11_20_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI5FISK_2_LC_11_20_2  (
            .in0(N__16712),
            .in1(N__15396),
            .in2(N__12102),
            .in3(N__12099),
            .lcout(\this_vga_signals.g1_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_0_LC_11_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_0_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_0_LC_11_20_3 .LUT_INIT=16'b1111100101100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_m2_0_LC_11_20_3  (
            .in0(N__16424),
            .in1(N__16707),
            .in2(N__12081),
            .in3(N__12066),
            .lcout(\this_vga_signals.g0_1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_11_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_11_20_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_17_LC_11_20_4  (
            .in0(N__12713),
            .in1(N__16425),
            .in2(N__16742),
            .in3(N__12654),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_3_d_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIHM8LF_3_LC_11_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIHM8LF_3_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIHM8LF_3_LC_11_20_5 .LUT_INIT=16'b0101101001010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIHM8LF_3_LC_11_20_5  (
            .in0(N__15298),
            .in1(_gnd_net_),
            .in2(N__12054),
            .in3(N__12051),
            .lcout(),
            .ltout(\this_vga_signals.g2_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQC7Q91_2_LC_11_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQC7Q91_2_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQC7Q91_2_LC_11_20_6 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQC7Q91_2_LC_11_20_6  (
            .in0(N__15393),
            .in1(N__13377),
            .in2(N__12045),
            .in3(N__13293),
            .lcout(),
            .ltout(\this_vga_signals.g3_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_11_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_11_20_7 .LUT_INIT=16'b1011001111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_0_LC_11_20_7  (
            .in0(N__15297),
            .in1(N__13211),
            .in2(N__12246),
            .in3(N__12747),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNII65L3_9_LC_11_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNII65L3_9_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNII65L3_9_LC_11_21_0 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNII65L3_9_LC_11_21_0  (
            .in0(N__14597),
            .in1(N__14680),
            .in2(N__14181),
            .in3(N__22956),
            .lcout(M_this_vga_ramdac_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_11_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_11_21_1 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_11_21_1  (
            .in0(N__12280),
            .in1(N__12321),
            .in2(N__13998),
            .in3(N__13826),
            .lcout(),
            .ltout(\this_vga_signals.M_hcounter_d7lt7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_11_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_11_21_2 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_11_21_2  (
            .in0(N__12327),
            .in1(N__14596),
            .in2(N__12237),
            .in3(N__14679),
            .lcout(\this_vga_signals.M_hcounter_d7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_11_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_11_21_3 .LUT_INIT=16'b0001001001001000;
    LogicCell40 \this_vga_signals.un4_haddress_if_m2_0_LC_11_21_3  (
            .in0(N__14040),
            .in1(N__13827),
            .in2(N__14101),
            .in3(N__13463),
            .lcout(\this_vga_signals.if_m2_0 ),
            .ltout(\this_vga_signals.if_m2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_11_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_11_21_4 .LUT_INIT=16'b0010010001001101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_11_21_4  (
            .in0(N__13464),
            .in1(N__14093),
            .in2(N__12234),
            .in3(N__13830),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_0_1_LC_11_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_0_1_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_0_1_LC_11_21_5 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_0_1_LC_11_21_5  (
            .in0(N__12281),
            .in1(N__13088),
            .in2(N__13999),
            .in3(N__13147),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un89_sum_c3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNII3DE13_2_LC_11_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNII3DE13_2_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNII3DE13_2_LC_11_21_6 .LUT_INIT=16'b0110010110100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNII3DE13_2_LC_11_21_6  (
            .in0(N__13148),
            .in1(N__14041),
            .in2(N__12231),
            .in3(N__13120),
            .lcout(),
            .ltout(\this_vga_signals.haddress_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI7BUL75_2_LC_11_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI7BUL75_2_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI7BUL75_2_LC_11_21_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI7BUL75_2_LC_11_21_7  (
            .in0(N__13155),
            .in1(N__15558),
            .in2(N__12228),
            .in3(N__13089),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_11_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_11_22_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_11_22_0  (
            .in0(N__13880),
            .in1(N__14158),
            .in2(_gnd_net_),
            .in3(N__13932),
            .lcout(\this_vga_signals.M_hcounter_d7lto7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_11_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_11_22_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__14027),
            .in2(_gnd_net_),
            .in3(N__14073),
            .lcout(\this_vga_signals.un2_hsynclto3_0 ),
            .ltout(\this_vga_signals.un2_hsynclto3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_0_LC_11_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_0_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_0_LC_11_22_3 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI58GD1_0_0_LC_11_22_3  (
            .in0(N__13990),
            .in1(N__12287),
            .in2(N__12315),
            .in3(N__13825),
            .lcout(),
            .ltout(\this_vga_signals.un2_hsynclto6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIKCQ82_7_LC_11_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIKCQ82_7_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIKCQ82_7_LC_11_22_4 .LUT_INIT=16'b1100110010001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIKCQ82_7_LC_11_22_4  (
            .in0(N__13881),
            .in1(N__14159),
            .in2(N__12312),
            .in3(N__13933),
            .lcout(\this_vga_signals.un2_hsynclt8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_11_22_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_11_22_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_11_22_7  (
            .in0(N__15618),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15817),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_23_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__12282),
            .in2(N__13994),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_11_23_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_11_23_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_11_23_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_11_23_1  (
            .in0(N__19060),
            .in1(N__14038),
            .in2(_gnd_net_),
            .in3(N__12255),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__34556),
            .ce(),
            .sr(N__12378));
    defparam \this_vga_signals.M_hcounter_q_3_LC_11_23_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_11_23_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_11_23_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_11_23_2  (
            .in0(N__19057),
            .in1(N__14088),
            .in2(_gnd_net_),
            .in3(N__12252),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__34556),
            .ce(),
            .sr(N__12378));
    defparam \this_vga_signals.M_hcounter_q_4_LC_11_23_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_11_23_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_11_23_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_11_23_3  (
            .in0(N__19061),
            .in1(N__13824),
            .in2(_gnd_net_),
            .in3(N__12249),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__34556),
            .ce(),
            .sr(N__12378));
    defparam \this_vga_signals.M_hcounter_q_5_LC_11_23_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_11_23_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_11_23_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_11_23_4  (
            .in0(N__19058),
            .in1(N__13882),
            .in2(_gnd_net_),
            .in3(N__12405),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__34556),
            .ce(),
            .sr(N__12378));
    defparam \this_vga_signals.M_hcounter_q_6_LC_11_23_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_11_23_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_11_23_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_11_23_5  (
            .in0(N__19062),
            .in1(N__13937),
            .in2(_gnd_net_),
            .in3(N__12402),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__34556),
            .ce(),
            .sr(N__12378));
    defparam \this_vga_signals.M_hcounter_q_7_LC_11_23_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_11_23_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_11_23_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_11_23_6  (
            .in0(N__19059),
            .in1(N__14171),
            .in2(_gnd_net_),
            .in3(N__12399),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__34556),
            .ce(),
            .sr(N__12378));
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_23_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_23_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_11_23_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_11_23_7  (
            .in0(N__19063),
            .in1(N__14671),
            .in2(_gnd_net_),
            .in3(N__12396),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__34556),
            .ce(),
            .sr(N__12378));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_11_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_11_24_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_11_24_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_11_24_0  (
            .in0(_gnd_net_),
            .in1(N__14591),
            .in2(_gnd_net_),
            .in3(N__12393),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34567),
            .ce(N__12390),
            .sr(N__12373));
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_12_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_12_17_0 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_26_LC_12_17_0  (
            .in0(N__16477),
            .in1(N__12726),
            .in2(N__16776),
            .in3(N__12653),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_3_d_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_3_LC_12_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_3_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_3_LC_12_17_1 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_3_LC_12_17_1  (
            .in0(N__16478),
            .in1(N__12678),
            .in2(_gnd_net_),
            .in3(N__12546),
            .lcout(\this_vga_signals.g0_i_x4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_x0_LC_12_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_x0_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_x0_LC_12_17_2 .LUT_INIT=16'b1011111011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_x0_LC_12_17_2  (
            .in0(N__15263),
            .in1(N__12782),
            .in2(N__13308),
            .in3(N__12420),
            .lcout(),
            .ltout(\this_vga_signals.g0_3_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_ns_LC_12_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_ns_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_ns_LC_12_17_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_ns_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__13389),
            .in2(N__12339),
            .in3(N__12411),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_0_a2_LC_12_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_0_a2_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_0_a2_LC_12_17_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_0_a2_LC_12_17_4  (
            .in0(N__13388),
            .in1(N__12783),
            .in2(N__15291),
            .in3(N__13306),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_12_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_12_17_5 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_1_LC_12_17_5  (
            .in0(N__15361),
            .in1(N__13070),
            .in2(_gnd_net_),
            .in3(N__12738),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_12_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_12_17_6 .LUT_INIT=16'b1000111011101000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_LC_12_17_6  (
            .in0(N__15463),
            .in1(N__15425),
            .in2(N__12468),
            .in3(N__12465),
            .lcout(\this_vga_signals.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIMRO4P_3_LC_12_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIMRO4P_3_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIMRO4P_3_LC_12_18_0 .LUT_INIT=16'b1001011010011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIMRO4P_3_LC_12_18_0  (
            .in0(N__13369),
            .in1(N__15234),
            .in2(N__12450),
            .in3(N__12441),
            .lcout(),
            .ltout(\this_vga_signals.g1_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIUC6F91_1_LC_12_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIUC6F91_1_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIUC6F91_1_LC_12_18_1 .LUT_INIT=16'b0000011001100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIUC6F91_1_LC_12_18_1  (
            .in0(N__15405),
            .in1(N__15456),
            .in2(N__12429),
            .in3(N__13294),
            .lcout(\this_vga_signals.g0_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_12_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_12_18_2 .LUT_INIT=16'b0001001000100001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_12_18_2  (
            .in0(N__13367),
            .in1(N__15230),
            .in2(N__12776),
            .in3(N__13270),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_1_LC_12_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_1_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_1_LC_12_18_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_a2_1_LC_12_18_3  (
            .in0(N__16455),
            .in1(_gnd_net_),
            .in2(N__13296),
            .in3(N__15226),
            .lcout(\this_vga_signals.g0_2_0_a2_1 ),
            .ltout(\this_vga_signals.g0_2_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_x1_LC_12_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_x1_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_x1_LC_12_18_4 .LUT_INIT=16'b0110111101101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_x1_LC_12_18_4  (
            .in0(N__12772),
            .in1(N__13275),
            .in2(N__12414),
            .in3(N__15235),
            .lcout(\this_vga_signals.g0_3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_13_x0_LC_12_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_13_x0_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_13_x0_LC_12_18_5 .LUT_INIT=16'b0110100100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_13_x0_LC_12_18_5  (
            .in0(N__12674),
            .in1(N__13368),
            .in2(N__15271),
            .in3(N__12538),
            .lcout(),
            .ltout(\this_vga_signals.g0_13_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_13_ns_LC_12_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_13_ns_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_13_ns_LC_12_18_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_13_ns_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__12660),
            .in2(N__12741),
            .in3(N__13274),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x0_LC_12_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x0_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x0_LC_12_18_7 .LUT_INIT=16'b1010010011100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x0_LC_12_18_7  (
            .in0(N__12582),
            .in1(N__15225),
            .in2(N__16484),
            .in3(N__12537),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_12_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_12_19_0 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_14_LC_12_19_0  (
            .in0(N__16394),
            .in1(N__12732),
            .in2(N__16775),
            .in3(N__12711),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_3_d_2 ),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_3_d_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_13_x1_LC_12_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_13_x1_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_13_x1_LC_12_19_1 .LUT_INIT=16'b1100011000111001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_13_x1_LC_12_19_1  (
            .in0(N__12540),
            .in1(N__15240),
            .in2(N__12663),
            .in3(N__13361),
            .lcout(\this_vga_signals.g0_13_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_ns_LC_12_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_ns_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_ns_LC_12_19_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_ns_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__12647),
            .in2(N__12510),
            .in3(N__12615),
            .lcout(\this_vga_signals.mult1_un61_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIANU4Q_3_LC_12_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIANU4Q_3_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIANU4Q_3_LC_12_19_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIANU4Q_3_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__15241),
            .in2(N__12609),
            .in3(N__13362),
            .lcout(\this_vga_signals.M_vcounter_q_RNIANU4QZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x1_LC_12_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x1_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x1_LC_12_19_4 .LUT_INIT=16'b0110010011100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_x1_LC_12_19_4  (
            .in0(N__12597),
            .in1(N__16366),
            .in2(N__15272),
            .in3(N__12539),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNITVMCU_3_LC_12_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNITVMCU_3_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNITVMCU_3_LC_12_19_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNITVMCU_3_LC_12_19_5  (
            .in0(N__12501),
            .in1(N__13363),
            .in2(N__15302),
            .in3(N__13276),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_RNITVMCUZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI2KDQ22_3_LC_12_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI2KDQ22_3_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI2KDQ22_3_LC_12_19_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI2KDQ22_3_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__12495),
            .in2(N__12486),
            .in3(N__12483),
            .lcout(),
            .ltout(\this_vga_signals.g2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI0FHHA4_2_LC_12_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI0FHHA4_2_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI0FHHA4_2_LC_12_19_7 .LUT_INIT=16'b1010111001010001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI0FHHA4_2_LC_12_19_7  (
            .in0(N__13071),
            .in1(N__15387),
            .in2(N__13059),
            .in3(N__13212),
            .lcout(\this_vga_signals.g0_0_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_12_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_12_20_0 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_LC_12_20_0  (
            .in0(N__13050),
            .in1(N__17068),
            .in2(N__13032),
            .in3(N__13011),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_axb1_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_12_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_12_20_1 .LUT_INIT=16'b0011100111001001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_12_20_1  (
            .in0(N__12966),
            .in1(N__16764),
            .in2(N__12993),
            .in3(N__12801),
            .lcout(\this_vga_signals.g0_i_x4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_4_1_LC_12_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_4_1_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_4_1_LC_12_20_2 .LUT_INIT=16'b0001011111101000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_4_1_LC_12_20_2  (
            .in0(N__15267),
            .in1(N__12768),
            .in2(N__16451),
            .in3(N__13384),
            .lcout(),
            .ltout(\this_vga_signals.g0_i_x4_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_4_LC_12_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_4_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_4_LC_12_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_4_LC_12_20_3  (
            .in0(N__15404),
            .in1(N__12990),
            .in2(N__12984),
            .in3(N__13269),
            .lcout(\this_vga_signals.g0_i_x4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_12_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_12_20_4 .LUT_INIT=16'b0100100011011110;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_0_LC_12_20_4  (
            .in0(N__16385),
            .in1(N__12965),
            .in2(N__16777),
            .in3(N__12880),
            .lcout(\this_vga_signals.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_12_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_12_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_12_20_5  (
            .in0(N__15274),
            .in1(N__13366),
            .in2(N__16481),
            .in3(N__13268),
            .lcout(\this_vga_signals.g0_2_0_a2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_12_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_12_20_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_12_20_6  (
            .in0(N__13365),
            .in1(_gnd_net_),
            .in2(N__13295),
            .in3(N__12767),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a2_LC_12_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a2_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a2_LC_12_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_0_a2_LC_12_20_7  (
            .in0(N__15273),
            .in1(N__13364),
            .in2(N__16480),
            .in3(N__13264),
            .lcout(\this_vga_signals.N_4_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_12_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_12_21_0 .LUT_INIT=16'b0011100101100011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_12_21_0  (
            .in0(N__13828),
            .in1(N__13492),
            .in2(N__14102),
            .in3(N__13465),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_12_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_12_21_1 .LUT_INIT=16'b0010010011011011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_12_21_1  (
            .in0(N__14100),
            .in1(N__14042),
            .in2(N__13197),
            .in3(N__13440),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI49VKF_9_LC_12_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI49VKF_9_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI49VKF_9_LC_12_21_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI49VKF_9_LC_12_21_2  (
            .in0(N__13173),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15559),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_12_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_12_21_3 .LUT_INIT=16'b1110000100011110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_12_21_3  (
            .in0(N__13179),
            .in1(N__13172),
            .in2(N__13497),
            .in3(N__13164),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_0_LC_12_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_0_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_0_LC_12_21_4 .LUT_INIT=16'b1010101001110001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_0_LC_12_21_4  (
            .in0(N__14043),
            .in1(N__14000),
            .in2(N__13158),
            .in3(N__13087),
            .lcout(\this_vga_signals.mult1_un82_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIIHKHP3_9_LC_12_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIIHKHP3_9_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIIHKHP3_9_LC_12_21_5 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIIHKHP3_9_LC_12_21_5  (
            .in0(N__15560),
            .in1(N__13149),
            .in2(N__13134),
            .in3(N__13121),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_12_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_12_21_6 .LUT_INIT=16'b0011011001101100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_12_21_6  (
            .in0(N__13829),
            .in1(N__13493),
            .in2(N__14103),
            .in3(N__13466),
            .lcout(\this_vga_signals.mult1_un75_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_12_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_12_22_0 .LUT_INIT=16'b1010111010001010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_12_22_0  (
            .in0(N__14120),
            .in1(N__13413),
            .in2(N__13884),
            .in3(N__13931),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_12_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_12_22_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(N__13878),
            .in2(N__13500),
            .in3(N__13809),
            .lcout(\this_vga_signals.mult1_un68_sum_axb2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x1_LC_12_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x1_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x1_LC_12_22_2 .LUT_INIT=16'b0010111110001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x1_LC_12_22_2  (
            .in0(N__13808),
            .in1(N__13412),
            .in2(N__13883),
            .in3(N__13930),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_x1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_ns_LC_12_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_ns_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_ns_LC_12_22_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_ns_LC_12_22_3  (
            .in0(_gnd_net_),
            .in1(N__14121),
            .in2(N__13482),
            .in3(N__13401),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_12_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_12_22_4 .LUT_INIT=16'b0000000001010010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_12_22_4  (
            .in0(N__13877),
            .in1(N__13395),
            .in2(N__13479),
            .in3(N__14109),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_12_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_12_22_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(N__14087),
            .in2(N__13443),
            .in3(N__13810),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI18DB6_9_LC_12_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI18DB6_9_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI18DB6_9_LC_12_22_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI18DB6_9_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(N__13434),
            .in2(_gnd_net_),
            .in3(N__15561),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_12_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_12_23_0 .LUT_INIT=16'b1001010111010111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_12_23_0  (
            .in0(N__14663),
            .in1(N__14160),
            .in2(N__14601),
            .in3(N__13924),
            .lcout(\this_vga_signals.SUM_3 ),
            .ltout(\this_vga_signals.SUM_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x0_LC_12_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x0_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x0_LC_12_23_1 .LUT_INIT=16'b0101101000010010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_x0_LC_12_23_1  (
            .in0(N__13926),
            .in1(N__13869),
            .in2(N__13404),
            .in3(N__13805),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_12_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_12_23_2 .LUT_INIT=16'b0010100000000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_12_23_2  (
            .in0(N__14665),
            .in1(N__14164),
            .in2(N__14602),
            .in3(N__13927),
            .lcout(\this_vga_signals.N_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_12_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_12_23_3 .LUT_INIT=16'b0101011010010101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_12_23_3  (
            .in0(N__13925),
            .in1(N__14587),
            .in2(N__14173),
            .in3(N__14664),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ),
            .ltout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_LC_12_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_LC_12_23_4 .LUT_INIT=16'b0000001000001110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_LC_12_23_4  (
            .in0(N__13806),
            .in1(N__13879),
            .in2(N__14112),
            .in3(N__13928),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI3O9R_1_LC_12_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI3O9R_1_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI3O9R_1_LC_12_23_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI3O9R_1_LC_12_23_6  (
            .in0(N__14089),
            .in1(N__14039),
            .in2(_gnd_net_),
            .in3(N__14001),
            .lcout(),
            .ltout(\this_vga_signals.un4_hsynclt4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIFPJM1_5_LC_12_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIFPJM1_5_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIFPJM1_5_LC_12_23_7 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIFPJM1_5_LC_12_23_7  (
            .in0(N__13929),
            .in1(N__13870),
            .in2(N__13833),
            .in3(N__13807),
            .lcout(\this_vga_signals.un4_hsynclt8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_3_0_0_LC_12_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_3_0_0_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_3_0_0_LC_12_24_4 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a3_3_0_0_LC_12_24_4  (
            .in0(N__33492),
            .in1(N__34757),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_N_419_i_i_0_a3_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_i_2_LC_12_25_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_2_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_2_LC_12_25_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_i_2_LC_12_25_1  (
            .in0(N__18241),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33443),
            .lcout(N_91_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_i_1_LC_12_25_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_1_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_1_LC_12_25_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_i_1_LC_12_25_6  (
            .in0(_gnd_net_),
            .in1(N__32912),
            .in2(_gnd_net_),
            .in3(N__18240),
            .lcout(N_93_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI43UU_6_LC_13_13_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI43UU_6_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI43UU_6_LC_13_13_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \this_ppu.M_state_q_RNI43UU_6_LC_13_13_6  (
            .in0(N__13740),
            .in1(N__29990),
            .in2(N__30164),
            .in3(N__31089),
            .lcout(M_this_ppu_sprites_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI43UU_2_6_LC_13_15_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI43UU_2_6_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI43UU_2_6_LC_13_15_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \this_ppu.M_state_q_RNI43UU_2_6_LC_13_15_6  (
            .in0(N__14523),
            .in1(N__30000),
            .in2(N__30162),
            .in3(N__31116),
            .lcout(M_this_ppu_sprites_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_13_17_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_13_17_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_13_17_0  (
            .in0(N__18997),
            .in1(N__15429),
            .in2(N__19131),
            .in3(N__19123),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__34487),
            .ce(),
            .sr(N__14723));
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_17_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_17_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_13_17_1  (
            .in0(N__18999),
            .in1(N__15457),
            .in2(_gnd_net_),
            .in3(N__14277),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__34487),
            .ce(),
            .sr(N__14723));
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_17_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_17_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_13_17_2  (
            .in0(N__18998),
            .in1(N__15360),
            .in2(_gnd_net_),
            .in3(N__14274),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__34487),
            .ce(),
            .sr(N__14723));
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_17_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_17_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_13_17_3  (
            .in0(N__19000),
            .in1(N__15236),
            .in2(_gnd_net_),
            .in3(N__14271),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__34487),
            .ce(),
            .sr(N__14723));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_17_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__16479),
            .in2(_gnd_net_),
            .in3(N__14268),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_17_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__16760),
            .in2(_gnd_net_),
            .in3(N__14244),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_17_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__16608),
            .in2(_gnd_net_),
            .in3(N__14208),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_17_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__17072),
            .in2(_gnd_net_),
            .in3(N__14184),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_18_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__17171),
            .in2(_gnd_net_),
            .in3(N__14874),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_13_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_13_18_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__20102),
            .in2(_gnd_net_),
            .in3(N__14871),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_13_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_13_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_13_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14825),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34498),
            .ce(N__14768),
            .sr(N__14724));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_13_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_13_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14795),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34516),
            .ce(N__14769),
            .sr(N__14728));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIR18F4_9_LC_13_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIR18F4_9_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIR18F4_9_LC_13_21_0 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIR18F4_9_LC_13_21_0  (
            .in0(N__14690),
            .in1(N__14631),
            .in2(N__14622),
            .in3(N__14607),
            .lcout(this_vga_signals_hsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_13_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_13_21_3 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_13_21_3  (
            .in0(N__15832),
            .in1(N__15895),
            .in2(N__15875),
            .in3(N__19113),
            .lcout(\this_vga_signals.M_pcounter_q_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_13_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_13_21_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_13_21_5 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_1_LC_13_21_5  (
            .in0(N__15834),
            .in1(N__15896),
            .in2(N__15876),
            .in3(N__19115),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34526),
            .ce(N__19009),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_13_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_13_21_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_13_21_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_0_LC_13_21_6  (
            .in0(N__19114),
            .in1(N__15833),
            .in2(_gnd_net_),
            .in3(N__15714),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34526),
            .ce(N__19009),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_13_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_13_21_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_13_21_7  (
            .in0(N__15831),
            .in1(N__15713),
            .in2(_gnd_net_),
            .in3(N__19112),
            .lcout(\this_vga_signals.M_pcounter_q_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_13_22_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_13_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__15805),
            .in2(_gnd_net_),
            .in3(N__16233),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_i_0_LC_13_25_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_0_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_0_LC_13_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_i_0_LC_13_25_5  (
            .in0(N__33750),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18239),
            .lcout(N_95_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_14_17_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_14_17_1 .LUT_INIT=16'b0010011000100110;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_14_17_1  (
            .in0(N__18730),
            .in1(N__18773),
            .in2(N__18840),
            .in3(_gnd_net_),
            .lcout(\this_vga_ramdac.N_24_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_17_2 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_17_2  (
            .in0(N__15455),
            .in1(N__15421),
            .in2(N__15365),
            .in3(N__15197),
            .lcout(\this_vga_signals.M_vcounter_d7lt8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI43UU_0_6_LC_14_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI43UU_0_6_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI43UU_0_6_LC_14_17_4 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \this_ppu.M_state_q_RNI43UU_0_6_LC_14_17_4  (
            .in0(N__15150),
            .in1(N__29941),
            .in2(N__30163),
            .in3(N__31161),
            .lcout(M_this_ppu_sprites_addr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_14_17_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_14_17_6 .LUT_INIT=16'b0110010100101011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_14_17_6  (
            .in0(N__18883),
            .in1(N__18832),
            .in2(N__18784),
            .in3(N__18729),
            .lcout(\this_vga_ramdac.m19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_14_17_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_14_17_7 .LUT_INIT=16'b0011001100101111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_14_17_7  (
            .in0(N__18731),
            .in1(N__18884),
            .in2(N__18839),
            .in3(N__18777),
            .lcout(\this_vga_ramdac.m6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_14_18_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_14_18_1 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_14_18_1  (
            .in0(N__14904),
            .in1(N__16263),
            .in2(N__14891),
            .in3(N__22870),
            .lcout(\this_vga_ramdac.N_2862_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34488),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.G_330_LC_14_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.G_330_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.G_330_LC_14_18_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.G_330_LC_14_18_3  (
            .in0(N__15701),
            .in1(N__16279),
            .in2(_gnd_net_),
            .in3(N__34104),
            .lcout(\this_vga_signals.GZ0Z_330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_14_18_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_14_18_4 .LUT_INIT=16'b0100011100100101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_14_18_4  (
            .in0(N__18871),
            .in1(N__18820),
            .in2(N__18785),
            .in3(N__18715),
            .lcout(\this_vga_ramdac.i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_1_LC_14_18_5 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_1_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_1_LC_14_18_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clk.M_counter_q_1_LC_14_18_5  (
            .in0(N__15702),
            .in1(N__16280),
            .in2(_gnd_net_),
            .in3(N__34105),
            .lcout(this_pixel_clk_M_counter_q_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34488),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_14_18_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_14_18_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_14_18_6  (
            .in0(N__16110),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15791),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_14_19_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_14_19_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_14_19_0 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_14_19_0  (
            .in0(N__15672),
            .in1(N__16255),
            .in2(N__15653),
            .in3(N__22859),
            .lcout(\this_vga_ramdac.N_2863_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34499),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_14_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_14_19_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_14_19_2 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_2_LC_14_19_2  (
            .in0(N__15728),
            .in1(_gnd_net_),
            .in2(N__15849),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_this_vga_signals_pixel_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34499),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_14_19_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_14_19_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_14_19_3 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_14_19_3  (
            .in0(N__22862),
            .in1(N__15761),
            .in2(N__16266),
            .in3(N__15636),
            .lcout(\this_vga_ramdac.N_2867_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34499),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_14_19_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_14_19_4 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_14_19_4  (
            .in0(N__15627),
            .in1(N__16259),
            .in2(N__15614),
            .in3(N__22861),
            .lcout(\this_vga_ramdac.N_2866_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34499),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_2_RNIH7PG8_LC_14_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_2_RNIH7PG8_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_2_RNIH7PG8_LC_14_19_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_2_RNIH7PG8_LC_14_19_5  (
            .in0(N__15597),
            .in1(N__15845),
            .in2(_gnd_net_),
            .in3(N__15727),
            .lcout(M_pcounter_q_ret_2_RNIH7PG8),
            .ltout(M_pcounter_q_ret_2_RNIH7PG8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_14_19_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_14_19_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_14_19_6 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_q_ret_LC_14_19_6  (
            .in0(N__15790),
            .in1(N__15591),
            .in2(N__15525),
            .in3(N__22863),
            .lcout(\this_vga_ramdac.M_this_vga_ramdac_en_reto_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34499),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_14_19_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_14_19_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_14_19_7 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_14_19_7  (
            .in0(N__22860),
            .in1(N__16109),
            .in2(N__16265),
            .in3(N__16125),
            .lcout(\this_vga_ramdac.N_2864_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34499),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI0F523_0_6_LC_14_20_2.C_ON=1'b0;
    defparam M_this_state_q_RNI0F523_0_6_LC_14_20_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI0F523_0_6_LC_14_20_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 M_this_state_q_RNI0F523_0_6_LC_14_20_2 (
            .in0(N__22901),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(dma_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_14_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_14_20_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_14_20_4  (
            .in0(N__15897),
            .in1(N__15882),
            .in2(_gnd_net_),
            .in3(N__19007),
            .lcout(\this_vga_signals.N_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_14_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_14_20_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_14_20_6  (
            .in0(N__15874),
            .in1(N__15855),
            .in2(_gnd_net_),
            .in3(N__19008),
            .lcout(\this_vga_signals.N_3_0 ),
            .ltout(\this_vga_signals.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_LC_14_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_14_20_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_14_20_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15837),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_pcounter_q_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34508),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_14_21_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_14_21_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_14_21_2  (
            .in0(N__15804),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15765),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_14_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_14_21_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_14_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15729),
            .lcout(\this_vga_signals.M_pcounter_q_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34517),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_14_23_3.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_14_23_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_14_23_3.LUT_INIT=16'b0101000011011000;
    LogicCell40 M_this_data_count_q_13_LC_14_23_3 (
            .in0(N__18586),
            .in1(N__20463),
            .in2(N__16182),
            .in3(N__34125),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34535),
            .ce(N__18483),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_10_LC_14_24_3.C_ON=1'b0;
    defparam M_this_data_count_q_10_LC_14_24_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_14_24_3.LUT_INIT=16'b0101000011011000;
    LogicCell40 M_this_data_count_q_10_LC_14_24_3 (
            .in0(N__18585),
            .in1(N__18280),
            .in2(N__16206),
            .in3(N__34124),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34542),
            .ce(N__18476),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_c_0_LC_14_25_0.C_ON=1'b1;
    defparam M_this_data_count_q_cry_c_0_LC_14_25_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_c_0_LC_14_25_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 M_this_data_count_q_cry_c_0_LC_14_25_0 (
            .in0(_gnd_net_),
            .in1(N__18339),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(M_this_data_count_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_14_25_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_14_25_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_14_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_0_THRU_LUT4_0_LC_14_25_1 (
            .in0(_gnd_net_),
            .in1(N__17705),
            .in2(N__18411),
            .in3(N__16149),
            .lcout(M_this_data_count_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_0),
            .carryout(M_this_data_count_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_14_25_2.C_ON=1'b1;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_14_25_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_14_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_1_THRU_LUT4_0_LC_14_25_2 (
            .in0(_gnd_net_),
            .in1(N__18428),
            .in2(N__17805),
            .in3(N__16146),
            .lcout(M_this_data_count_q_cry_1_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_1),
            .carryout(M_this_data_count_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_14_25_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_14_25_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_14_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_2_THRU_LUT4_0_LC_14_25_3 (
            .in0(_gnd_net_),
            .in1(N__17709),
            .in2(N__18450),
            .in3(N__16143),
            .lcout(M_this_data_count_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_2),
            .carryout(M_this_data_count_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_14_25_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_14_25_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_14_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_3_THRU_LUT4_0_LC_14_25_4 (
            .in0(_gnd_net_),
            .in1(N__16947),
            .in2(N__17806),
            .in3(N__16140),
            .lcout(M_this_data_count_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_3),
            .carryout(M_this_data_count_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_14_25_5.C_ON=1'b1;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_14_25_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_14_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_4_THRU_LUT4_0_LC_14_25_5 (
            .in0(_gnd_net_),
            .in1(N__17713),
            .in2(N__16923),
            .in3(N__16137),
            .lcout(M_this_data_count_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_4),
            .carryout(M_this_data_count_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_6_LC_14_25_6.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_6_LC_14_25_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_6_LC_14_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_6_LC_14_25_6 (
            .in0(_gnd_net_),
            .in1(N__16965),
            .in2(N__17804),
            .in3(N__16134),
            .lcout(M_this_data_count_q_s_6),
            .ltout(),
            .carryin(M_this_data_count_q_cry_5),
            .carryout(M_this_data_count_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_14_25_7.C_ON=1'b1;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_14_25_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_14_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_6_THRU_LUT4_0_LC_14_25_7 (
            .in0(_gnd_net_),
            .in1(N__17714),
            .in2(N__16899),
            .in3(N__16131),
            .lcout(M_this_data_count_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_6),
            .carryout(M_this_data_count_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_7_THRU_LUT4_0_LC_14_26_0.C_ON=1'b1;
    defparam M_this_data_count_q_cry_7_THRU_LUT4_0_LC_14_26_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_7_THRU_LUT4_0_LC_14_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_7_THRU_LUT4_0_LC_14_26_0 (
            .in0(_gnd_net_),
            .in1(N__16821),
            .in2(N__17897),
            .in3(N__16128),
            .lcout(M_this_data_count_q_cry_7_THRU_CO),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(M_this_data_count_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_14_26_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_14_26_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_14_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_8_THRU_LUT4_0_LC_14_26_1 (
            .in0(_gnd_net_),
            .in1(N__17817),
            .in2(N__17454),
            .in3(N__16209),
            .lcout(M_this_data_count_q_cry_8_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_8),
            .carryout(M_this_data_count_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_10_LC_14_26_2.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_10_LC_14_26_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_10_LC_14_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_10_LC_14_26_2 (
            .in0(_gnd_net_),
            .in1(N__18386),
            .in2(N__17895),
            .in3(N__16194),
            .lcout(M_this_data_count_q_s_10),
            .ltout(),
            .carryin(M_this_data_count_q_cry_9),
            .carryout(M_this_data_count_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_14_26_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_14_26_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_14_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_10_THRU_LUT4_0_LC_14_26_3 (
            .in0(_gnd_net_),
            .in1(N__17810),
            .in2(N__18365),
            .in3(N__16191),
            .lcout(M_this_data_count_q_cry_10_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_10),
            .carryout(M_this_data_count_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_14_26_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_14_26_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_14_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_11_THRU_LUT4_0_LC_14_26_4 (
            .in0(_gnd_net_),
            .in1(N__16860),
            .in2(N__17896),
            .in3(N__16188),
            .lcout(M_this_data_count_q_cry_11_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_11),
            .carryout(M_this_data_count_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_13_LC_14_26_5.C_ON=1'b0;
    defparam M_this_data_count_q_RNO_0_13_LC_14_26_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_13_LC_14_26_5.LUT_INIT=16'b1010101001010101;
    LogicCell40 M_this_data_count_q_RNO_0_13_LC_14_26_5 (
            .in0(N__16844),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16185),
            .lcout(M_this_data_count_q_s_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_610_0_i_LC_14_26_7 .C_ON=1'b0;
    defparam \this_vga_signals.N_610_0_i_LC_14_26_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_610_0_i_LC_14_26_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \this_vga_signals.N_610_0_i_LC_14_26_7  (
            .in0(N__20600),
            .in1(N__19409),
            .in2(_gnd_net_),
            .in3(N__34109),
            .lcout(N_610_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_i_4_LC_14_27_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_4_LC_14_27_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_4_LC_14_27_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_i_4_LC_14_27_1  (
            .in0(N__32543),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18237),
            .lcout(N_87_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_i_7_LC_14_27_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_7_LC_14_27_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_i_7_LC_14_27_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_i_7_LC_14_27_7  (
            .in0(N__33657),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18238),
            .lcout(N_81_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_15_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_15_17_1 .LUT_INIT=16'b0001000100010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_15_17_1  (
            .in0(N__16611),
            .in1(N__16766),
            .in2(N__16506),
            .in3(N__16456),
            .lcout(\this_vga_signals.un4_lvisibility_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_7_LC_15_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_7_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_7_LC_15_17_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_state_q_7_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__30152),
            .in2(_gnd_net_),
            .in3(N__34118),
            .lcout(\this_ppu.M_state_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34476),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_15_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_15_17_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_15_17_4  (
            .in0(N__16765),
            .in1(N__16610),
            .in2(N__17178),
            .in3(N__17047),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_d7lto8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_15_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_15_17_5 .LUT_INIT=16'b1100110010001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_15_17_5  (
            .in0(N__16502),
            .in1(N__20110),
            .in2(N__16494),
            .in3(N__16457),
            .lcout(\this_vga_signals.M_vcounter_d8 ),
            .ltout(\this_vga_signals.M_vcounter_d8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_15_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_15_17_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__18974),
            .in2(N__16296),
            .in3(N__19119),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_0_LC_15_18_3 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_0_LC_15_18_3 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_0_LC_15_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clk.M_counter_q_0_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16281),
            .lcout(this_pixel_clk_M_counter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34482),
            .ce(),
            .sr(N__34024));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_15_19_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_15_19_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_15_19_0 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_15_19_0  (
            .in0(N__18684),
            .in1(N__16264),
            .in2(N__16229),
            .in3(N__22826),
            .lcout(\this_vga_ramdac.N_2865_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34489),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_15_19_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_15_19_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_15_19_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_15_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIDU2V1_6_LC_15_21_2.C_ON=1'b0;
    defparam M_this_state_q_RNIDU2V1_6_LC_15_21_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIDU2V1_6_LC_15_21_2.LUT_INIT=16'b1111111111110001;
    LogicCell40 M_this_state_q_RNIDU2V1_6_LC_15_21_2 (
            .in0(N__16794),
            .in1(N__16806),
            .in2(N__20496),
            .in3(N__23703),
            .lcout(),
            .ltout(dma_ac0_5_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI0F523_6_LC_15_21_3.C_ON=1'b0;
    defparam M_this_state_q_RNI0F523_6_LC_15_21_3.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI0F523_6_LC_15_21_3.LUT_INIT=16'b0000110000000000;
    LogicCell40 M_this_state_q_RNI0F523_6_LC_15_21_3 (
            .in0(_gnd_net_),
            .in1(N__16800),
            .in2(N__16212),
            .in3(N__19317),
            .lcout(dma_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_tr27_i_o3_LC_15_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_tr27_i_o3_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_tr27_i_o3_LC_15_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_tr27_i_o3_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__18306),
            .in2(_gnd_net_),
            .in3(N__35793),
            .lcout(N_160_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIOE1S_11_LC_15_22_0.C_ON=1'b0;
    defparam M_this_state_q_RNIOE1S_11_LC_15_22_0.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIOE1S_11_LC_15_22_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_state_q_RNIOE1S_11_LC_15_22_0 (
            .in0(N__19691),
            .in1(N__18304),
            .in2(N__24965),
            .in3(N__20342),
            .lcout(M_this_state_q_RNIOE1SZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un20_i_a2_x_3_LC_15_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un20_i_a2_x_3_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un20_i_a2_x_3_LC_15_22_1 .LUT_INIT=16'b0000000100000001;
    LogicCell40 \this_vga_signals.un20_i_a2_x_3_LC_15_22_1  (
            .in0(N__18305),
            .in1(N__28120),
            .in2(N__23750),
            .in3(_gnd_net_),
            .lcout(un20_i_a2_x_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIG01L_12_LC_15_22_6.C_ON=1'b0;
    defparam M_this_state_q_RNIG01L_12_LC_15_22_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIG01L_12_LC_15_22_6.LUT_INIT=16'b0000000000010001;
    LogicCell40 M_this_state_q_RNIG01L_12_LC_15_22_6 (
            .in0(N__35579),
            .in1(N__28119),
            .in2(_gnd_net_),
            .in3(N__20410),
            .lcout(M_this_state_q_RNIG01LZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_326_i_i_a2_LC_15_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.N_326_i_i_a2_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_326_i_i_a2_LC_15_23_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.N_326_i_i_a2_LC_15_23_7  (
            .in0(_gnd_net_),
            .in1(N__19313),
            .in2(_gnd_net_),
            .in3(N__20492),
            .lcout(N_278),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_419_i_i_0_1_LC_15_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.N_419_i_i_0_1_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_419_i_i_0_1_LC_15_24_1 .LUT_INIT=16'b0000101000110011;
    LogicCell40 \this_vga_signals.N_419_i_i_0_1_LC_15_24_1  (
            .in0(N__19872),
            .in1(N__19395),
            .in2(N__19436),
            .in3(N__20416),
            .lcout(),
            .ltout(\this_vga_signals.N_419_i_i_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_qe_0_i_LC_15_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_qe_0_i_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_qe_0_i_LC_15_24_2 .LUT_INIT=16'b1111111110110000;
    LogicCell40 \this_vga_signals.M_this_data_count_qe_0_i_LC_15_24_2  (
            .in0(N__19396),
            .in1(N__20512),
            .in2(N__16788),
            .in3(N__34114),
            .lcout(M_this_data_count_qe_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_a3_0_9_LC_15_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_a3_0_9_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_a3_0_9_LC_15_24_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_a3_0_9_LC_15_24_4  (
            .in0(N__33487),
            .in1(N__20415),
            .in2(N__34770),
            .in3(N__19871),
            .lcout(N_212),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_6_LC_15_25_0.C_ON=1'b0;
    defparam M_this_data_count_q_6_LC_15_25_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_15_25_0.LUT_INIT=16'b0010001011100010;
    LogicCell40 M_this_data_count_q_6_LC_15_25_0 (
            .in0(N__16785),
            .in1(N__18568),
            .in2(N__19569),
            .in3(N__34123),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34543),
            .ce(N__18477),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d55_9_LC_15_25_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d55_9_LC_15_25_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d55_9_LC_15_25_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_d55_9_LC_15_25_1  (
            .in0(N__16964),
            .in1(N__16918),
            .in2(N__16898),
            .in3(N__16945),
            .lcout(\this_vga_signals.M_this_state_d55Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_4_LC_15_25_2.C_ON=1'b0;
    defparam M_this_data_count_q_4_LC_15_25_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_15_25_2.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_4_LC_15_25_2 (
            .in0(N__16946),
            .in1(N__16953),
            .in2(_gnd_net_),
            .in3(N__18566),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34543),
            .ce(N__18477),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_5_LC_15_25_3.C_ON=1'b0;
    defparam M_this_data_count_q_5_LC_15_25_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_15_25_3.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_5_LC_15_25_3 (
            .in0(N__16932),
            .in1(N__18565),
            .in2(_gnd_net_),
            .in3(N__16919),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34543),
            .ce(N__18477),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_7_LC_15_25_4.C_ON=1'b0;
    defparam M_this_data_count_q_7_LC_15_25_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_15_25_4.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_7_LC_15_25_4 (
            .in0(N__16905),
            .in1(N__18567),
            .in2(_gnd_net_),
            .in3(N__16894),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34543),
            .ce(N__18477),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_3_LC_15_25_5.C_ON=1'b0;
    defparam M_this_data_count_q_3_LC_15_25_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_15_25_5.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_3_LC_15_25_5 (
            .in0(N__16878),
            .in1(N__18564),
            .in2(_gnd_net_),
            .in3(N__18449),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34543),
            .ce(N__18477),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_11_LC_15_26_2.C_ON=1'b0;
    defparam M_this_data_count_q_11_LC_15_26_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_15_26_2.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_11_LC_15_26_2 (
            .in0(N__18366),
            .in1(N__18558),
            .in2(_gnd_net_),
            .in3(N__16872),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34549),
            .ce(N__18491),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_12_LC_15_26_3.C_ON=1'b0;
    defparam M_this_data_count_q_12_LC_15_26_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_15_26_3.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_12_LC_15_26_3 (
            .in0(N__18559),
            .in1(N__16866),
            .in2(_gnd_net_),
            .in3(N__16859),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34549),
            .ce(N__18491),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d55_8_LC_15_26_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d55_8_LC_15_26_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d55_8_LC_15_26_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_d55_8_LC_15_26_4  (
            .in0(N__16858),
            .in1(N__17449),
            .in2(N__16845),
            .in3(N__16819),
            .lcout(\this_vga_signals.M_this_state_d55Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_8_LC_15_26_5.C_ON=1'b0;
    defparam M_this_data_count_q_8_LC_15_26_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_15_26_5.LUT_INIT=16'b0000100100001001;
    LogicCell40 M_this_data_count_q_8_LC_15_26_5 (
            .in0(N__16820),
            .in1(N__16827),
            .in2(N__18579),
            .in3(_gnd_net_),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34549),
            .ce(N__18491),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_2_LC_15_26_7.C_ON=1'b0;
    defparam M_this_data_count_q_2_LC_15_26_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_15_26_7.LUT_INIT=16'b0101000000000101;
    LogicCell40 M_this_data_count_q_2_LC_15_26_7 (
            .in0(N__18560),
            .in1(_gnd_net_),
            .in2(N__17469),
            .in3(N__18429),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34549),
            .ce(N__18491),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_9_LC_15_27_0.C_ON=1'b0;
    defparam M_this_data_count_q_9_LC_15_27_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_15_27_0.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_9_LC_15_27_0 (
            .in0(N__17460),
            .in1(N__18569),
            .in2(_gnd_net_),
            .in3(N__17453),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34557),
            .ce(N__18498),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI43UU_1_6_LC_16_15_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI43UU_1_6_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI43UU_1_6_LC_16_15_4 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \this_ppu.M_state_q_RNI43UU_1_6_LC_16_15_4  (
            .in0(N__17433),
            .in1(N__29978),
            .in2(N__30145),
            .in3(N__31137),
            .lcout(M_this_ppu_sprites_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_LC_16_17_0 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_LC_16_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.line_clk.M_last_q_LC_16_17_0 .LUT_INIT=16'b1011000011010000;
    LogicCell40 \this_ppu.line_clk.M_last_q_LC_16_17_0  (
            .in0(N__17190),
            .in1(N__17177),
            .in2(N__20004),
            .in3(N__17048),
            .lcout(\this_ppu.M_last_q ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34473),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIKM001_1_LC_16_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIKM001_1_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIKM001_1_LC_16_18_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_ppu.M_count_q_RNIKM001_1_LC_16_18_1  (
            .in0(N__19150),
            .in1(N__18057),
            .in2(N__19227),
            .in3(N__18633),
            .lcout(\this_ppu.M_count_d_0_sqmuxa_1_7 ),
            .ltout(\this_ppu.M_count_d_0_sqmuxa_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_7_LC_16_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_7_LC_16_18_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_7_LC_16_18_2 .LUT_INIT=16'b0101111101001100;
    LogicCell40 \this_ppu.M_count_q_7_LC_16_18_2  (
            .in0(N__25931),
            .in1(N__17496),
            .in2(N__17193),
            .in3(N__28642),
            .lcout(\this_ppu.M_count_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34475),
            .ce(),
            .sr(N__34021));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICHRV3_8_LC_16_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICHRV3_8_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICHRV3_8_LC_16_18_4 .LUT_INIT=16'b1011000011010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICHRV3_8_LC_16_18_4  (
            .in0(N__17189),
            .in1(N__17176),
            .in2(N__20000),
            .in3(N__17073),
            .lcout(M_this_vga_signals_line_clk_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_19_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__19191),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\this_ppu.un1_M_count_q_1_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_19_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__19151),
            .in2(N__17602),
            .in3(N__16968),
            .lcout(\this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_0_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_19_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__17550),
            .in2(N__18075),
            .in3(N__18033),
            .lcout(\this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_1_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_19_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__19219),
            .in2(N__17603),
            .in3(N__18030),
            .lcout(\this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_2_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_19_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__17554),
            .in2(N__18120),
            .in3(N__18027),
            .lcout(\this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_3_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_19_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__18137),
            .in2(N__17604),
            .in3(N__18024),
            .lcout(\this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_4_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_19_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__17558),
            .in2(N__18102),
            .in3(N__17502),
            .lcout(\this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_5_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_7_LC_16_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_16_19_7 .LUT_INIT=16'b1100110000110110;
    LogicCell40 \this_ppu.M_count_q_RNO_0_7_LC_16_19_7  (
            .in0(N__25925),
            .in1(N__18645),
            .in2(N__28668),
            .in3(N__17499),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_5_LC_16_20_0 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_5_LC_16_20_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_5_LC_16_20_0 .LUT_INIT=16'b1010000010000010;
    LogicCell40 \this_ppu.M_count_q_5_LC_16_20_0  (
            .in0(N__19253),
            .in1(N__17490),
            .in2(N__18138),
            .in3(N__19288),
            .lcout(\this_ppu.M_count_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34486),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_6_LC_16_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_6_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_6_LC_16_20_2 .LUT_INIT=16'b1010000010000010;
    LogicCell40 \this_ppu.M_count_q_6_LC_16_20_2  (
            .in0(N__19254),
            .in1(N__17484),
            .in2(N__18098),
            .in3(N__19289),
            .lcout(\this_ppu.M_count_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34486),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_4_LC_16_20_4 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_4_LC_16_20_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_4_LC_16_20_4 .LUT_INIT=16'b1010100000000010;
    LogicCell40 \this_ppu.M_count_q_4_LC_16_20_4  (
            .in0(N__19252),
            .in1(N__17478),
            .in2(N__19290),
            .in3(N__18116),
            .lcout(\this_ppu.M_count_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34486),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_2_LC_16_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_2_LC_16_20_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_2_LC_16_20_5 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_2_LC_16_20_5  (
            .in0(N__18071),
            .in1(N__19284),
            .in2(N__18147),
            .in3(N__19251),
            .lcout(\this_ppu.M_count_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34486),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIDE0G_2_LC_16_20_6 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIDE0G_2_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIDE0G_2_LC_16_20_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_count_q_RNIDE0G_2_LC_16_20_6  (
            .in0(N__18133),
            .in1(N__18115),
            .in2(N__18097),
            .in3(N__18070),
            .lcout(\this_ppu.M_count_d_1_sqmuxa_1_i_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_9_LC_16_20_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_9_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_9_LC_16_20_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_9_LC_16_20_7  (
            .in0(N__21023),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18666),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34486),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_2_LC_16_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_2_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_2_LC_16_21_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_i_o3_0_2_LC_16_21_0  (
            .in0(N__21678),
            .in1(N__21727),
            .in2(_gnd_net_),
            .in3(N__21634),
            .lcout(N_465_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_10_LC_16_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_10_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_10_LC_16_21_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_i_o3_0_10_LC_16_21_1  (
            .in0(N__21635),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19344),
            .lcout(this_vga_signals_M_this_state_q_ns_i_o3_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_16_21_2 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_16_21_2 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_16_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18048),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34497),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_6_LC_16_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_6_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_6_LC_16_21_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_6_LC_16_21_4  (
            .in0(N__26373),
            .in1(N__21213),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_8_LC_16_22_0.C_ON=1'b0;
    defparam M_this_state_q_8_LC_16_22_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_8_LC_16_22_0.LUT_INIT=16'b0000110000001000;
    LogicCell40 M_this_state_q_8_LC_16_22_0 (
            .in0(N__20865),
            .in1(N__23702),
            .in2(N__20937),
            .in3(N__20809),
            .lcout(M_this_state_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34505),
            .ce(),
            .sr(N__34012));
    defparam \this_vga_signals.un20_i_a2_sx_3_LC_16_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un20_i_a2_sx_3_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un20_i_a2_sx_3_LC_16_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \this_vga_signals.un20_i_a2_sx_3_LC_16_22_1  (
            .in0(N__18302),
            .in1(N__19338),
            .in2(N__19692),
            .in3(N__23728),
            .lcout(),
            .ltout(\this_vga_signals.un20_i_a2_sxZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un20_i_a2_3_LC_16_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un20_i_a2_3_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un20_i_a2_3_LC_16_22_2 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \this_vga_signals.un20_i_a2_3_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18036),
            .in3(N__28118),
            .lcout(),
            .ltout(\this_vga_signals.N_322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_11_0_i_LC_16_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_11_0_i_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_11_0_i_LC_16_22_3 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_11_0_i_LC_16_22_3  (
            .in0(N__19296),
            .in1(N__23729),
            .in2(N__18318),
            .in3(N__35713),
            .lcout(un1_M_this_state_q_11_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_10_LC_16_22_4.C_ON=1'b0;
    defparam M_this_state_q_10_LC_16_22_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_10_LC_16_22_4.LUT_INIT=16'b0101010100010000;
    LogicCell40 M_this_state_q_10_LC_16_22_4 (
            .in0(N__35714),
            .in1(N__20610),
            .in2(N__18315),
            .in3(N__18303),
            .lcout(M_this_state_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34505),
            .ce(),
            .sr(N__34012));
    defparam M_this_state_q_2_LC_16_23_0.C_ON=1'b0;
    defparam M_this_state_q_2_LC_16_23_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_16_23_0.LUT_INIT=16'b0000000011111000;
    LogicCell40 M_this_state_q_2_LC_16_23_0 (
            .in0(N__18627),
            .in1(N__28567),
            .in2(N__24995),
            .in3(N__35812),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34513),
            .ce(),
            .sr(N__34011));
    defparam M_this_substate_q_LC_16_23_1.C_ON=1'b0;
    defparam M_this_substate_q_LC_16_23_1.SEQ_MODE=4'b1000;
    defparam M_this_substate_q_LC_16_23_1.LUT_INIT=16'b1100000011101010;
    LogicCell40 M_this_substate_q_LC_16_23_1 (
            .in0(N__19545),
            .in1(N__19526),
            .in2(N__18615),
            .in3(N__24228),
            .lcout(M_this_substate_qZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34513),
            .ce(),
            .sr(N__34011));
    defparam M_this_state_q_9_LC_16_23_2.C_ON=1'b0;
    defparam M_this_state_q_9_LC_16_23_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_9_LC_16_23_2.LUT_INIT=16'b1111111011111010;
    LogicCell40 M_this_state_q_9_LC_16_23_2 (
            .in0(N__18281),
            .in1(N__20519),
            .in2(N__18251),
            .in3(N__19343),
            .lcout(M_this_state_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34513),
            .ce(),
            .sr(N__34011));
    defparam M_this_state_q_11_LC_16_23_4.C_ON=1'b0;
    defparam M_this_state_q_11_LC_16_23_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_11_LC_16_23_4.LUT_INIT=16'b1111110011111110;
    LogicCell40 M_this_state_q_11_LC_16_23_4 (
            .in0(N__19668),
            .in1(N__19562),
            .in2(N__35248),
            .in3(N__21650),
            .lcout(M_this_state_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34513),
            .ce(),
            .sr(N__34011));
    defparam M_this_state_q_5_LC_16_23_5.C_ON=1'b0;
    defparam M_this_state_q_5_LC_16_23_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_16_23_5.LUT_INIT=16'b1101010111000000;
    LogicCell40 M_this_state_q_5_LC_16_23_5 (
            .in0(N__35810),
            .in1(N__19361),
            .in2(N__26670),
            .in3(N__20420),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34513),
            .ce(),
            .sr(N__34011));
    defparam M_this_state_q_1_LC_16_23_6.C_ON=1'b0;
    defparam M_this_state_q_1_LC_16_23_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_16_23_6.LUT_INIT=16'b1010000011101100;
    LogicCell40 M_this_state_q_1_LC_16_23_6 (
            .in0(N__19360),
            .in1(N__26318),
            .in2(N__19527),
            .in3(N__35811),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34513),
            .ce(),
            .sr(N__34011));
    defparam M_this_state_q_12_LC_16_23_7.C_ON=1'b0;
    defparam M_this_state_q_12_LC_16_23_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_12_LC_16_23_7.LUT_INIT=16'b0101010101000000;
    LogicCell40 M_this_state_q_12_LC_16_23_7 (
            .in0(N__35809),
            .in1(N__19667),
            .in2(N__21654),
            .in3(N__28126),
            .lcout(M_this_state_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34513),
            .ce(),
            .sr(N__34011));
    defparam M_this_state_q_RNO_0_2_LC_16_24_0.C_ON=1'b0;
    defparam M_this_state_q_RNO_0_2_LC_16_24_0.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_0_2_LC_16_24_0.LUT_INIT=16'b0000100000000000;
    LogicCell40 M_this_state_q_RNO_0_2_LC_16_24_0 (
            .in0(N__26725),
            .in1(N__19543),
            .in2(N__28415),
            .in3(N__18610),
            .lcout(M_this_state_qc_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_1_4_LC_16_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_1_4_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_1_4_LC_16_24_2 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_1_4_LC_16_24_2  (
            .in0(N__26726),
            .in1(_gnd_net_),
            .in2(N__28416),
            .in3(N__18611),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_q_ns_0_i_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_16_24_3.C_ON=1'b0;
    defparam M_this_state_q_4_LC_16_24_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_16_24_3.LUT_INIT=16'b0101110100001100;
    LogicCell40 M_this_state_q_4_LC_16_24_3 (
            .in0(N__35813),
            .in1(N__28579),
            .in2(N__18618),
            .in3(N__35578),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34524),
            .ce(),
            .sr(N__34010));
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_1_LC_16_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_1_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_1_LC_16_24_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o2_1_LC_16_24_4  (
            .in0(N__26727),
            .in1(N__28414),
            .in2(N__28584),
            .in3(N__18609),
            .lcout(N_484_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_419_i_i_0_a2_LC_16_25_3 .C_ON=1'b0;
    defparam \this_vga_signals.N_419_i_i_0_a2_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_419_i_i_0_a2_LC_16_25_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.N_419_i_i_0_a2_LC_16_25_3  (
            .in0(N__21649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20579),
            .lcout(\this_vga_signals.N_279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_0_LC_16_25_4.C_ON=1'b0;
    defparam M_this_data_count_q_0_LC_16_25_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_16_25_4.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_0_LC_16_25_4 (
            .in0(_gnd_net_),
            .in1(N__18587),
            .in2(_gnd_net_),
            .in3(N__18338),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34533),
            .ce(N__18484),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_1_LC_16_25_7.C_ON=1'b0;
    defparam M_this_data_count_q_1_LC_16_25_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_16_25_7.LUT_INIT=16'b0101000000000101;
    LogicCell40 M_this_data_count_q_1_LC_16_25_7 (
            .in0(N__18588),
            .in1(_gnd_net_),
            .in2(N__18510),
            .in3(N__18407),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34533),
            .ce(N__18484),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d55_6_LC_16_26_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d55_6_LC_16_26_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d55_6_LC_16_26_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_this_state_d55_6_LC_16_26_1  (
            .in0(_gnd_net_),
            .in1(N__18445),
            .in2(_gnd_net_),
            .in3(N__18427),
            .lcout(\this_vga_signals.M_this_state_d55Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d55_7_LC_16_26_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d55_7_LC_16_26_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d55_7_LC_16_26_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_d55_7_LC_16_26_5  (
            .in0(N__18403),
            .in1(N__18387),
            .in2(N__18364),
            .in3(N__18334),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_d55Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d55_LC_16_26_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d55_LC_16_26_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d55_LC_16_26_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_state_d55_LC_16_26_6  (
            .in0(N__18906),
            .in1(N__18900),
            .in2(N__18894),
            .in3(N__18891),
            .lcout(M_this_state_d55),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_17_16_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_17_16_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_17_16_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__20988),
            .in2(_gnd_net_),
            .in3(N__21042),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34474),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_17_16_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_17_16_6 .LUT_INIT=16'b0010001110010111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_17_16_6  (
            .in0(N__18885),
            .in1(N__18831),
            .in2(N__18789),
            .in3(N__18732),
            .lcout(\this_vga_ramdac.m16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_6_LC_17_17_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_6_LC_17_17_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_6_LC_17_17_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_6_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__20990),
            .in2(_gnd_net_),
            .in3(N__18672),
            .lcout(\this_reset_cond.M_stage_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34477),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_5_LC_17_17_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_5_LC_17_17_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_5_LC_17_17_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_5_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__20989),
            .in2(_gnd_net_),
            .in3(N__19740),
            .lcout(\this_reset_cond.M_stage_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34477),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_8_LC_17_17_5 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_8_LC_17_17_5 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_8_LC_17_17_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_8_LC_17_17_5  (
            .in0(N__20992),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18651),
            .lcout(\this_reset_cond.M_stage_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34477),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_7_LC_17_17_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_7_LC_17_17_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_7_LC_17_17_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_7_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__20991),
            .in2(_gnd_net_),
            .in3(N__18657),
            .lcout(\this_reset_cond.M_stage_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34477),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIL508_7_LC_17_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIL508_7_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIL508_7_LC_17_18_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_count_q_RNIL508_7_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__18644),
            .in2(_gnd_net_),
            .in3(N__19189),
            .lcout(\this_ppu.M_count_d_1_sqmuxa_1_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_0_LC_17_18_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_0_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_0_LC_17_18_3 .LUT_INIT=16'b1101000011111111;
    LogicCell40 \this_ppu.M_state_q_0_LC_17_18_3  (
            .in0(N__29358),
            .in1(N__29403),
            .in2(N__29471),
            .in3(N__18921),
            .lcout(\this_ppu.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34483),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI4GQN4_0_LC_17_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI4GQN4_0_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI4GQN4_0_LC_17_18_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_ppu.M_state_q_RNI4GQN4_0_LC_17_18_6  (
            .in0(N__29402),
            .in1(N__29456),
            .in2(_gnd_net_),
            .in3(N__29357),
            .lcout(\this_ppu.N_132_0 ),
            .ltout(\this_ppu.N_132_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_0_LC_17_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_0_LC_17_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_0_LC_17_18_7 .LUT_INIT=16'b0000011000000000;
    LogicCell40 \this_ppu.M_count_q_0_LC_17_18_7  (
            .in0(N__19190),
            .in1(N__25930),
            .in2(N__19194),
            .in3(N__18920),
            .lcout(\this_ppu.M_count_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34483),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNIL33N6_1_LC_17_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNIL33N6_1_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNIL33N6_1_LC_17_19_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNIL33N6_1_LC_17_19_0  (
            .in0(N__19133),
            .in1(N__19176),
            .in2(_gnd_net_),
            .in3(N__20147),
            .lcout(\this_vga_signals.un1_M_hcounter_d7_1_0 ),
            .ltout(\this_vga_signals.un1_M_hcounter_d7_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_0_LC_17_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_0_LC_17_19_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_0_LC_17_19_1 .LUT_INIT=16'b0010011000101010;
    LogicCell40 \this_vga_signals.M_lcounter_q_0_LC_17_19_1  (
            .in0(N__20133),
            .in1(N__19054),
            .in2(N__19164),
            .in3(N__19134),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_1_LC_17_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_1_LC_17_19_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_1_LC_17_19_2 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_1_LC_17_19_2  (
            .in0(N__19152),
            .in1(N__19283),
            .in2(N__19161),
            .in3(N__19250),
            .lcout(\this_ppu.M_count_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI01PG1_0_1_LC_17_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI01PG1_0_1_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI01PG1_0_1_LC_17_19_3 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_ppu.M_state_q_RNI01PG1_0_1_LC_17_19_3  (
            .in0(N__25846),
            .in1(N__25921),
            .in2(_gnd_net_),
            .in3(N__34106),
            .lcout(\this_ppu.N_1157_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_17_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_17_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_1_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__20132),
            .in2(_gnd_net_),
            .in3(N__19132),
            .lcout(),
            .ltout(\this_vga_signals.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_1_LC_17_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_1_LC_17_19_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_1_LC_17_19_6 .LUT_INIT=16'b0101011100100000;
    LogicCell40 \this_vga_signals.M_lcounter_q_1_LC_17_19_6  (
            .in0(N__19053),
            .in1(N__18930),
            .in2(N__18924),
            .in3(N__20148),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34490),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI4HJ86_0_LC_17_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI4HJ86_0_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI4HJ86_0_LC_17_20_5 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \this_ppu.M_state_q_RNI4HJ86_0_LC_17_20_5  (
            .in0(N__29472),
            .in1(N__18919),
            .in2(N__29434),
            .in3(N__29370),
            .lcout(\this_ppu.N_1157_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI4L615_0_LC_17_20_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI4L615_0_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI4L615_0_LC_17_20_6 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \this_ppu.M_state_q_RNI4L615_0_LC_17_20_6  (
            .in0(N__29371),
            .in1(N__29427),
            .in2(N__25932),
            .in3(N__29473),
            .lcout(\this_ppu.un16_0 ),
            .ltout(\this_ppu.un16_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_3_LC_17_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_3_LC_17_20_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_3_LC_17_20_7 .LUT_INIT=16'b1100100100000000;
    LogicCell40 \this_ppu.M_count_q_3_LC_17_20_7  (
            .in0(N__19263),
            .in1(N__19220),
            .in2(N__19257),
            .in3(N__19249),
            .lcout(\this_ppu.M_count_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34500),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_1_LC_17_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_1_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_1_LC_17_21_1 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_1_LC_17_21_1  (
            .in0(N__26138),
            .in1(N__24984),
            .in2(N__32971),
            .in3(N__35755),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_start_data_delay_out_m_0_LC_17_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_start_data_delay_out_m_0_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_start_data_delay_out_m_0_LC_17_21_2 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \this_vga_signals.M_this_start_data_delay_out_m_0_LC_17_21_2  (
            .in0(N__23690),
            .in1(N__20924),
            .in2(N__20893),
            .in3(N__20801),
            .lcout(\this_vga_signals.M_this_state_q_ns_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_0_LC_17_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_0_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o2_0_LC_17_21_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o2_0_LC_17_21_3  (
            .in0(N__20800),
            .in1(_gnd_net_),
            .in2(N__20934),
            .in3(N__20885),
            .lcout(N_459_0),
            .ltout(N_459_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_0_0_LC_17_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_0_0_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_0_0_LC_17_21_4 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o3_0_0_LC_17_21_4  (
            .in0(N__21728),
            .in1(_gnd_net_),
            .in2(N__19200),
            .in3(_gnd_net_),
            .lcout(N_462_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_17_21_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_17_21_5 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_17_21_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_17_21_5  (
            .in0(N__20802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20881),
            .lcout(this_start_data_delay_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34509),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_LC_17_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_LC_17_21_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o3_1_LC_17_21_6  (
            .in0(N__20886),
            .in1(N__20920),
            .in2(_gnd_net_),
            .in3(N__20799),
            .lcout(N_458_0),
            .ltout(N_458_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_419_i_i_0_o2_LC_17_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.N_419_i_i_0_o2_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_419_i_i_0_o2_LC_17_21_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vga_signals.N_419_i_i_0_o2_LC_17_21_7  (
            .in0(N__32954),
            .in1(N__20552),
            .in2(N__19197),
            .in3(N__33670),
            .lcout(\this_vga_signals.N_169_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_2_0_LC_17_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_2_0_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_2_0_LC_17_22_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o3_2_0_LC_17_22_0  (
            .in0(N__20334),
            .in1(N__24961),
            .in2(N__35609),
            .in3(N__26292),
            .lcout(),
            .ltout(N_496_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_1_0_LC_17_22_1.C_ON=1'b0;
    defparam M_this_state_q_RNO_1_0_LC_17_22_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_1_0_LC_17_22_1.LUT_INIT=16'b0111010111110101;
    LogicCell40 M_this_state_q_RNO_1_0_LC_17_22_1 (
            .in0(N__35716),
            .in1(N__19440),
            .in2(N__19413),
            .in3(N__20414),
            .lcout(),
            .ltout(M_this_state_qsr_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNO_0_0_LC_17_22_2.C_ON=1'b0;
    defparam M_this_state_q_RNO_0_0_LC_17_22_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNO_0_0_LC_17_22_2.LUT_INIT=16'b0100000001010000;
    LogicCell40 M_this_state_q_RNO_0_0_LC_17_22_2 (
            .in0(N__19659),
            .in1(N__19410),
            .in2(N__19380),
            .in3(N__20609),
            .lcout(),
            .ltout(M_this_state_qsr_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_0_LC_17_22_3.C_ON=1'b0;
    defparam M_this_state_q_0_LC_17_22_3.SEQ_MODE=4'b1001;
    defparam M_this_state_q_0_LC_17_22_3.LUT_INIT=16'b1101111100001111;
    LogicCell40 M_this_state_q_0_LC_17_22_3 (
            .in0(N__19377),
            .in1(N__21744),
            .in2(N__19371),
            .in3(N__21679),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34518),
            .ce(),
            .sr(N__34014));
    defparam M_this_state_q_3_LC_17_22_4.C_ON=1'b0;
    defparam M_this_state_q_3_LC_17_22_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_17_22_4.LUT_INIT=16'b0000000011101010;
    LogicCell40 M_this_state_q_3_LC_17_22_4 (
            .in0(N__20335),
            .in1(N__19368),
            .in2(N__26760),
            .in3(N__35717),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34518),
            .ce(),
            .sr(N__34014));
    defparam \this_vga_signals.M_this_external_address_d_0_sqmuxa_1_3_LC_17_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_0_sqmuxa_1_3_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_0_sqmuxa_1_3_LC_17_22_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_this_external_address_d_0_sqmuxa_1_3_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(N__23673),
            .in2(_gnd_net_),
            .in3(N__20333),
            .lcout(\this_vga_signals.N_159_0 ),
            .ltout(\this_vga_signals.N_159_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_12_0_m2_LC_17_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_12_0_m2_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_12_0_m2_LC_17_22_6 .LUT_INIT=16'b1110111111100000;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_12_0_m2_LC_17_22_6  (
            .in0(N__24933),
            .in1(N__26291),
            .in2(N__19347),
            .in3(N__35715),
            .lcout(\this_vga_signals.N_166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un22_i_a2_0_o2_LC_17_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.un22_i_a2_0_o2_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un22_i_a2_0_o2_LC_17_23_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.un22_i_a2_0_o2_LC_17_23_0  (
            .in0(_gnd_net_),
            .in1(N__19689),
            .in2(_gnd_net_),
            .in3(N__19339),
            .lcout(N_168_0),
            .ltout(N_168_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_d_0_sqmuxa_1_2_LC_17_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_d_0_sqmuxa_1_2_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_d_0_sqmuxa_1_2_LC_17_23_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_d_0_sqmuxa_1_2_LC_17_23_1  (
            .in0(N__20409),
            .in1(N__26290),
            .in2(N__19299),
            .in3(N__20270),
            .lcout(\this_vga_signals.M_this_external_address_d_0_sqmuxa_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_11_LC_17_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_11_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_11_LC_17_23_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o3_1_11_LC_17_23_6  (
            .in0(_gnd_net_),
            .in1(N__20607),
            .in2(_gnd_net_),
            .in3(N__19690),
            .lcout(N_456_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_0_0_LC_17_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_0_0_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_0_0_LC_17_23_7 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a3_0_0_LC_17_23_7  (
            .in0(N__32916),
            .in1(N__33672),
            .in2(N__20553),
            .in3(N__24199),
            .lcout(N_500),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_0_LC_17_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_0_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_0_LC_17_24_0 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_0_LC_17_24_0  (
            .in0(N__33800),
            .in1(N__27399),
            .in2(N__32598),
            .in3(N__27350),
            .lcout(M_this_sprites_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d_2_sqmuxa_LC_17_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d_2_sqmuxa_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d_2_sqmuxa_LC_17_24_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_this_state_d_2_sqmuxa_LC_17_24_4  (
            .in0(N__24218),
            .in1(N__34740),
            .in2(_gnd_net_),
            .in3(N__24200),
            .lcout(M_this_state_d_2_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_0_0_1_LC_17_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_0_0_1_LC_17_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_0_0_1_LC_17_24_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a3_0_0_1_LC_17_24_5  (
            .in0(N__28407),
            .in1(N__26708),
            .in2(N__28583),
            .in3(N__19544),
            .lcout(this_vga_signals_M_this_state_q_ns_0_a3_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_2_LC_17_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_2_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_2_LC_17_24_6 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_2_LC_17_24_6  (
            .in0(N__35781),
            .in1(N__22133),
            .in2(N__33491),
            .in3(N__24960),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3_0_LC_17_25_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3_0_LC_17_25_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3_0_LC_17_25_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3_0_LC_17_25_2  (
            .in0(N__33799),
            .in1(N__32799),
            .in2(N__32409),
            .in3(N__32588),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_o3_1_0_o2_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_18_15_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_18_15_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_18_15_1  (
            .in0(N__19512),
            .in1(N__19491),
            .in2(_gnd_net_),
            .in3(N__30458),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_18_15_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_18_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_18_15_2  (
            .in0(N__30455),
            .in1(N__19476),
            .in2(_gnd_net_),
            .in3(N__19455),
            .lcout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_18_15_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_18_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_18_15_3  (
            .in0(N__19851),
            .in1(N__19833),
            .in2(_gnd_net_),
            .in3(N__30457),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_18_15_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_18_15_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_18_15_4  (
            .in0(N__30456),
            .in1(N__19815),
            .in2(_gnd_net_),
            .in3(N__19797),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_18_15_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_18_15_5 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_18_15_5  (
            .in0(N__28999),
            .in1(N__24588),
            .in2(N__19776),
            .in3(N__19773),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_18_15_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_18_15_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_18_15_6  (
            .in0(N__24589),
            .in1(N__19767),
            .in2(N__19761),
            .in3(N__19758),
            .lcout(M_this_ppu_vram_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_18_16_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_18_16_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_18_16_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__21021),
            .in2(_gnd_net_),
            .in3(N__19752),
            .lcout(\this_reset_cond.M_stage_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34478),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_4_LC_18_16_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_4_LC_18_16_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_4_LC_18_16_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_4_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__21022),
            .in2(_gnd_net_),
            .in3(N__19746),
            .lcout(\this_reset_cond.M_stage_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34478),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_18_17_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_18_17_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_18_17_1  (
            .in0(N__30418),
            .in1(N__19734),
            .in2(_gnd_net_),
            .in3(N__19716),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_18_17_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_18_17_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_18_17_2  (
            .in0(N__29003),
            .in1(N__24593),
            .in2(N__19695),
            .in3(N__25038),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_18_17_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_18_17_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_18_17_3  (
            .in0(N__24594),
            .in1(N__20154),
            .in2(N__20223),
            .in3(N__20631),
            .lcout(M_this_ppu_vram_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_13_LC_18_17_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_13_LC_18_17_4 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_13_LC_18_17_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \this_sprites_ram.mem_radreg_13_LC_18_17_4  (
            .in0(N__31002),
            .in1(N__30108),
            .in2(N__20220),
            .in3(N__29999),
            .lcout(\this_sprites_ram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34484),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_18_17_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_18_17_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_18_17_7  (
            .in0(N__30419),
            .in1(N__20193),
            .in2(_gnd_net_),
            .in3(N__20172),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_7_LC_18_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_7_LC_18_18_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_7_LC_18_18_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_haddress_q_7_LC_18_18_0  (
            .in0(N__20622),
            .in1(N__25135),
            .in2(N__25258),
            .in3(N__25185),
            .lcout(M_this_ppu_map_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34491),
            .ce(),
            .sr(N__23129));
    defparam \this_ppu.M_haddress_q_5_LC_18_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_5_LC_18_18_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_5_LC_18_18_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_haddress_q_5_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__25243),
            .in2(_gnd_net_),
            .in3(N__20620),
            .lcout(M_this_ppu_map_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34491),
            .ce(),
            .sr(N__23129));
    defparam \this_ppu.M_haddress_q_6_LC_18_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_6_LC_18_18_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_6_LC_18_18_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \this_ppu.M_haddress_q_6_LC_18_18_2  (
            .in0(N__20621),
            .in1(_gnd_net_),
            .in2(N__25257),
            .in3(N__25184),
            .lcout(M_this_ppu_map_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34491),
            .ce(),
            .sr(N__23129));
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_18_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_18_18_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_18_18_4  (
            .in0(N__20146),
            .in1(N__20131),
            .in2(_gnd_net_),
            .in3(N__20109),
            .lcout(\this_vga_signals.line_clk_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_3_LC_18_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_3_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_3_LC_18_19_6 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_3_LC_18_19_6  (
            .in0(N__32800),
            .in1(N__27404),
            .in2(N__33658),
            .in3(N__27368),
            .lcout(M_this_sprites_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_a3_0_6_LC_18_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_a3_0_6_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_a3_0_6_LC_18_21_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_a3_0_6_LC_18_21_0  (
            .in0(N__33471),
            .in1(N__20433),
            .in2(N__34705),
            .in3(N__19862),
            .lcout(N_210),
            .ltout(N_210_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_12_0_o3_LC_18_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_12_0_o3_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_12_0_o3_LC_18_21_1 .LUT_INIT=16'b0000101000001111;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_12_0_o3_LC_18_21_1  (
            .in0(N__20434),
            .in1(_gnd_net_),
            .in2(N__20274),
            .in3(N__20354),
            .lcout(),
            .ltout(\this_vga_signals.N_167_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_12_0_i_LC_18_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_12_0_i_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_12_0_i_LC_18_21_2 .LUT_INIT=16'b0100111100001111;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_12_0_i_LC_18_21_2  (
            .in0(N__20435),
            .in1(N__20271),
            .in2(N__20259),
            .in3(N__23763),
            .lcout(un1_M_this_state_q_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_6_LC_18_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_6_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_6_LC_18_21_3 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_6_LC_18_21_3  (
            .in0(N__35765),
            .in1(N__21168),
            .in2(N__25014),
            .in3(N__32393),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_13_LC_18_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_13_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_13_LC_18_21_4 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_13_LC_18_21_4  (
            .in0(N__31783),
            .in1(N__26357),
            .in2(N__32403),
            .in3(N__35763),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_5_LC_18_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_5_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_5_LC_18_21_5 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_5_LC_18_21_5  (
            .in0(N__35764),
            .in1(N__21427),
            .in2(N__25013),
            .in3(N__34684),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_0_LC_18_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_0_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_0_LC_18_21_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_0_LC_18_21_7  (
            .in0(N__26358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24332),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_5_LC_18_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_5_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_5_LC_18_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_5_LC_18_22_0  (
            .in0(_gnd_net_),
            .in1(N__21428),
            .in2(_gnd_net_),
            .in3(N__26356),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_5_LC_18_22_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_5_LC_18_22_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_5_LC_18_22_1.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_5_LC_18_22_1 (
            .in0(N__20256),
            .in1(N__27721),
            .in2(N__20250),
            .in3(N__21369),
            .lcout(M_this_sprites_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34527),
            .ce(),
            .sr(N__34017));
    defparam M_this_sprites_address_q_6_LC_18_22_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_6_LC_18_22_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_6_LC_18_22_4.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_sprites_address_q_6_LC_18_22_4 (
            .in0(N__27722),
            .in1(N__20247),
            .in2(N__20241),
            .in3(N__21135),
            .lcout(M_this_sprites_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34527),
            .ce(),
            .sr(N__34017));
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_7_LC_18_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_7_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_i_o3_0_7_LC_18_23_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_i_o3_0_7_LC_18_23_1  (
            .in0(N__20487),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21648),
            .lcout(),
            .ltout(this_vga_signals_M_this_state_q_ns_i_o3_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_18_23_2.C_ON=1'b0;
    defparam M_this_state_q_7_LC_18_23_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_18_23_2.LUT_INIT=16'b0000000011011100;
    LogicCell40 M_this_state_q_7_LC_18_23_2 (
            .in0(N__20608),
            .in1(N__23697),
            .in2(N__20556),
            .in3(N__35782),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34536),
            .ce(),
            .sr(N__34015));
    defparam \this_vga_signals.M_this_state_d_0_sqmuxa_i_LC_18_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d_0_sqmuxa_i_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d_0_sqmuxa_i_LC_18_23_4 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \this_vga_signals.M_this_state_d_0_sqmuxa_i_LC_18_23_4  (
            .in0(N__20429),
            .in1(N__20936),
            .in2(N__20895),
            .in3(N__20816),
            .lcout(N_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d_2_sqmuxa_0_LC_18_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d_2_sqmuxa_0_LC_18_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d_2_sqmuxa_0_LC_18_23_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.M_this_state_d_2_sqmuxa_0_LC_18_23_6  (
            .in0(N__32917),
            .in1(N__33671),
            .in2(N__33483),
            .in3(N__20551),
            .lcout(this_vga_signals_M_this_state_d_2_sqmuxa_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_6_LC_18_23_7.C_ON=1'b0;
    defparam M_this_state_q_6_LC_18_23_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_18_23_7.LUT_INIT=16'b1111111011111100;
    LogicCell40 M_this_state_q_6_LC_18_23_7 (
            .in0(N__20488),
            .in1(N__20459),
            .in2(N__23769),
            .in3(N__20523),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34536),
            .ce(),
            .sr(N__34015));
    defparam \this_vga_signals.un1_M_this_state_q_14_LC_18_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_14_LC_18_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_14_LC_18_24_0 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_14_LC_18_24_0  (
            .in0(N__20458),
            .in1(N__20436),
            .in2(N__27360),
            .in3(N__20358),
            .lcout(\this_vga_signals.un1_M_this_state_q_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_4_LC_18_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_4_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_4_LC_18_24_1 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_4_LC_18_24_1  (
            .in0(N__27445),
            .in1(N__35779),
            .in2(N__32594),
            .in3(N__25002),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_9_LC_18_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_9_LC_18_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_9_LC_18_24_3 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_9_LC_18_24_3  (
            .in0(N__22377),
            .in1(N__35780),
            .in2(N__33482),
            .in3(N__26375),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_LC_18_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_LC_18_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_LC_18_24_7 .LUT_INIT=16'b0000001100000111;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_LC_18_24_7  (
            .in0(N__23677),
            .in1(N__35778),
            .in2(N__23767),
            .in3(N__20343),
            .lcout(\this_vga_signals.M_this_sprites_ram_write_data_sn_N_4_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_19_15_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_19_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_19_15_4  (
            .in0(N__20313),
            .in1(N__20292),
            .in2(_gnd_net_),
            .in3(N__30459),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_11_LC_19_15_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_11_LC_19_15_7 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_11_LC_19_15_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \this_sprites_ram.mem_radreg_11_LC_19_15_7  (
            .in0(N__30081),
            .in1(N__30021),
            .in2(N__20760),
            .in3(N__30978),
            .lcout(\this_sprites_ram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34479),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_19_16_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_19_16_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_19_16_0 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_19_16_0  (
            .in0(N__21048),
            .in1(N__30372),
            .in2(N__24600),
            .in3(N__20673),
            .lcout(M_this_ppu_vram_data_3),
            .ltout(M_this_ppu_vram_data_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.vram_en_i_a2_0_LC_19_16_1 .C_ON=1'b0;
    defparam \this_ppu.vram_en_i_a2_0_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.vram_en_i_a2_0_LC_19_16_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.vram_en_i_a2_0_LC_19_16_1  (
            .in0(N__20708),
            .in1(N__21776),
            .in2(N__20697),
            .in3(N__20687),
            .lcout(\this_ppu.N_156 ),
            .ltout(\this_ppu.N_156_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI22N1G_5_LC_19_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI22N1G_5_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI22N1G_5_LC_19_16_2 .LUT_INIT=16'b1100111111001100;
    LogicCell40 \this_ppu.M_state_q_RNI22N1G_5_LC_19_16_2  (
            .in0(_gnd_net_),
            .in1(N__30006),
            .in2(N__20676),
            .in3(N__23504),
            .lcout(M_this_ppu_vram_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_6_LC_19_16_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_6_LC_19_16_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_6_LC_19_16_3 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \this_ppu.M_state_q_6_LC_19_16_3  (
            .in0(N__23505),
            .in1(N__23365),
            .in2(N__23784),
            .in3(N__22871),
            .lcout(\this_ppu.M_state_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34485),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_19_16_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_19_16_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_19_16_4 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_19_16_4  (
            .in0(N__24595),
            .in1(N__21093),
            .in2(N__29004),
            .in3(N__22995),
            .lcout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_19_17_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_19_17_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_19_17_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_19_17_0  (
            .in0(N__30424),
            .in1(N__20667),
            .in2(_gnd_net_),
            .in3(N__20649),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIRHU1G_1_LC_19_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIRHU1G_1_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIRHU1G_1_LC_19_17_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNIRHU1G_1_LC_19_17_3  (
            .in0(N__25517),
            .in1(N__25569),
            .in2(_gnd_net_),
            .in3(N__22605),
            .lcout(\this_ppu.un1_M_haddress_q_3_c2 ),
            .ltout(\this_ppu.un1_M_haddress_q_3_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI81A2G_4_LC_19_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI81A2G_4_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI81A2G_4_LC_19_17_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNI81A2G_4_LC_19_17_4  (
            .in0(N__25302),
            .in1(N__25382),
            .in2(N__20625),
            .in3(N__25464),
            .lcout(\this_ppu.un1_M_haddress_q_3_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_17_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_17_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_17_6  (
            .in0(N__30423),
            .in1(N__21126),
            .in2(_gnd_net_),
            .in3(N__21108),
            .lcout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_19_17_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_19_17_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_19_17_7  (
            .in0(N__21087),
            .in1(N__21066),
            .in2(_gnd_net_),
            .in3(N__30425),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_19_18_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_19_18_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_19_18_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_19_18_0  (
            .in0(_gnd_net_),
            .in1(N__21030),
            .in2(_gnd_net_),
            .in3(N__20943),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34501),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_19_18_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_19_18_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_19_18_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_19_18_3  (
            .in0(N__21029),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34501),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIGL6V4_0_LC_19_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIGL6V4_0_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIGL6V4_0_LC_19_18_4 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \this_ppu.M_state_q_RNIGL6V4_0_LC_19_18_4  (
            .in0(N__29474),
            .in1(N__29372),
            .in2(N__29435),
            .in3(N__34111),
            .lcout(\this_ppu.M_state_q_RNIGL6V4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_4_LC_19_20_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_4_LC_19_20_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_4_LC_19_20_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_4_LC_19_20_5 (
            .in0(N__32593),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34519),
            .ce(N__34163),
            .sr(N__34025));
    defparam \this_vga_signals.M_this_state_q_tr32_i_o3_LC_19_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_tr32_i_o3_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_tr32_i_o3_LC_19_21_1 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \this_vga_signals.M_this_state_q_tr32_i_o3_LC_19_21_1  (
            .in0(N__28133),
            .in1(N__20935),
            .in2(N__20894),
            .in3(N__20817),
            .lcout(N_156_0),
            .ltout(N_156_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_29_LC_19_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_29_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_29_LC_19_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_29_LC_19_21_2  (
            .in0(N__35435),
            .in1(N__34750),
            .in2(N__20775),
            .in3(N__34987),
            .lcout(N_35_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_RNO_1_LC_19_21_5.C_ON=1'b0;
    defparam M_this_substate_q_RNO_1_LC_19_21_5.SEQ_MODE=4'b0000;
    defparam M_this_substate_q_RNO_1_LC_19_21_5.LUT_INIT=16'b0100010000000000;
    LogicCell40 M_this_substate_q_RNO_1_LC_19_21_5 (
            .in0(N__21732),
            .in1(N__21689),
            .in2(_gnd_net_),
            .in3(N__21639),
            .lcout(M_this_substate_q_RNOZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI13IA1_1_1_LC_19_21_6.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI13IA1_1_1_LC_19_21_6.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI13IA1_1_1_LC_19_21_6.LUT_INIT=16'b1111111100000010;
    LogicCell40 M_this_oam_address_q_RNI13IA1_1_1_LC_19_21_6 (
            .in0(N__35080),
            .in1(N__34986),
            .in2(N__35467),
            .in3(N__34115),
            .lcout(N_1142_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNIQ61C7_0_LC_19_22_0.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNIQ61C7_0_LC_19_22_0.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNIQ61C7_0_LC_19_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNIQ61C7_0_LC_19_22_0 (
            .in0(_gnd_net_),
            .in1(N__24281),
            .in2(N__21606),
            .in3(N__21605),
            .lcout(M_this_sprites_address_q_RNIQ61C7Z0Z_0),
            .ltout(),
            .carryin(bfn_19_22_0_),
            .carryout(un1_M_this_sprites_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_19_22_1.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_19_22_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_19_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_19_22_1 (
            .in0(_gnd_net_),
            .in1(N__26097),
            .in2(_gnd_net_),
            .in3(N__21591),
            .lcout(un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_0),
            .carryout(un1_M_this_sprites_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_19_22_2.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_19_22_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_19_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_19_22_2 (
            .in0(_gnd_net_),
            .in1(N__22132),
            .in2(_gnd_net_),
            .in3(N__21588),
            .lcout(un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_1),
            .carryout(un1_M_this_sprites_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_19_22_3.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_19_22_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_19_22_3.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_19_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24038),
            .in3(N__21585),
            .lcout(un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_2),
            .carryout(un1_M_this_sprites_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_19_22_4.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_19_22_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_19_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_19_22_4 (
            .in0(_gnd_net_),
            .in1(N__27466),
            .in2(_gnd_net_),
            .in3(N__21582),
            .lcout(un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_3),
            .carryout(un1_M_this_sprites_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_19_22_5.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_19_22_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_19_22_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_19_22_5 (
            .in0(_gnd_net_),
            .in1(N__21401),
            .in2(_gnd_net_),
            .in3(N__21363),
            .lcout(un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_4),
            .carryout(un1_M_this_sprites_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_19_22_6.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_19_22_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_19_22_6.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_19_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21186),
            .in3(N__21129),
            .lcout(un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_5),
            .carryout(un1_M_this_sprites_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_19_22_7.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_19_22_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_19_22_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_19_22_7 (
            .in0(_gnd_net_),
            .in1(N__21860),
            .in2(_gnd_net_),
            .in3(N__21765),
            .lcout(un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_6),
            .carryout(un1_M_this_sprites_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_19_23_0.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_19_23_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_19_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_19_23_0 (
            .in0(_gnd_net_),
            .in1(N__26433),
            .in2(_gnd_net_),
            .in3(N__21762),
            .lcout(un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0),
            .ltout(),
            .carryin(bfn_19_23_0_),
            .carryout(un1_M_this_sprites_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_19_23_1.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_19_23_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_19_23_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_19_23_1 (
            .in0(_gnd_net_),
            .in1(N__22373),
            .in2(_gnd_net_),
            .in3(N__21759),
            .lcout(un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_8),
            .carryout(un1_M_this_sprites_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_19_23_2.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_19_23_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_19_23_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_19_23_2 (
            .in0(_gnd_net_),
            .in1(N__24688),
            .in2(_gnd_net_),
            .in3(N__21756),
            .lcout(un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_9),
            .carryout(un1_M_this_sprites_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_19_23_3.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_19_23_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_19_23_3.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_19_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31861),
            .in3(N__21753),
            .lcout(un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_10),
            .carryout(un1_M_this_sprites_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_19_23_4.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_19_23_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_19_23_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_19_23_4 (
            .in0(_gnd_net_),
            .in1(N__31940),
            .in2(_gnd_net_),
            .in3(N__21750),
            .lcout(un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_11),
            .carryout(un1_M_this_sprites_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_19_23_5.C_ON=1'b0;
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_19_23_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_19_23_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_19_23_5 (
            .in0(_gnd_net_),
            .in1(N__31724),
            .in2(_gnd_net_),
            .in3(N__21747),
            .lcout(un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_5_220_LC_19_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_5_220_LC_19_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_a3_5_220_LC_19_23_7 .LUT_INIT=16'b0000001100000111;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_a3_5_220_LC_19_23_7  (
            .in0(N__26735),
            .in1(N__28561),
            .in2(N__26666),
            .in3(N__28394),
            .lcout(M_this_state_d25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_9_LC_19_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_9_LC_19_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_9_LC_19_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_9_LC_19_24_0  (
            .in0(_gnd_net_),
            .in1(N__22418),
            .in2(_gnd_net_),
            .in3(N__25003),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_9_LC_19_24_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_9_LC_19_24_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_9_LC_19_24_1.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_sprites_address_q_9_LC_19_24_1 (
            .in0(N__27685),
            .in1(N__22587),
            .in2(N__22581),
            .in3(N__22578),
            .lcout(M_this_sprites_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34550),
            .ce(),
            .sr(N__34016));
    defparam \this_vga_signals.M_this_sprites_address_q_m_2_LC_19_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_2_LC_19_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_2_LC_19_24_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_2_LC_19_24_3  (
            .in0(_gnd_net_),
            .in1(N__22111),
            .in2(_gnd_net_),
            .in3(N__26376),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_2_LC_19_24_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_2_LC_19_24_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_2_LC_19_24_4.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_2_LC_19_24_4 (
            .in0(N__22314),
            .in1(N__27683),
            .in2(N__22305),
            .in3(N__22302),
            .lcout(M_this_sprites_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34550),
            .ce(),
            .sr(N__34016));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_3_LC_19_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_3_LC_19_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_3_LC_19_24_6 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_3_LC_19_24_6  (
            .in0(N__35851),
            .in1(N__24029),
            .in2(N__32832),
            .in3(N__25004),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_3_LC_19_24_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_3_LC_19_24_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_3_LC_19_24_7.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_sprites_address_q_3_LC_19_24_7 (
            .in0(N__27684),
            .in1(N__23940),
            .in2(N__22056),
            .in3(N__22053),
            .lcout(M_this_sprites_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34550),
            .ce(),
            .sr(N__34016));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_7_LC_19_25_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_7_LC_19_25_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_7_LC_19_25_3 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_7_LC_19_25_3  (
            .in0(N__35852),
            .in1(N__21839),
            .in2(N__33818),
            .in3(N__26374),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_7_LC_19_25_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_7_LC_19_25_4.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_7_LC_19_25_4.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_7_LC_19_25_4 (
            .in0(N__21798),
            .in1(N__27702),
            .in2(N__22044),
            .in3(N__22041),
            .lcout(M_this_sprites_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34558),
            .ce(),
            .sr(N__34013));
    defparam \this_vga_signals.M_this_sprites_address_q_m_7_LC_19_25_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_7_LC_19_25_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_7_LC_19_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_7_LC_19_25_5  (
            .in0(_gnd_net_),
            .in1(N__21838),
            .in2(_gnd_net_),
            .in3(N__25005),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_20_15_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_20_15_0 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_20_15_0  (
            .in0(N__23034),
            .in1(N__21792),
            .in2(N__24599),
            .in3(N__24546),
            .lcout(M_this_ppu_vram_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_20_15_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_20_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_wclke_3_LC_20_15_5  (
            .in0(N__31970),
            .in1(N__31863),
            .in2(N__31779),
            .in3(N__31649),
            .lcout(\this_sprites_ram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_20_15_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_20_15_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_20_15_7  (
            .in0(N__23061),
            .in1(N__23046),
            .in2(_gnd_net_),
            .in3(N__30460),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_20_16_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_20_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_20_16_1  (
            .in0(N__30464),
            .in1(N__23028),
            .in2(_gnd_net_),
            .in3(N__23013),
            .lcout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI42KTA_0_LC_20_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI42KTA_0_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI42KTA_0_LC_20_16_2 .LUT_INIT=16'b1111111100101010;
    LogicCell40 \this_ppu.M_state_q_RNI42KTA_0_LC_20_16_2  (
            .in0(N__28663),
            .in1(N__22988),
            .in2(N__22930),
            .in3(N__34112),
            .lcout(\this_ppu.M_state_q_RNI42KTAZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_1_LC_20_16_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_20_16_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.M_state_q_RNO_0_1_LC_20_16_5  (
            .in0(N__30019),
            .in1(N__23506),
            .in2(_gnd_net_),
            .in3(N__28664),
            .lcout(),
            .ltout(\this_ppu.N_150_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_1_LC_20_16_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_1_LC_20_16_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_1_LC_20_16_6 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \this_ppu.M_state_q_1_LC_20_16_6  (
            .in0(N__23507),
            .in1(N__23366),
            .in2(N__22875),
            .in3(N__22872),
            .lcout(\this_ppu.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34492),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI70261_2_LC_20_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI70261_2_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI70261_2_LC_20_17_0 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_ppu.M_haddress_q_RNI70261_2_LC_20_17_0  (
            .in0(N__29997),
            .in1(N__25098),
            .in2(N__30082),
            .in3(N__25462),
            .lcout(M_this_ppu_sprites_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_2_LC_20_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_2_LC_20_17_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_2_LC_20_17_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_haddress_q_2_LC_20_17_1  (
            .in0(N__22607),
            .in1(N__25468),
            .in2(N__25580),
            .in3(N__25520),
            .lcout(M_this_ppu_vram_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34502),
            .ce(),
            .sr(N__23130));
    defparam \this_ppu.M_haddress_q_1_LC_20_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_1_LC_20_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_1_LC_20_17_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_haddress_q_1_LC_20_17_2  (
            .in0(N__25519),
            .in1(N__25573),
            .in2(_gnd_net_),
            .in3(N__22606),
            .lcout(M_this_ppu_vram_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34502),
            .ce(),
            .sr(N__23130));
    defparam \this_ppu.M_haddress_q_0_LC_20_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_0_LC_20_17_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_0_LC_20_17_3 .LUT_INIT=16'b0101101001010110;
    LogicCell40 \this_ppu.M_haddress_q_0_LC_20_17_3  (
            .in0(N__25572),
            .in1(N__23508),
            .in2(N__30018),
            .in3(N__23370),
            .lcout(M_this_ppu_vram_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34502),
            .ce(),
            .sr(N__23130));
    defparam \this_ppu.M_haddress_q_RNI88B5_0_LC_20_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI88B5_0_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI88B5_0_LC_20_17_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \this_ppu.M_haddress_q_RNI88B5_0_LC_20_17_4  (
            .in0(N__28031),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25570),
            .lcout(),
            .ltout(\this_ppu.un2_hscroll_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIVK7O_0_LC_20_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIVK7O_0_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIVK7O_0_LC_20_17_5 .LUT_INIT=16'b1010101010001011;
    LogicCell40 \this_ppu.M_haddress_q_RNIVK7O_0_LC_20_17_5  (
            .in0(N__25571),
            .in1(N__30055),
            .in2(N__23349),
            .in3(N__29998),
            .lcout(M_this_ppu_sprites_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_3_LC_20_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_3_LC_20_17_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_3_LC_20_17_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_haddress_q_3_LC_20_17_6  (
            .in0(N__25383),
            .in1(N__25463),
            .in2(_gnd_net_),
            .in3(N__23138),
            .lcout(M_this_ppu_map_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34502),
            .ce(),
            .sr(N__23130));
    defparam \this_ppu.M_haddress_q_4_LC_20_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_4_LC_20_17_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_4_LC_20_17_7 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_haddress_q_4_LC_20_17_7  (
            .in0(N__23139),
            .in1(N__25384),
            .in2(N__25312),
            .in3(N__25469),
            .lcout(M_this_ppu_map_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34502),
            .ce(),
            .sr(N__23130));
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_20_18_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_20_18_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_wclke_3_LC_20_18_0  (
            .in0(N__31969),
            .in1(N__31862),
            .in2(N__31790),
            .in3(N__31645),
            .lcout(\this_sprites_ram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_4_LC_20_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_4_LC_20_18_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_idx_q_4_LC_20_18_2 .LUT_INIT=16'b0110000010100000;
    LogicCell40 \this_ppu.M_oam_idx_q_4_LC_20_18_2  (
            .in0(N__23393),
            .in1(N__23820),
            .in2(N__23910),
            .in3(N__23478),
            .lcout(\this_ppu.M_oam_idx_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34510),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_2_LC_20_18_3 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_2_LC_20_18_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_idx_q_2_LC_20_18_3 .LUT_INIT=16'b0010100010100000;
    LogicCell40 \this_ppu.M_oam_idx_q_2_LC_20_18_3  (
            .in0(N__23906),
            .in1(N__23864),
            .in2(N__23456),
            .in3(N__23886),
            .lcout(M_this_ppu_oam_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34510),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_1_LC_20_18_4.C_ON=1'b0;
    defparam M_this_oam_address_q_1_LC_20_18_4.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_1_LC_20_18_4.LUT_INIT=16'b0010100010100000;
    LogicCell40 M_this_oam_address_q_1_LC_20_18_4 (
            .in0(N__30682),
            .in1(N__35189),
            .in2(N__35418),
            .in3(N__34982),
            .lcout(M_this_oam_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34510),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI01PG1_1_LC_20_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI01PG1_1_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI01PG1_1_LC_20_18_5 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \this_ppu.M_state_q_RNI01PG1_1_LC_20_18_5  (
            .in0(N__25910),
            .in1(N__25856),
            .in2(_gnd_net_),
            .in3(N__34108),
            .lcout(\this_ppu.N_1046_0 ),
            .ltout(\this_ppu.N_1046_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_3_LC_20_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_3_LC_20_18_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_idx_q_3_LC_20_18_6 .LUT_INIT=16'b0011000011000000;
    LogicCell40 \this_ppu.M_oam_idx_q_3_LC_20_18_6  (
            .in0(_gnd_net_),
            .in1(N__23819),
            .in2(N__23511),
            .in3(N__23477),
            .lcout(M_this_ppu_oam_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34510),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_0_LC_20_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_0_LC_20_19_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_idx_q_0_LC_20_19_0 .LUT_INIT=16'b1011010000000000;
    LogicCell40 \this_ppu.M_oam_idx_q_0_LC_20_19_0  (
            .in0(N__26012),
            .in1(N__25951),
            .in2(N__23420),
            .in3(N__23905),
            .lcout(M_this_ppu_oam_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34520),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_5_LC_20_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_5_LC_20_19_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_5_LC_20_19_1 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \this_ppu.M_state_q_5_LC_20_19_1  (
            .in0(N__34120),
            .in1(_gnd_net_),
            .in2(N__25953),
            .in3(N__26011),
            .lcout(\this_ppu.M_state_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34520),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_3_LC_20_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_3_LC_20_19_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_3_LC_20_19_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_state_q_3_LC_20_19_2  (
            .in0(_gnd_net_),
            .in1(N__23376),
            .in2(_gnd_net_),
            .in3(N__34119),
            .lcout(\this_ppu.M_state_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34520),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIGJUB2_3_LC_20_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIGJUB2_3_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIGJUB2_3_LC_20_19_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.M_state_q_RNIGJUB2_3_LC_20_19_3  (
            .in0(N__25947),
            .in1(N__23413),
            .in2(_gnd_net_),
            .in3(N__26010),
            .lcout(\this_ppu.un1_M_oam_idx_q_1_c1 ),
            .ltout(\this_ppu.un1_M_oam_idx_q_1_c1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_RNIHI6C2_2_LC_20_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_RNIHI6C2_2_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_idx_q_RNIHI6C2_2_LC_20_19_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \this_ppu.M_oam_idx_q_RNIHI6C2_2_LC_20_19_4  (
            .in0(N__23862),
            .in1(_gnd_net_),
            .in2(N__23481),
            .in3(N__23449),
            .lcout(\this_ppu.un1_M_oam_idx_q_1_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_RNI3VF_4_LC_20_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_RNI3VF_4_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_idx_q_RNI3VF_4_LC_20_19_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_ppu.M_oam_idx_q_RNI3VF_4_LC_20_19_5  (
            .in0(N__23448),
            .in1(N__23412),
            .in2(N__23394),
            .in3(N__23861),
            .lcout(\this_ppu.N_144_4 ),
            .ltout(\this_ppu.N_144_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_4_LC_20_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_4_LC_20_19_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_4_LC_20_19_6 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \this_ppu.M_state_q_4_LC_20_19_6  (
            .in0(N__25994),
            .in1(N__23821),
            .in2(N__23379),
            .in3(N__34121),
            .lcout(\this_ppu.M_state_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34520),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_idx_q_1_LC_20_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_oam_idx_q_1_LC_20_19_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_idx_q_1_LC_20_19_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_ppu.M_oam_idx_q_1_LC_20_19_7  (
            .in0(N__23904),
            .in1(N__23863),
            .in2(_gnd_net_),
            .in3(N__23885),
            .lcout(M_this_ppu_oam_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34520),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_6_LC_20_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_6_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_6_LC_20_20_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_ppu.M_state_q_RNO_0_6_LC_20_20_3  (
            .in0(N__23825),
            .in1(N__23790),
            .in2(N__25995),
            .in3(N__34110),
            .lcout(\this_ppu.N_144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_en_iv_0_LC_20_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_en_iv_0_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_en_iv_0_LC_20_21_1 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_en_iv_0_LC_20_21_1  (
            .in0(N__23768),
            .in1(N__23701),
            .in2(_gnd_net_),
            .in3(N__35783),
            .lcout(M_this_sprites_ram_write_en_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_12_LC_20_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_12_LC_20_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_12_LC_20_21_2 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_12_LC_20_21_2  (
            .in0(N__35784),
            .in1(N__31967),
            .in2(N__34761),
            .in3(N__26379),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_2_LC_20_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_2_LC_20_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_2_LC_20_21_3 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_2_LC_20_21_3  (
            .in0(N__33454),
            .in1(N__27400),
            .in2(N__32389),
            .in3(N__27369),
            .lcout(M_this_sprites_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_0_LC_20_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_0_LC_20_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_8_m_0_LC_20_21_7 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_8_m_0_LC_20_21_7  (
            .in0(N__24282),
            .in1(N__25012),
            .in2(N__33833),
            .in3(N__35785),
            .lcout(\this_vga_signals.M_this_sprites_address_d_8_mZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_20_22_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_20_22_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_20_22_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_sprites_ram.mem_mem_4_0_wclke_3_LC_20_22_0  (
            .in0(N__31947),
            .in1(N__31626),
            .in2(N__31753),
            .in3(N__31845),
            .lcout(\this_sprites_ram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_11_LC_20_22_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_11_LC_20_22_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_11_LC_20_22_1.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_11_LC_20_22_1 (
            .in0(N__26748),
            .in1(N__27725),
            .in2(N__24249),
            .in3(N__23535),
            .lcout(M_this_sprites_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34544),
            .ce(),
            .sr(N__34022));
    defparam M_this_sprites_address_q_13_LC_20_22_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_13_LC_20_22_2.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_13_LC_20_22_2.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_sprites_address_q_13_LC_20_22_2 (
            .in0(N__27727),
            .in1(N__23529),
            .in2(N__23922),
            .in3(N__23517),
            .lcout(M_this_sprites_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34544),
            .ce(),
            .sr(N__34022));
    defparam M_this_sprites_address_q_12_LC_20_22_3.C_ON=1'b0;
    defparam M_this_sprites_address_q_12_LC_20_22_3.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_12_LC_20_22_3.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_12_LC_20_22_3 (
            .in0(N__24507),
            .in1(N__27726),
            .in2(N__23934),
            .in3(N__24501),
            .lcout(M_this_sprites_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34544),
            .ce(),
            .sr(N__34022));
    defparam M_this_sprites_address_q_0_LC_20_22_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_0_LC_20_22_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_0_LC_20_22_5.LUT_INIT=16'b1111101011111110;
    LogicCell40 M_this_sprites_address_q_0_LC_20_22_5 (
            .in0(N__24495),
            .in1(N__24489),
            .in2(N__24483),
            .in3(N__27724),
            .lcout(M_this_sprites_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34544),
            .ce(),
            .sr(N__34022));
    defparam \this_vga_signals.M_this_sprites_address_q_m_11_LC_20_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_11_LC_20_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_11_LC_20_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_11_LC_20_23_1  (
            .in0(_gnd_net_),
            .in1(N__24985),
            .in2(_gnd_net_),
            .in3(N__31844),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_RNO_0_LC_20_23_3.C_ON=1'b0;
    defparam M_this_substate_q_RNO_0_LC_20_23_3.SEQ_MODE=4'b0000;
    defparam M_this_substate_q_RNO_0_LC_20_23_3.LUT_INIT=16'b1100101000000000;
    LogicCell40 M_this_substate_q_RNO_0_LC_20_23_3 (
            .in0(N__28557),
            .in1(N__28464),
            .in2(N__24648),
            .in3(N__24237),
            .lcout(M_this_substate_q_s_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_8_LC_20_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_8_LC_20_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_8_LC_20_23_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_8_LC_20_23_5  (
            .in0(_gnd_net_),
            .in1(N__24986),
            .in2(_gnd_net_),
            .in3(N__26419),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_data_ibuf_RNIC68K4_5_LC_20_23_6.C_ON=1'b0;
    defparam port_data_ibuf_RNIC68K4_5_LC_20_23_6.SEQ_MODE=4'b0000;
    defparam port_data_ibuf_RNIC68K4_5_LC_20_23_6.LUT_INIT=16'b0000000001111111;
    LogicCell40 port_data_ibuf_RNIC68K4_5_LC_20_23_6 (
            .in0(N__24219),
            .in1(N__24204),
            .in2(N__34762),
            .in3(N__34107),
            .lcout(N_1152_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_3_LC_20_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_3_LC_20_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_3_LC_20_23_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_3_LC_20_23_7  (
            .in0(_gnd_net_),
            .in1(N__23999),
            .in2(_gnd_net_),
            .in3(N__26384),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_12_LC_20_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_12_LC_20_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_12_LC_20_24_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_12_LC_20_24_4  (
            .in0(N__24997),
            .in1(N__31968),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_13_LC_20_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_13_LC_20_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_13_LC_20_24_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_13_LC_20_24_5  (
            .in0(_gnd_net_),
            .in1(N__24996),
            .in2(_gnd_net_),
            .in3(N__31749),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_10_LC_20_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_10_LC_20_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_10_LC_20_24_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_10_LC_20_24_6  (
            .in0(N__24998),
            .in1(N__24690),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_10_LC_20_24_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_10_LC_20_24_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_10_LC_20_24_7.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_10_LC_20_24_7 (
            .in0(N__24654),
            .in1(N__27703),
            .in2(N__24888),
            .in3(N__24885),
            .lcout(M_this_sprites_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34559),
            .ce(),
            .sr(N__34018));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_10_LC_20_25_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_10_LC_20_25_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_10_LC_20_25_0 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_10_LC_20_25_0  (
            .in0(N__24689),
            .in1(N__32823),
            .in2(N__26385),
            .in3(N__35850),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_RNO_3_LC_20_25_1.C_ON=1'b0;
    defparam M_this_substate_q_RNO_3_LC_20_25_1.SEQ_MODE=4'b0000;
    defparam M_this_substate_q_RNO_3_LC_20_25_1.LUT_INIT=16'b0000000001010101;
    LogicCell40 M_this_substate_q_RNO_3_LC_20_25_1 (
            .in0(N__26731),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28364),
            .lcout(M_this_substate_q_RNOZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_m_4_LC_20_25_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_4_LC_20_25_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_4_LC_20_25_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_4_LC_20_25_3  (
            .in0(_gnd_net_),
            .in1(N__27441),
            .in2(_gnd_net_),
            .in3(N__26383),
            .lcout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_21_15_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_21_15_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_21_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_21_15_1  (
            .in0(N__30453),
            .in1(N__24636),
            .in2(_gnd_net_),
            .in3(N__24621),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_21_15_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_21_15_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_21_15_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_21_15_2  (
            .in0(N__28989),
            .in1(N__24587),
            .in2(N__24549),
            .in3(N__24513),
            .lcout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_15_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_15_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_15_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_15_5  (
            .in0(N__30454),
            .in1(N__24540),
            .in2(_gnd_net_),
            .in3(N__24525),
            .lcout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_hscroll_cry_0_c_inv_LC_21_16_0 .C_ON=1'b1;
    defparam \this_ppu.un2_hscroll_cry_0_c_inv_LC_21_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_hscroll_cry_0_c_inv_LC_21_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un2_hscroll_cry_0_c_inv_LC_21_16_0  (
            .in0(_gnd_net_),
            .in1(N__25568),
            .in2(N__25113),
            .in3(N__28030),
            .lcout(\this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ),
            .ltout(),
            .carryin(bfn_21_16_0_),
            .carryout(\this_ppu.un2_hscroll_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_21_16_1 .C_ON=1'b1;
    defparam \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_21_16_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_21_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_21_16_1  (
            .in0(_gnd_net_),
            .in1(N__25502),
            .in2(N__25029),
            .in3(N__25104),
            .lcout(\this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0 ),
            .ltout(),
            .carryin(\this_ppu.un2_hscroll_cry_0 ),
            .carryout(\this_ppu.un2_hscroll_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_21_16_2 .C_ON=1'b0;
    defparam \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_21_16_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_21_16_2  (
            .in0(N__27931),
            .in1(N__25461),
            .in2(_gnd_net_),
            .in3(N__25101),
            .lcout(\this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_21_16_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_21_16_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_wclke_3_LC_21_16_3  (
            .in0(N__31988),
            .in1(N__31886),
            .in2(N__31799),
            .in3(N__31660),
            .lcout(\this_sprites_ram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIPG425_1_LC_21_16_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIPG425_1_LC_21_16_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIPG425_1_LC_21_16_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIPG425_1_LC_21_16_7  (
            .in0(N__28672),
            .in1(N__28715),
            .in2(_gnd_net_),
            .in3(N__29327),
            .lcout(\this_ppu.un1_M_vaddress_q_2_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_21_17_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_21_17_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_21_17_0  (
            .in0(N__30449),
            .in1(N__25068),
            .in2(_gnd_net_),
            .in3(N__25050),
            .lcout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_21_17_1 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_21_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_21_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30927),
            .lcout(M_this_oam_ram_read_data_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_21_17_2 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_21_17_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_oam_ram.mem_mem_0_0_RNISG75_LC_21_17_2  (
            .in0(N__27980),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_oam_ram_read_data_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc1_LC_21_17_5 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc1_LC_21_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc1_LC_21_17_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc1_LC_21_17_5  (
            .in0(_gnd_net_),
            .in1(N__30871),
            .in2(_gnd_net_),
            .in3(N__30928),
            .lcout(\this_ppu.un1_M_haddress_q_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI4S061_1_LC_21_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI4S061_1_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI4S061_1_LC_21_17_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_ppu.M_haddress_q_RNI4S061_1_LC_21_17_6  (
            .in0(N__29991),
            .in1(N__25020),
            .in2(N__30153),
            .in3(N__25518),
            .lcout(M_this_ppu_sprites_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_21_18_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_21_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_21_18_0  (
            .in0(_gnd_net_),
            .in1(N__28044),
            .in2(N__28032),
            .in3(N__25567),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_0 ),
            .ltout(),
            .carryin(bfn_21_18_0_),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_21_18_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_21_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_21_18_1  (
            .in0(_gnd_net_),
            .in1(N__27993),
            .in2(N__27981),
            .in3(N__25501),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_0 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_21_18_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_21_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_21_18_2  (
            .in0(_gnd_net_),
            .in1(N__27948),
            .in2(N__27936),
            .in3(N__25460),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_1 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_21_18_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_21_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_21_18_3  (
            .in0(_gnd_net_),
            .in1(N__27896),
            .in2(N__25425),
            .in3(N__25381),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_0 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_2 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_21_18_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_21_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_21_18_4  (
            .in0(_gnd_net_),
            .in1(N__28283),
            .in2(N__25347),
            .in3(N__25301),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_3 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_21_18_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_21_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_21_18_5  (
            .in0(_gnd_net_),
            .in1(N__28269),
            .in2(N__28083),
            .in3(N__25256),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_4 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_21_18_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_21_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_21_18_6  (
            .in0(_gnd_net_),
            .in1(N__28257),
            .in2(N__31056),
            .in3(N__25192),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_3 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_5 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_21_18_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_21_18_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_21_18_7  (
            .in0(N__25139),
            .in1(N__30747),
            .in2(N__28245),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_4 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_6 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIFEE22_LC_21_19_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIFEE22_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIFEE22_LC_21_19_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIFEE22_LC_21_19_0  (
            .in0(N__28227),
            .in1(N__28089),
            .in2(_gnd_net_),
            .in3(N__26016),
            .lcout(\this_ppu.vscroll8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_2_LC_21_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_2_LC_21_19_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_2_LC_21_19_2 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \this_ppu.M_state_q_2_LC_21_19_2  (
            .in0(N__25830),
            .in1(N__34122),
            .in2(N__25926),
            .in3(N__26013),
            .lcout(\this_ppu.M_state_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34528),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_20_LC_21_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_20_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_20_LC_21_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_20_LC_21_19_4  (
            .in0(N__35340),
            .in1(N__35165),
            .in2(N__25824),
            .in3(N__34994),
            .lcout(N_48_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_28_LC_21_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_28_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_28_LC_21_19_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_28_LC_21_19_6  (
            .in0(N__35341),
            .in1(N__35164),
            .in2(N__32592),
            .in3(N__34995),
            .lcout(M_this_oam_ram_write_data_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_2_LC_21_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_2_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_2_LC_21_19_7 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \this_ppu.M_state_q_RNO_0_2_LC_21_19_7  (
            .in0(N__25952),
            .in1(N__25911),
            .in2(_gnd_net_),
            .in3(N__25857),
            .lcout(\this_ppu.N_148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_20_LC_21_20_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_20_LC_21_20_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_20_LC_21_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_20_LC_21_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32578),
            .lcout(M_this_data_tmp_qZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34537),
            .ce(N__31449),
            .sr(N__34027));
    defparam M_this_oam_address_q_RNI13IA1_0_1_LC_21_21_0.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI13IA1_0_1_LC_21_21_0.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI13IA1_0_1_LC_21_21_0.LUT_INIT=16'b1111111100100000;
    LogicCell40 M_this_oam_address_q_RNI13IA1_0_1_LC_21_21_0 (
            .in0(N__35119),
            .in1(N__35400),
            .in2(N__35003),
            .in3(N__34116),
            .lcout(N_1134_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_8_LC_21_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_8_LC_21_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_8_LC_21_21_1 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_8_LC_21_21_1  (
            .in0(N__26434),
            .in1(N__26378),
            .in2(N__32985),
            .in3(N__35787),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d21_6_LC_21_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d21_6_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d21_6_LC_21_21_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_d21_6_LC_21_21_3  (
            .in0(N__28527),
            .in1(N__28214),
            .in2(N__28167),
            .in3(N__28191),
            .lcout(\this_vga_signals.M_this_state_d21Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_21_21_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_21_21_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_21_21_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_5_0_wclke_3_LC_21_21_5  (
            .in0(N__31627),
            .in1(N__31948),
            .in2(N__31754),
            .in3(N__31846),
            .lcout(\this_sprites_ram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d22_LC_21_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d22_LC_21_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d22_LC_21_22_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vga_signals.M_this_state_d22_LC_21_22_0  (
            .in0(N__28502),
            .in1(N__28395),
            .in2(N__26682),
            .in3(N__28454),
            .lcout(M_this_state_d22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_11_LC_21_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_11_LC_21_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_d_5_m_11_LC_21_22_5 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_d_5_m_11_LC_21_22_5  (
            .in0(N__31843),
            .in1(N__26377),
            .in2(N__32568),
            .in3(N__35846),
            .lcout(\this_vga_signals.M_this_sprites_address_d_5_mZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d24_LC_21_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d24_LC_21_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d24_LC_21_22_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.M_this_state_d24_LC_21_22_7  (
            .in0(N__26739),
            .in1(N__26681),
            .in2(N__28329),
            .in3(N__28503),
            .lcout(\this_vga_signals.M_this_state_dZ0Z24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_9_LC_21_23_0.C_ON=1'b0;
    defparam M_this_external_address_q_9_LC_21_23_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_9_LC_21_23_0.LUT_INIT=16'b1110110001001100;
    LogicCell40 M_this_external_address_q_9_LC_21_23_0 (
            .in0(N__35610),
            .in1(N__32019),
            .in2(N__35871),
            .in3(N__32926),
            .lcout(M_this_external_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34560),
            .ce(),
            .sr(N__34023));
    defparam M_this_sprites_address_q_8_LC_21_23_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_8_LC_21_23_2.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_8_LC_21_23_2.LUT_INIT=16'b1111110111111100;
    LogicCell40 M_this_sprites_address_q_8_LC_21_23_2 (
            .in0(N__27729),
            .in1(N__26640),
            .in2(N__26631),
            .in3(N__26622),
            .lcout(M_this_sprites_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34560),
            .ce(),
            .sr(N__34023));
    defparam \this_vga_signals.M_this_sprites_address_q_m_1_LC_21_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_m_1_LC_21_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_m_1_LC_21_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_m_1_LC_21_23_4  (
            .in0(_gnd_net_),
            .in1(N__26044),
            .in2(_gnd_net_),
            .in3(N__26352),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_q_mZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_1_LC_21_23_5.C_ON=1'b0;
    defparam M_this_sprites_address_q_1_LC_21_23_5.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_1_LC_21_23_5.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_1_LC_21_23_5 (
            .in0(N__26250),
            .in1(N__27728),
            .in2(N__26238),
            .in3(N__26235),
            .lcout(M_this_sprites_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34560),
            .ce(),
            .sr(N__34023));
    defparam M_this_sprites_address_q_4_LC_21_24_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_4_LC_21_24_0.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_4_LC_21_24_0.LUT_INIT=16'b1111101111111010;
    LogicCell40 M_this_sprites_address_q_4_LC_21_24_0 (
            .in0(N__27738),
            .in1(N__27723),
            .in2(N__27654),
            .in3(N__27645),
            .lcout(M_this_sprites_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34568),
            .ce(),
            .sr(N__34020));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_LC_21_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_LC_21_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_LC_21_24_5 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_1_LC_21_24_5  (
            .in0(N__32955),
            .in1(N__27405),
            .in2(N__34739),
            .in3(N__27361),
            .lcout(M_this_sprites_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_7_LC_22_14_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_7_LC_22_14_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_7_LC_22_14_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_7_LC_22_14_1 (
            .in0(N__33630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34493),
            .ce(N__34198),
            .sr(N__34036));
    defparam \this_ppu.M_state_q_RNI53UU_6_LC_22_15_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI53UU_6_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI53UU_6_LC_22_15_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \this_ppu.M_state_q_RNI53UU_6_LC_22_15_0  (
            .in0(N__27222),
            .in1(N__30017),
            .in2(N__31041),
            .in3(N__30112),
            .lcout(M_this_ppu_sprites_addr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIFH3G1_1_LC_22_15_1 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIFH3G1_1_LC_22_15_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIFH3G1_1_LC_22_15_1 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_ppu.M_vaddress_q_RNIFH3G1_1_LC_22_15_1  (
            .in0(N__30016),
            .in1(N__29040),
            .in2(N__30136),
            .in3(N__28711),
            .lcout(M_this_ppu_sprites_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_1_LC_22_15_2 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_1_LC_22_15_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_1_LC_22_15_2 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \this_ppu.M_vaddress_q_1_LC_22_15_2  (
            .in0(N__29326),
            .in1(_gnd_net_),
            .in2(N__28721),
            .in3(N__28676),
            .lcout(\this_ppu.M_vaddress_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34503),
            .ce(),
            .sr(N__29264));
    defparam \this_ppu.M_vaddress_q_5_LC_22_15_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_5_LC_22_15_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_5_LC_22_15_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_ppu.M_vaddress_q_5_LC_22_15_4  (
            .in0(N__27881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27851),
            .lcout(M_this_ppu_map_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34503),
            .ce(),
            .sr(N__29264));
    defparam \this_ppu.M_vaddress_q_6_LC_22_15_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_6_LC_22_15_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_6_LC_22_15_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_vaddress_q_6_LC_22_15_6  (
            .in0(N__27882),
            .in1(N__27801),
            .in2(_gnd_net_),
            .in3(N__27852),
            .lcout(M_this_ppu_map_addr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34503),
            .ce(),
            .sr(N__29264));
    defparam \this_ppu.M_vaddress_q_7_LC_22_15_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_7_LC_22_15_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_7_LC_22_15_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \this_ppu.M_vaddress_q_7_LC_22_15_7  (
            .in0(N__27853),
            .in1(N__27880),
            .in2(N__27809),
            .in3(N__27760),
            .lcout(M_this_ppu_map_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34503),
            .ce(),
            .sr(N__29264));
    defparam \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_22_16_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_22_16_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_22_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_22_16_7  (
            .in0(N__29506),
            .in1(N__29556),
            .in2(N__29594),
            .in3(N__29630),
            .lcout(\this_ppu.un1_M_vaddress_q_2_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_22_17_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_22_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_22_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_22_17_0  (
            .in0(_gnd_net_),
            .in1(N__29213),
            .in2(N__29198),
            .in3(N__29302),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_7 ),
            .ltout(),
            .carryin(bfn_22_17_0_),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_22_17_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_22_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_22_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_22_17_1  (
            .in0(_gnd_net_),
            .in1(N__29147),
            .in2(N__31206),
            .in3(N__28716),
            .lcout(\this_ppu.M_vaddress_q_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_0 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_22_17_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_22_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_22_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_22_17_2  (
            .in0(_gnd_net_),
            .in1(N__29132),
            .in2(N__29118),
            .in3(N__29628),
            .lcout(\this_ppu.M_vaddress_q_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_1 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_22_17_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_22_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_22_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_22_17_3  (
            .in0(_gnd_net_),
            .in1(N__30332),
            .in2(N__31509),
            .in3(N__29555),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_5 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_2 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_22_17_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_22_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_22_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_22_17_4  (
            .in0(_gnd_net_),
            .in1(N__30314),
            .in2(N__30945),
            .in3(N__29505),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_6 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_3 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_22_17_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_22_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_22_17_5  (
            .in0(_gnd_net_),
            .in1(N__30296),
            .in2(N__31221),
            .in3(N__27857),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_7 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_4 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_22_17_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_22_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_22_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_22_17_6  (
            .in0(_gnd_net_),
            .in1(N__30278),
            .in2(N__31347),
            .in3(N__27808),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_8 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_5 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_22_17_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_22_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_22_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_22_17_7  (
            .in0(_gnd_net_),
            .in1(N__31392),
            .in2(N__30264),
            .in3(N__27764),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_9 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_6 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_22_18_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_22_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_22_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28092),
            .lcout(\this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc2_LC_22_18_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc2_LC_22_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc2_LC_22_18_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc2_LC_22_18_1  (
            .in0(N__30782),
            .in1(N__30879),
            .in2(_gnd_net_),
            .in3(N__30930),
            .lcout(\this_ppu.un1_M_haddress_q_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNO_0_4_LC_22_18_4.C_ON=1'b0;
    defparam M_this_oam_address_q_RNO_0_4_LC_22_18_4.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNO_0_4_LC_22_18_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_oam_address_q_RNO_0_4_LC_22_18_4 (
            .in0(N__35398),
            .in1(N__35175),
            .in2(N__34996),
            .in3(N__30590),
            .lcout(),
            .ltout(un1_M_this_oam_address_q_c3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_4_LC_22_18_5.C_ON=1'b0;
    defparam M_this_oam_address_q_4_LC_22_18_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_4_LC_22_18_5.LUT_INIT=16'b0010100010001000;
    LogicCell40 M_this_oam_address_q_4_LC_22_18_5 (
            .in0(N__30689),
            .in1(N__30181),
            .in2(N__28071),
            .in3(N__30634),
            .lcout(M_this_oam_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34529),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_7_LC_22_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_7_LC_22_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_7_LC_22_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_7_LC_22_18_6  (
            .in0(N__35397),
            .in1(N__35174),
            .in2(N__28068),
            .in3(N__34922),
            .lcout(N_65_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_0_c_LC_22_19_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_0_c_LC_22_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_0_c_LC_22_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_0_c_LC_22_19_0  (
            .in0(_gnd_net_),
            .in1(N__28043),
            .in2(N__28026),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_22_19_0_),
            .carryout(\this_ppu.un1_M_haddress_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_1_c_LC_22_19_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_1_c_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_1_c_LC_22_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_1_c_LC_22_19_1  (
            .in0(_gnd_net_),
            .in1(N__27992),
            .in2(N__27976),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_0 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_2_c_LC_22_19_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_2_c_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_2_c_LC_22_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_2_c_LC_22_19_2  (
            .in0(_gnd_net_),
            .in1(N__27947),
            .in2(N__27932),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_1 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_3_c_LC_22_19_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_3_c_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_3_c_LC_22_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_3_c_LC_22_19_3  (
            .in0(_gnd_net_),
            .in1(N__30929),
            .in2(N__27897),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_2 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_4_c_LC_22_19_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_4_c_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_4_c_LC_22_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_4_c_LC_22_19_4  (
            .in0(_gnd_net_),
            .in1(N__30878),
            .in2(N__28284),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_3 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_5_c_LC_22_19_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_5_c_LC_22_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_5_c_LC_22_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_5_c_LC_22_19_5  (
            .in0(_gnd_net_),
            .in1(N__28268),
            .in2(N__30786),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_4 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_6_c_LC_22_19_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_6_c_LC_22_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_6_c_LC_22_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_6_c_LC_22_19_6  (
            .in0(_gnd_net_),
            .in1(N__28256),
            .in2(N__30819),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_5 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_7_c_LC_22_19_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_7_c_LC_22_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_7_c_LC_22_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_7_c_LC_22_19_7  (
            .in0(_gnd_net_),
            .in1(N__28241),
            .in2(N__30840),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_6 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_RNI6VRP1_LC_22_20_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_RNI6VRP1_LC_22_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_RNI6VRP1_LC_22_20_0 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_7_c_RNI6VRP1_LC_22_20_0  (
            .in0(N__30957),
            .in1(N__31068),
            .in2(N__30243),
            .in3(N__28230),
            .lcout(\this_ppu.vscroll8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_2_LC_22_20_6.C_ON=1'b0;
    defparam M_this_oam_address_q_2_LC_22_20_6.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_2_LC_22_20_6.LUT_INIT=16'b0100010010001000;
    LogicCell40 M_this_oam_address_q_2_LC_22_20_6 (
            .in0(N__30585),
            .in1(N__30683),
            .in2(_gnd_net_),
            .in3(N__30552),
            .lcout(M_this_oam_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34545),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d21_6_x_LC_22_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d21_6_x_LC_22_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d21_6_x_LC_22_20_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_this_state_d21_6_x_LC_22_20_7  (
            .in0(N__28221),
            .in1(N__28187),
            .in2(_gnd_net_),
            .in3(N__28160),
            .lcout(M_this_state_d21_6_x),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNILT531_12_LC_22_21_4.C_ON=1'b0;
    defparam M_this_state_q_RNILT531_12_LC_22_21_4.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNILT531_12_LC_22_21_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_state_q_RNILT531_12_LC_22_21_4 (
            .in0(N__34935),
            .in1(N__28137),
            .in2(N__35469),
            .in3(N__35786),
            .lcout(un1_M_this_oam_address_q_c2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_13_LC_22_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_13_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_13_LC_22_21_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_13_LC_22_21_5  (
            .in0(N__35452),
            .in1(N__35098),
            .in2(N__28593),
            .in3(N__34936),
            .lcout(N_56_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_13_LC_22_22_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_13_LC_22_22_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_13_LC_22_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_13_LC_22_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34695),
            .lcout(M_this_data_tmp_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34561),
            .ce(N__32188),
            .sr(N__34026));
    defparam \this_vga_signals.M_this_state_d21_1_LC_22_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d21_1_LC_22_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d21_1_LC_22_23_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.M_this_state_d21_1_LC_22_23_0  (
            .in0(N__28501),
            .in1(N__28478),
            .in2(N__28455),
            .in3(N__28520),
            .lcout(M_this_state_d21_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_RNO_2_LC_22_23_3.C_ON=1'b0;
    defparam M_this_substate_q_RNO_2_LC_22_23_3.SEQ_MODE=4'b0000;
    defparam M_this_substate_q_RNO_2_LC_22_23_3.LUT_INIT=16'b0000000001000000;
    LogicCell40 M_this_substate_q_RNO_2_LC_22_23_3 (
            .in0(N__28519),
            .in1(N__28500),
            .in2(N__28479),
            .in3(N__28450),
            .lcout(M_this_substate_q_RNOZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d24_1_LC_22_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d24_1_LC_22_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d24_1_LC_22_24_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_this_state_d24_1_LC_22_24_5  (
            .in0(N__28441),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28382),
            .lcout(\this_vga_signals.M_this_state_d24Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_22_24_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_22_24_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_22_24_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_sprites_ram.mem_mem_7_0_wclke_3_LC_22_24_6  (
            .in0(N__31983),
            .in1(N__31875),
            .in2(N__31791),
            .in3(N__31659),
            .lcout(\this_sprites_ram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_3_LC_22_26_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_3_LC_22_26_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_3_LC_22_26_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_3_LC_22_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32801),
            .lcout(M_this_data_tmp_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34581),
            .ce(N__34187),
            .sr(N__34019));
    defparam M_this_data_tmp_q_esr_15_LC_23_13_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_15_LC_23_13_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_15_LC_23_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_15_LC_23_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33629),
            .lcout(M_this_data_tmp_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34494),
            .ce(N__32189),
            .sr(N__34039));
    defparam M_this_data_tmp_q_esr_6_LC_23_14_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_6_LC_23_14_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_6_LC_23_14_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_6_LC_23_14_6 (
            .in0(N__32348),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34504),
            .ce(N__34199),
            .sr(N__34037));
    defparam \this_vga_signals.M_this_oam_ram_write_data_15_LC_23_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_15_LC_23_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_15_LC_23_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_15_LC_23_15_3  (
            .in0(N__35466),
            .in1(N__35230),
            .in2(N__29076),
            .in3(N__34962),
            .lcout(M_this_oam_ram_write_data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_vscroll_cry_0_c_inv_LC_23_16_0 .C_ON=1'b1;
    defparam \this_ppu.un2_vscroll_cry_0_c_inv_LC_23_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_vscroll_cry_0_c_inv_LC_23_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un2_vscroll_cry_0_c_inv_LC_23_16_0  (
            .in0(_gnd_net_),
            .in1(N__29303),
            .in2(N__29049),
            .in3(N__29199),
            .lcout(\this_ppu.M_this_oam_ram_read_data_i_16 ),
            .ltout(),
            .carryin(bfn_23_16_0_),
            .carryout(\this_ppu.un2_vscroll_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_23_16_1 .C_ON=1'b1;
    defparam \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_23_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_23_16_1  (
            .in0(_gnd_net_),
            .in1(N__31167),
            .in2(N__28722),
            .in3(N__29034),
            .lcout(\this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0 ),
            .ltout(),
            .carryin(\this_ppu.un2_vscroll_cry_0 ),
            .carryout(\this_ppu.un2_vscroll_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_23_16_2 .C_ON=1'b0;
    defparam \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_23_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_23_16_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_23_16_2  (
            .in0(N__29116),
            .in1(N__29629),
            .in2(_gnd_net_),
            .in3(N__29031),
            .lcout(\this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_12_LC_23_16_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_12_LC_23_16_6 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_12_LC_23_16_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \this_sprites_ram.mem_radreg_12_LC_23_16_6  (
            .in0(N__30161),
            .in1(N__30020),
            .in2(N__29028),
            .in3(N__31020),
            .lcout(\this_sprites_ram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34521),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIIL4G1_2_LC_23_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIIL4G1_2_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIIL4G1_2_LC_23_17_0 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_ppu.M_vaddress_q_RNIIL4G1_2_LC_23_17_0  (
            .in0(N__30002),
            .in1(N__28956),
            .in2(N__30165),
            .in3(N__29631),
            .lcout(M_this_ppu_sprites_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_2_LC_23_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_2_LC_23_17_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_2_LC_23_17_1 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \this_ppu.M_vaddress_q_2_LC_23_17_1  (
            .in0(N__29633),
            .in1(N__28720),
            .in2(N__28677),
            .in3(N__29306),
            .lcout(\this_ppu.M_vaddress_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34530),
            .ce(),
            .sr(N__29265));
    defparam \this_ppu.M_vaddress_q_3_LC_23_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_3_LC_23_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_3_LC_23_17_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_vaddress_q_3_LC_23_17_2  (
            .in0(N__29600),
            .in1(N__29557),
            .in2(_gnd_net_),
            .in3(N__29632),
            .lcout(M_this_ppu_map_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34530),
            .ce(),
            .sr(N__29265));
    defparam \this_ppu.M_vaddress_q_RNINGCA_0_LC_23_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNINGCA_0_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNINGCA_0_LC_23_17_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_ppu.M_vaddress_q_RNINGCA_0_LC_23_17_3  (
            .in0(_gnd_net_),
            .in1(N__29193),
            .in2(_gnd_net_),
            .in3(N__29304),
            .lcout(),
            .ltout(\this_ppu.un2_vscroll_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIS5A21_0_LC_23_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIS5A21_0_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIS5A21_0_LC_23_17_4 .LUT_INIT=16'b1100110010001101;
    LogicCell40 \this_ppu.M_vaddress_q_RNIS5A21_0_LC_23_17_4  (
            .in0(N__30160),
            .in1(N__29319),
            .in2(N__30024),
            .in3(N__30001),
            .lcout(M_this_ppu_sprites_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_4_LC_23_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_4_LC_23_17_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_4_LC_23_17_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \this_ppu.M_vaddress_q_4_LC_23_17_5  (
            .in0(N__29634),
            .in1(N__29601),
            .in2(N__29564),
            .in3(N__29507),
            .lcout(M_this_ppu_map_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34530),
            .ce(),
            .sr(N__29265));
    defparam \this_ppu.M_vaddress_q_0_LC_23_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_0_LC_23_17_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_0_LC_23_17_6 .LUT_INIT=16'b1010011010101010;
    LogicCell40 \this_ppu.M_vaddress_q_0_LC_23_17_6  (
            .in0(N__29305),
            .in1(N__29481),
            .in2(N__29436),
            .in3(N__29379),
            .lcout(M_this_ppu_vram_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34530),
            .ce(),
            .sr(N__29265));
    defparam M_this_oam_address_q_0_LC_23_18_5.C_ON=1'b0;
    defparam M_this_oam_address_q_0_LC_23_18_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_0_LC_23_18_5.LUT_INIT=16'b0101101000000000;
    LogicCell40 M_this_oam_address_q_0_LC_23_18_5 (
            .in0(N__34921),
            .in1(_gnd_net_),
            .in2(N__35229),
            .in3(N__30690),
            .lcout(M_this_oam_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34538),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_4_LC_23_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_4_LC_23_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_4_LC_23_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_4_LC_23_18_6  (
            .in0(N__35399),
            .in1(N__35176),
            .in2(N__29241),
            .in3(N__34920),
            .lcout(N_71_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_0_c_LC_23_19_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_0_c_LC_23_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_0_c_LC_23_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_0_c_LC_23_19_0  (
            .in0(_gnd_net_),
            .in1(N__29214),
            .in2(N__29197),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_23_19_0_),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_1_c_LC_23_19_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_1_c_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_1_c_LC_23_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_1_c_LC_23_19_1  (
            .in0(_gnd_net_),
            .in1(N__29148),
            .in2(N__31205),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_0 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_2_c_LC_23_19_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_2_c_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_2_c_LC_23_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_2_c_LC_23_19_2  (
            .in0(_gnd_net_),
            .in1(N__29133),
            .in2(N__29117),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_1 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_3_c_LC_23_19_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_3_c_LC_23_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_3_c_LC_23_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_3_c_LC_23_19_3  (
            .in0(_gnd_net_),
            .in1(N__31545),
            .in2(N__30336),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_2 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_4_c_LC_23_19_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_4_c_LC_23_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_4_c_LC_23_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_4_c_LC_23_19_4  (
            .in0(_gnd_net_),
            .in1(N__31257),
            .in2(N__30318),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_3 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_5_c_LC_23_19_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_5_c_LC_23_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_5_c_LC_23_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_5_c_LC_23_19_5  (
            .in0(_gnd_net_),
            .in1(N__31290),
            .in2(N__30300),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_4 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_6_c_LC_23_19_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_6_c_LC_23_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_6_c_LC_23_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_6_c_LC_23_19_6  (
            .in0(_gnd_net_),
            .in1(N__31373),
            .in2(N__30282),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_5 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_LC_23_19_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_LC_23_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_LC_23_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_7_c_LC_23_19_7  (
            .in0(_gnd_net_),
            .in1(N__30263),
            .in2(N__31416),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_6 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_7_THRU_LUT4_0_LC_23_20_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_THRU_LUT4_0_LC_23_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_THRU_LUT4_0_LC_23_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_7_THRU_LUT4_0_LC_23_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30246),
            .lcout(\this_ppu.un1_M_vaddress_q_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_10_LC_23_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_10_LC_23_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_10_LC_23_20_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_10_LC_23_20_1  (
            .in0(N__35430),
            .in1(N__35169),
            .in2(N__30501),
            .in3(N__34937),
            .lcout(N_61_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_3_LC_23_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_3_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_3_LC_23_20_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_3_LC_23_20_2  (
            .in0(N__34938),
            .in1(N__30222),
            .in2(N__35228),
            .in3(N__35444),
            .lcout(N_73_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_5_LC_23_20_4.C_ON=1'b0;
    defparam M_this_oam_address_q_5_LC_23_20_4.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_5_LC_23_20_4.LUT_INIT=16'b0010100010100000;
    LogicCell40 M_this_oam_address_q_5_LC_23_20_4 (
            .in0(N__30685),
            .in1(N__30191),
            .in2(N__30710),
            .in3(N__30537),
            .lcout(M_this_oam_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34551),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_3_LC_23_20_5.C_ON=1'b0;
    defparam M_this_oam_address_q_3_LC_23_20_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_3_LC_23_20_5.LUT_INIT=16'b0111100000000000;
    LogicCell40 M_this_oam_address_q_3_LC_23_20_5 (
            .in0(N__30551),
            .in1(N__30586),
            .in2(N__30635),
            .in3(N__30684),
            .lcout(M_this_oam_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34551),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNO_0_5_LC_23_20_6.C_ON=1'b0;
    defparam M_this_oam_address_q_RNO_0_5_LC_23_20_6.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNO_0_5_LC_23_20_6.LUT_INIT=16'b1000100000000000;
    LogicCell40 M_this_oam_address_q_RNO_0_5_LC_23_20_6 (
            .in0(N__30621),
            .in1(N__30581),
            .in2(_gnd_net_),
            .in3(N__30550),
            .lcout(un1_M_this_oam_address_q_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_19_LC_23_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_19_LC_23_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_19_LC_23_20_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_19_LC_23_20_7  (
            .in0(N__35445),
            .in1(N__35170),
            .in2(N__31488),
            .in3(N__34939),
            .lcout(N_50_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_21_LC_23_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_21_LC_23_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_21_LC_23_21_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_21_LC_23_21_0  (
            .in0(N__35431),
            .in1(N__35120),
            .in2(N__30510),
            .in3(N__34950),
            .lcout(N_46_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_21_LC_23_21_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_21_LC_23_21_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_21_LC_23_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_21_LC_23_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34706),
            .lcout(M_this_data_tmp_qZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34562),
            .ce(N__31445),
            .sr(N__34029));
    defparam M_this_data_tmp_q_esr_10_LC_23_22_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_10_LC_23_22_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_10_LC_23_22_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_10_LC_23_22_6 (
            .in0(N__33444),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34569),
            .ce(N__32183),
            .sr(N__34028));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_24_15_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_24_15_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_24_15_2  (
            .in0(N__30489),
            .in1(N__30477),
            .in2(_gnd_net_),
            .in3(N__30465),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_15_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_15_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_15_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_15_5  (
            .in0(N__31989),
            .in1(N__31890),
            .in2(N__31800),
            .in3(N__31671),
            .lcout(\this_sprites_ram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_24_16_4 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_24_16_4 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_24_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_LC_24_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31201),
            .lcout(M_this_oam_ram_read_data_i_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un9lto7_5_LC_24_17_0 .C_ON=1'b0;
    defparam \this_ppu.un9lto7_5_LC_24_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un9lto7_5_LC_24_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.un9lto7_5_LC_24_17_0  (
            .in0(N__31148),
            .in1(N__31127),
            .in2(N__31109),
            .in3(N__31079),
            .lcout(\this_ppu.un9lto7Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc3_LC_24_17_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc3_LC_24_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc3_LC_24_17_1 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc3_LC_24_17_1  (
            .in0(N__30774),
            .in1(N__30870),
            .in2(N__30815),
            .in3(N__30915),
            .lcout(\this_ppu.un1_M_haddress_q_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un9lto7_4_LC_24_17_3 .C_ON=1'b0;
    defparam \this_ppu.un9lto7_4_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un9lto7_4_LC_24_17_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.un9lto7_4_LC_24_17_3  (
            .in0(N__31031),
            .in1(N__31013),
            .in2(N__30995),
            .in3(N__30968),
            .lcout(\this_ppu.un9lto7Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc1_LC_24_18_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc1_LC_24_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc1_LC_24_18_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \this_ppu.un1_oam_data_axbxc1_LC_24_18_1  (
            .in0(N__31541),
            .in1(_gnd_net_),
            .in2(N__31256),
            .in3(_gnd_net_),
            .lcout(\this_ppu.un1_M_vaddress_q_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_ac0_1_LC_24_18_3 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_ac0_1_LC_24_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_ac0_1_LC_24_18_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_ac0_1_LC_24_18_3  (
            .in0(N__30905),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30861),
            .lcout(),
            .ltout(\this_ppu.un1_oam_data_1_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc4_LC_24_18_4 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc4_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc4_LC_24_18_4 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc4_LC_24_18_4  (
            .in0(N__30830),
            .in1(N__30811),
            .in2(N__30789),
            .in3(N__30775),
            .lcout(\this_ppu.un1_M_haddress_q_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_6_LC_24_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_6_LC_24_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_6_LC_24_18_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_6_LC_24_18_5  (
            .in0(N__35439),
            .in1(N__35184),
            .in2(N__30738),
            .in3(N__34923),
            .lcout(N_67_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_ac0_1_LC_24_18_6 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_ac0_1_LC_24_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_ac0_1_LC_24_18_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.un1_oam_data_ac0_1_LC_24_18_6  (
            .in0(_gnd_net_),
            .in1(N__31249),
            .in2(_gnd_net_),
            .in3(N__31540),
            .lcout(),
            .ltout(\this_ppu.un1_oam_data_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc4_LC_24_18_7 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc4_LC_24_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc4_LC_24_18_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \this_ppu.un1_oam_data_axbxc4_LC_24_18_7  (
            .in0(N__31415),
            .in1(N__31374),
            .in2(N__31395),
            .in3(N__31289),
            .lcout(\this_ppu.un1_M_vaddress_q_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_22_LC_24_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_22_LC_24_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_22_LC_24_19_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_22_LC_24_19_0  (
            .in0(N__34892),
            .in1(N__31470),
            .in2(N__35233),
            .in3(N__35423),
            .lcout(M_this_oam_ram_write_data_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc3_LC_24_19_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc3_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc3_LC_24_19_1 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.un1_oam_data_axbxc3_LC_24_19_1  (
            .in0(N__31248),
            .in1(N__31282),
            .in2(N__31372),
            .in3(N__31536),
            .lcout(\this_ppu.un1_M_vaddress_q_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_31_LC_24_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_31_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_31_LC_24_19_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_31_LC_24_19_2  (
            .in0(N__34890),
            .in1(N__33668),
            .in2(N__35231),
            .in3(N__35421),
            .lcout(M_this_oam_ram_write_data_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_18_LC_24_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_18_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_18_LC_24_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_18_LC_24_19_3  (
            .in0(N__35420),
            .in1(N__35200),
            .in2(N__31479),
            .in3(N__34893),
            .lcout(N_52_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_16_LC_24_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_16_LC_24_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_16_LC_24_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_16_LC_24_19_4  (
            .in0(N__34891),
            .in1(N__31494),
            .in2(N__35232),
            .in3(N__35422),
            .lcout(M_this_oam_ram_write_data_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_i_o3_LC_24_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_i_o3_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_i_o3_LC_24_19_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_i_o3_LC_24_19_5  (
            .in0(N__35419),
            .in1(N__35190),
            .in2(_gnd_net_),
            .in3(N__34889),
            .lcout(N_158_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc2_LC_24_19_6 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc2_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc2_LC_24_19_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.un1_oam_data_axbxc2_LC_24_19_6  (
            .in0(N__31535),
            .in1(N__31278),
            .in2(_gnd_net_),
            .in3(N__31247),
            .lcout(\this_ppu.un1_M_vaddress_q_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_24_19_7 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_24_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_24_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31534),
            .lcout(M_this_oam_ram_read_data_i_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_16_LC_24_20_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_16_LC_24_20_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_16_LC_24_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_16_LC_24_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33825),
            .lcout(M_this_data_tmp_qZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34563),
            .ce(N__31438),
            .sr(N__34031));
    defparam M_this_data_tmp_q_esr_19_LC_24_20_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_19_LC_24_20_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_19_LC_24_20_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_19_LC_24_20_2 (
            .in0(N__32835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34563),
            .ce(N__31438),
            .sr(N__34031));
    defparam M_this_data_tmp_q_esr_18_LC_24_20_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_18_LC_24_20_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_18_LC_24_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_18_LC_24_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33472),
            .lcout(M_this_data_tmp_qZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34563),
            .ce(N__31438),
            .sr(N__34031));
    defparam M_this_data_tmp_q_esr_22_LC_24_20_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_22_LC_24_20_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_22_LC_24_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_22_LC_24_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32331),
            .lcout(M_this_data_tmp_qZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34563),
            .ce(N__31438),
            .sr(N__34031));
    defparam M_this_data_tmp_q_esr_23_LC_24_20_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_23_LC_24_20_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_23_LC_24_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_23_LC_24_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33669),
            .lcout(M_this_data_tmp_qZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34563),
            .ce(N__31438),
            .sr(N__34031));
    defparam M_this_data_tmp_q_esr_17_LC_24_20_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_17_LC_24_20_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_17_LC_24_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_17_LC_24_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32981),
            .lcout(M_this_data_tmp_qZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34563),
            .ce(N__31438),
            .sr(N__34031));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_17_LC_24_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_17_LC_24_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_17_LC_24_21_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_17_LC_24_21_1  (
            .in0(N__35429),
            .in1(N__35122),
            .in2(N__31464),
            .in3(N__34953),
            .lcout(N_54_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI13IA1_1_LC_24_21_4.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI13IA1_1_LC_24_21_4.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI13IA1_1_LC_24_21_4.LUT_INIT=16'b1111111101000000;
    LogicCell40 M_this_oam_address_q_RNI13IA1_1_LC_24_21_4 (
            .in0(N__34951),
            .in1(N__35427),
            .in2(N__35183),
            .in3(N__34117),
            .lcout(N_1126_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_30_LC_24_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_30_LC_24_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_30_LC_24_21_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_30_LC_24_21_5  (
            .in0(N__35428),
            .in1(N__35121),
            .in2(N__32352),
            .in3(N__34952),
            .lcout(M_this_oam_ram_write_data_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_0_c_LC_24_22_0.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_0_c_LC_24_22_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_0_c_LC_24_22_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_external_address_q_cry_0_c_LC_24_22_0 (
            .in0(_gnd_net_),
            .in1(N__33296),
            .in2(N__33272),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_24_22_0_),
            .carryout(un1_M_this_external_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_0_THRU_LUT4_0_LC_24_22_1.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_0_THRU_LUT4_0_LC_24_22_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_0_THRU_LUT4_0_LC_24_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_external_address_q_cry_0_THRU_LUT4_0_LC_24_22_1 (
            .in0(_gnd_net_),
            .in1(N__33222),
            .in2(_gnd_net_),
            .in3(N__31566),
            .lcout(un1_M_this_external_address_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_0),
            .carryout(un1_M_this_external_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_1_THRU_LUT4_0_LC_24_22_2.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_1_THRU_LUT4_0_LC_24_22_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_1_THRU_LUT4_0_LC_24_22_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_external_address_q_cry_1_THRU_LUT4_0_LC_24_22_2 (
            .in0(_gnd_net_),
            .in1(N__33173),
            .in2(_gnd_net_),
            .in3(N__31563),
            .lcout(un1_M_this_external_address_q_cry_1_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_1),
            .carryout(un1_M_this_external_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_2_THRU_LUT4_0_LC_24_22_3.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_2_THRU_LUT4_0_LC_24_22_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_2_THRU_LUT4_0_LC_24_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_external_address_q_cry_2_THRU_LUT4_0_LC_24_22_3 (
            .in0(_gnd_net_),
            .in1(N__33125),
            .in2(_gnd_net_),
            .in3(N__31560),
            .lcout(un1_M_this_external_address_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_2),
            .carryout(un1_M_this_external_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_3_THRU_LUT4_0_LC_24_22_4.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_3_THRU_LUT4_0_LC_24_22_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_3_THRU_LUT4_0_LC_24_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_external_address_q_cry_3_THRU_LUT4_0_LC_24_22_4 (
            .in0(_gnd_net_),
            .in1(N__33084),
            .in2(_gnd_net_),
            .in3(N__31557),
            .lcout(un1_M_this_external_address_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_3),
            .carryout(un1_M_this_external_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_4_THRU_LUT4_0_LC_24_22_5.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_4_THRU_LUT4_0_LC_24_22_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_4_THRU_LUT4_0_LC_24_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_external_address_q_cry_4_THRU_LUT4_0_LC_24_22_5 (
            .in0(_gnd_net_),
            .in1(N__33038),
            .in2(_gnd_net_),
            .in3(N__31554),
            .lcout(un1_M_this_external_address_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_4),
            .carryout(un1_M_this_external_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_5_THRU_LUT4_0_LC_24_22_6.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_5_THRU_LUT4_0_LC_24_22_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_5_THRU_LUT4_0_LC_24_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_external_address_q_cry_5_THRU_LUT4_0_LC_24_22_6 (
            .in0(_gnd_net_),
            .in1(N__35519),
            .in2(_gnd_net_),
            .in3(N__31551),
            .lcout(un1_M_this_external_address_q_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_5),
            .carryout(un1_M_this_external_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_6_THRU_LUT4_0_LC_24_22_7.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_6_THRU_LUT4_0_LC_24_22_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_6_THRU_LUT4_0_LC_24_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_external_address_q_cry_6_THRU_LUT4_0_LC_24_22_7 (
            .in0(_gnd_net_),
            .in1(N__32635),
            .in2(_gnd_net_),
            .in3(N__31548),
            .lcout(un1_M_this_external_address_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_6),
            .carryout(un1_M_this_external_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_7_c_RNIU5OB_LC_24_23_0.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_7_c_RNIU5OB_LC_24_23_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_7_c_RNIU5OB_LC_24_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_7_c_RNIU5OB_LC_24_23_0 (
            .in0(_gnd_net_),
            .in1(N__33695),
            .in2(_gnd_net_),
            .in3(N__32046),
            .lcout(un1_M_this_external_address_q_cry_7_c_RNIU5OBZ0),
            .ltout(),
            .carryin(bfn_24_23_0_),
            .carryout(un1_M_this_external_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_8_c_RNI09PB_LC_24_23_1.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_8_c_RNI09PB_LC_24_23_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_8_c_RNI09PB_LC_24_23_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_8_c_RNI09PB_LC_24_23_1 (
            .in0(_gnd_net_),
            .in1(N__32033),
            .in2(_gnd_net_),
            .in3(N__32010),
            .lcout(un1_M_this_external_address_q_cry_8_c_RNI09PBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_8),
            .carryout(un1_M_this_external_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_9_c_RNI9RGK_LC_24_23_2.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_9_c_RNI9RGK_LC_24_23_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_9_c_RNI9RGK_LC_24_23_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_9_c_RNI9RGK_LC_24_23_2 (
            .in0(_gnd_net_),
            .in1(N__33317),
            .in2(_gnd_net_),
            .in3(N__32007),
            .lcout(un1_M_this_external_address_q_cry_9_c_RNI9RGKZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_9),
            .carryout(un1_M_this_external_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_10_c_RNIIOGB_LC_24_23_3.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_10_c_RNIIOGB_LC_24_23_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_10_c_RNIIOGB_LC_24_23_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_10_c_RNIIOGB_LC_24_23_3 (
            .in0(_gnd_net_),
            .in1(N__32684),
            .in2(_gnd_net_),
            .in3(N__32004),
            .lcout(un1_M_this_external_address_q_cry_10_c_RNIIOGBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_10),
            .carryout(un1_M_this_external_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_11_c_RNIKRHB_LC_24_23_4.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_11_c_RNIKRHB_LC_24_23_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_11_c_RNIKRHB_LC_24_23_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_11_c_RNIKRHB_LC_24_23_4 (
            .in0(_gnd_net_),
            .in1(N__32480),
            .in2(_gnd_net_),
            .in3(N__32001),
            .lcout(un1_M_this_external_address_q_cry_11_c_RNIKRHBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_11),
            .carryout(un1_M_this_external_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_12_c_RNIMUIB_LC_24_23_5.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_12_c_RNIMUIB_LC_24_23_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_12_c_RNIMUIB_LC_24_23_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_12_c_RNIMUIB_LC_24_23_5 (
            .in0(_gnd_net_),
            .in1(N__32444),
            .in2(_gnd_net_),
            .in3(N__31998),
            .lcout(un1_M_this_external_address_q_cry_12_c_RNIMUIBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_12),
            .carryout(un1_M_this_external_address_q_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_13_c_RNIO1KB_LC_24_23_6.C_ON=1'b1;
    defparam un1_M_this_external_address_q_cry_13_c_RNIO1KB_LC_24_23_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_13_c_RNIO1KB_LC_24_23_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_external_address_q_cry_13_c_RNIO1KB_LC_24_23_6 (
            .in0(_gnd_net_),
            .in1(N__32270),
            .in2(_gnd_net_),
            .in3(N__31995),
            .lcout(un1_M_this_external_address_q_cry_13_c_RNIO1KBZ0),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_13),
            .carryout(un1_M_this_external_address_q_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_external_address_q_cry_14_c_RNIQ4LB_LC_24_23_7.C_ON=1'b0;
    defparam un1_M_this_external_address_q_cry_14_c_RNIQ4LB_LC_24_23_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_external_address_q_cry_14_c_RNIQ4LB_LC_24_23_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_M_this_external_address_q_cry_14_c_RNIQ4LB_LC_24_23_7 (
            .in0(_gnd_net_),
            .in1(N__33524),
            .in2(_gnd_net_),
            .in3(N__31992),
            .lcout(un1_M_this_external_address_q_cry_14_c_RNIQ4LBZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_24_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_24_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_24_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_24_5  (
            .in0(N__31984),
            .in1(N__31885),
            .in2(N__31795),
            .in3(N__31667),
            .lcout(\this_sprites_ram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_8_LC_26_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_8_LC_26_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_8_LC_26_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_8_LC_26_16_6  (
            .in0(N__35247),
            .in1(N__35483),
            .in2(N__32109),
            .in3(N__35002),
            .lcout(M_this_oam_ram_write_data_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_8_LC_26_16_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_8_LC_26_16_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_8_LC_26_16_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_8_LC_26_16_7 (
            .in0(N__33826),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34548),
            .ce(N__32184),
            .sr(N__34040));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_0_LC_26_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_0_LC_26_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_0_LC_26_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_0_LC_26_17_0  (
            .in0(N__35486),
            .in1(N__35239),
            .in2(N__32094),
            .in3(N__34990),
            .lcout(N_79_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_0_LC_26_17_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_0_LC_26_17_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_0_LC_26_17_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_0_LC_26_17_1 (
            .in0(N__33813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34552),
            .ce(N__34200),
            .sr(N__34038));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_24_LC_26_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_24_LC_26_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_24_LC_26_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_24_LC_26_17_2  (
            .in0(N__35484),
            .in1(N__35246),
            .in2(N__35004),
            .in3(N__33814),
            .lcout(N_43_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_1_LC_26_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_1_LC_26_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_1_LC_26_17_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_1_LC_26_17_3  (
            .in0(N__34988),
            .in1(N__32064),
            .in2(N__35250),
            .in3(N__35485),
            .lcout(N_77_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_1_LC_26_17_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_1_LC_26_17_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_1_LC_26_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_1_LC_26_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32987),
            .lcout(M_this_data_tmp_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34552),
            .ce(N__34200),
            .sr(N__34038));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_12_LC_26_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_12_LC_26_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_12_LC_26_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_12_LC_26_17_7  (
            .in0(N__34989),
            .in1(N__32220),
            .in2(N__35249),
            .in3(N__35487),
            .lcout(N_58_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_14_LC_26_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_14_LC_26_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_14_LC_26_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_14_LC_26_18_2  (
            .in0(N__35441),
            .in1(N__35186),
            .in2(N__32202),
            .in3(N__34980),
            .lcout(M_this_oam_ram_write_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_9_LC_26_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_9_LC_26_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_9_LC_26_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_9_LC_26_18_3  (
            .in0(N__34978),
            .in1(N__35443),
            .in2(N__32211),
            .in3(N__35188),
            .lcout(N_63_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_2_LC_26_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_2_LC_26_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_2_LC_26_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_2_LC_26_18_4  (
            .in0(N__35442),
            .in1(N__35187),
            .in2(N__32859),
            .in3(N__34981),
            .lcout(N_75_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_11_LC_26_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_11_LC_26_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_11_LC_26_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_11_LC_26_18_6  (
            .in0(N__35440),
            .in1(N__35185),
            .in2(N__32229),
            .in3(N__34979),
            .lcout(M_this_oam_ram_write_data_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_11_LC_26_19_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_11_LC_26_19_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_11_LC_26_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_11_LC_26_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32831),
            .lcout(M_this_data_tmp_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34570),
            .ce(N__32190),
            .sr(N__34034));
    defparam M_this_data_tmp_q_esr_12_LC_26_19_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_12_LC_26_19_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_12_LC_26_19_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_12_LC_26_19_1 (
            .in0(N__32529),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34570),
            .ce(N__32190),
            .sr(N__34034));
    defparam M_this_data_tmp_q_esr_9_LC_26_19_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_9_LC_26_19_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_9_LC_26_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_9_LC_26_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32988),
            .lcout(M_this_data_tmp_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34570),
            .ce(N__32190),
            .sr(N__34034));
    defparam M_this_data_tmp_q_esr_14_LC_26_19_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_14_LC_26_19_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_14_LC_26_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_14_LC_26_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32388),
            .lcout(M_this_data_tmp_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34570),
            .ce(N__32190),
            .sr(N__34034));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_26_LC_26_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_26_LC_26_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_26_LC_26_20_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_26_LC_26_20_0  (
            .in0(N__35237),
            .in1(N__35481),
            .in2(N__33421),
            .in3(N__35001),
            .lcout(N_39_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_27_LC_26_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_27_LC_26_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_27_LC_26_20_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_27_LC_26_20_2  (
            .in0(N__35235),
            .in1(N__35480),
            .in2(N__32830),
            .in3(N__35000),
            .lcout(M_this_oam_ram_write_data_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_23_LC_26_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_23_LC_26_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_23_LC_26_20_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_23_LC_26_20_4  (
            .in0(N__35234),
            .in1(N__35479),
            .in2(N__33006),
            .in3(N__34999),
            .lcout(M_this_oam_ram_write_data_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_25_LC_26_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_25_LC_26_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_25_LC_26_20_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_25_LC_26_20_7  (
            .in0(N__34998),
            .in1(N__35482),
            .in2(N__32986),
            .in3(N__35236),
            .lcout(N_41_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_2_LC_26_21_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_2_LC_26_21_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_2_LC_26_21_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_2_LC_26_21_2 (
            .in0(N__33394),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34576),
            .ce(N__34162),
            .sr(N__34033));
    defparam M_this_external_address_q_11_LC_26_22_0.C_ON=1'b0;
    defparam M_this_external_address_q_11_LC_26_22_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_11_LC_26_22_0.LUT_INIT=16'b1110010011001100;
    LogicCell40 M_this_external_address_q_11_LC_26_22_0 (
            .in0(N__35634),
            .in1(N__32847),
            .in2(N__32834),
            .in3(N__35856),
            .lcout(M_this_external_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__34032));
    defparam M_this_external_address_q_7_LC_26_22_1.C_ON=1'b0;
    defparam M_this_external_address_q_7_LC_26_22_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_7_LC_26_22_1.LUT_INIT=16'b0000011101110000;
    LogicCell40 M_this_external_address_q_7_LC_26_22_1 (
            .in0(N__35855),
            .in1(N__35640),
            .in2(N__32636),
            .in3(N__32661),
            .lcout(M_this_external_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__34032));
    defparam M_this_external_address_q_12_LC_26_22_2.C_ON=1'b0;
    defparam M_this_external_address_q_12_LC_26_22_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_12_LC_26_22_2.LUT_INIT=16'b1110010011001100;
    LogicCell40 M_this_external_address_q_12_LC_26_22_2 (
            .in0(N__35635),
            .in1(N__32610),
            .in2(N__32547),
            .in3(N__35857),
            .lcout(M_this_external_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__34032));
    defparam M_this_external_address_q_13_LC_26_22_3.C_ON=1'b0;
    defparam M_this_external_address_q_13_LC_26_22_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_13_LC_26_22_3.LUT_INIT=16'b1111011110000000;
    LogicCell40 M_this_external_address_q_13_LC_26_22_3 (
            .in0(N__35853),
            .in1(N__35638),
            .in2(N__34694),
            .in3(N__32457),
            .lcout(M_this_external_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__34032));
    defparam M_this_external_address_q_14_LC_26_22_4.C_ON=1'b0;
    defparam M_this_external_address_q_14_LC_26_22_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_14_LC_26_22_4.LUT_INIT=16'b1110010011001100;
    LogicCell40 M_this_external_address_q_14_LC_26_22_4 (
            .in0(N__35636),
            .in1(N__32421),
            .in2(N__32407),
            .in3(N__35858),
            .lcout(M_this_external_address_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__34032));
    defparam M_this_external_address_q_8_LC_26_22_6.C_ON=1'b0;
    defparam M_this_external_address_q_8_LC_26_22_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_8_LC_26_22_6.LUT_INIT=16'b1110010011001100;
    LogicCell40 M_this_external_address_q_8_LC_26_22_6 (
            .in0(N__35637),
            .in1(N__33846),
            .in2(N__33834),
            .in3(N__35859),
            .lcout(M_this_external_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__34032));
    defparam M_this_external_address_q_15_LC_26_22_7.C_ON=1'b0;
    defparam M_this_external_address_q_15_LC_26_22_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_15_LC_26_22_7.LUT_INIT=16'b1111011110000000;
    LogicCell40 M_this_external_address_q_15_LC_26_22_7 (
            .in0(N__35854),
            .in1(N__35639),
            .in2(N__33637),
            .in3(N__33546),
            .lcout(M_this_external_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34584),
            .ce(),
            .sr(N__34032));
    defparam M_this_external_address_q_10_LC_26_23_0.C_ON=1'b0;
    defparam M_this_external_address_q_10_LC_26_23_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_10_LC_26_23_0.LUT_INIT=16'b1110010011001100;
    LogicCell40 M_this_external_address_q_10_LC_26_23_0 (
            .in0(N__35611),
            .in1(N__33501),
            .in2(N__33420),
            .in3(N__35864),
            .lcout(M_this_external_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__34030));
    defparam M_this_external_address_q_0_LC_26_23_1.C_ON=1'b0;
    defparam M_this_external_address_q_0_LC_26_23_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_0_LC_26_23_1.LUT_INIT=16'b0000011101110000;
    LogicCell40 M_this_external_address_q_0_LC_26_23_1 (
            .in0(N__35860),
            .in1(N__35615),
            .in2(N__33262),
            .in3(N__33303),
            .lcout(M_this_external_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__34030));
    defparam M_this_external_address_q_1_LC_26_23_2.C_ON=1'b0;
    defparam M_this_external_address_q_1_LC_26_23_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_1_LC_26_23_2.LUT_INIT=16'b0001010000111100;
    LogicCell40 M_this_external_address_q_1_LC_26_23_2 (
            .in0(N__35612),
            .in1(N__33234),
            .in2(N__33220),
            .in3(N__35865),
            .lcout(M_this_external_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__34030));
    defparam M_this_external_address_q_2_LC_26_23_3.C_ON=1'b0;
    defparam M_this_external_address_q_2_LC_26_23_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_2_LC_26_23_3.LUT_INIT=16'b0000011101110000;
    LogicCell40 M_this_external_address_q_2_LC_26_23_3 (
            .in0(N__35861),
            .in1(N__35616),
            .in2(N__33172),
            .in3(N__33192),
            .lcout(M_this_external_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__34030));
    defparam M_this_external_address_q_3_LC_26_23_4.C_ON=1'b0;
    defparam M_this_external_address_q_3_LC_26_23_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_3_LC_26_23_4.LUT_INIT=16'b0001010000111100;
    LogicCell40 M_this_external_address_q_3_LC_26_23_4 (
            .in0(N__35613),
            .in1(N__33144),
            .in2(N__33124),
            .in3(N__35866),
            .lcout(M_this_external_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__34030));
    defparam M_this_external_address_q_4_LC_26_23_5.C_ON=1'b0;
    defparam M_this_external_address_q_4_LC_26_23_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_4_LC_26_23_5.LUT_INIT=16'b0000011101110000;
    LogicCell40 M_this_external_address_q_4_LC_26_23_5 (
            .in0(N__35862),
            .in1(N__35617),
            .in2(N__33082),
            .in3(N__33096),
            .lcout(M_this_external_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__34030));
    defparam M_this_external_address_q_5_LC_26_23_6.C_ON=1'b0;
    defparam M_this_external_address_q_5_LC_26_23_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_5_LC_26_23_6.LUT_INIT=16'b0001010000111100;
    LogicCell40 M_this_external_address_q_5_LC_26_23_6 (
            .in0(N__35614),
            .in1(N__33054),
            .in2(N__33034),
            .in3(N__35867),
            .lcout(M_this_external_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__34030));
    defparam M_this_external_address_q_6_LC_26_23_7.C_ON=1'b0;
    defparam M_this_external_address_q_6_LC_26_23_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_6_LC_26_23_7.LUT_INIT=16'b0000011101110000;
    LogicCell40 M_this_external_address_q_6_LC_26_23_7 (
            .in0(N__35863),
            .in1(N__35618),
            .in2(N__35515),
            .in3(N__35538),
            .lcout(M_this_external_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34585),
            .ce(),
            .sr(N__34030));
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_5_LC_27_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_5_LC_27_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_i_5_LC_27_19_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_i_5_LC_27_19_0  (
            .in0(N__35468),
            .in1(N__35238),
            .in2(N__34605),
            .in3(N__34997),
            .lcout(N_69_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_5_LC_27_20_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_5_LC_27_20_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_5_LC_27_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_5_LC_27_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34664),
            .lcout(M_this_data_tmp_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34577),
            .ce(N__34188),
            .sr(N__34035));
endmodule // cu_top_0
